magic
tech sky130A
magscale 1 2
timestamp 1730699969
<< error_p >>
rect 3138 3262 3208 3292
<< nwell >>
rect -102 3892 3200 4460
<< pwell >>
rect -102 3332 3200 3890
rect -142 3232 3208 3262
<< nmos >>
rect 94 3542 124 3742
rect 414 3542 444 3742
rect 734 3542 764 3742
rect 1054 3542 1084 3742
rect 1374 3542 1404 3742
rect 1694 3542 1724 3742
rect 2014 3542 2044 3742
rect 2334 3542 2364 3742
rect 2654 3542 2684 3742
rect 2974 3542 3004 3742
<< pmos >>
rect 94 4040 124 4240
rect 414 4040 444 4240
rect 734 4040 764 4240
rect 1054 4040 1084 4240
rect 1374 4040 1404 4240
rect 1694 4040 1724 4240
rect 2014 4040 2044 4240
rect 2334 4040 2364 4240
rect 2654 4040 2684 4240
rect 2974 4040 3004 4240
<< ndiff >>
rect 36 3730 94 3742
rect 36 3554 48 3730
rect 82 3554 94 3730
rect 36 3542 94 3554
rect 124 3730 182 3742
rect 124 3554 136 3730
rect 170 3554 182 3730
rect 124 3542 182 3554
rect 356 3730 414 3742
rect 356 3554 368 3730
rect 402 3554 414 3730
rect 356 3542 414 3554
rect 444 3730 502 3742
rect 444 3554 456 3730
rect 490 3554 502 3730
rect 444 3542 502 3554
rect 676 3730 734 3742
rect 676 3554 688 3730
rect 722 3554 734 3730
rect 676 3542 734 3554
rect 764 3730 822 3742
rect 764 3554 776 3730
rect 810 3554 822 3730
rect 764 3542 822 3554
rect 996 3730 1054 3742
rect 996 3554 1008 3730
rect 1042 3554 1054 3730
rect 996 3542 1054 3554
rect 1084 3730 1142 3742
rect 1084 3554 1096 3730
rect 1130 3554 1142 3730
rect 1084 3542 1142 3554
rect 1316 3730 1374 3742
rect 1316 3554 1328 3730
rect 1362 3554 1374 3730
rect 1316 3542 1374 3554
rect 1404 3730 1462 3742
rect 1404 3554 1416 3730
rect 1450 3554 1462 3730
rect 1404 3542 1462 3554
rect 1636 3730 1694 3742
rect 1636 3554 1648 3730
rect 1682 3554 1694 3730
rect 1636 3542 1694 3554
rect 1724 3730 1782 3742
rect 1724 3554 1736 3730
rect 1770 3554 1782 3730
rect 1724 3542 1782 3554
rect 1956 3730 2014 3742
rect 1956 3554 1968 3730
rect 2002 3554 2014 3730
rect 1956 3542 2014 3554
rect 2044 3730 2102 3742
rect 2044 3554 2056 3730
rect 2090 3554 2102 3730
rect 2044 3542 2102 3554
rect 2276 3730 2334 3742
rect 2276 3554 2288 3730
rect 2322 3554 2334 3730
rect 2276 3542 2334 3554
rect 2364 3730 2422 3742
rect 2364 3554 2376 3730
rect 2410 3554 2422 3730
rect 2364 3542 2422 3554
rect 2596 3730 2654 3742
rect 2596 3554 2608 3730
rect 2642 3554 2654 3730
rect 2596 3542 2654 3554
rect 2684 3730 2742 3742
rect 2684 3554 2696 3730
rect 2730 3554 2742 3730
rect 2684 3542 2742 3554
rect 2916 3730 2974 3742
rect 2916 3554 2928 3730
rect 2962 3554 2974 3730
rect 2916 3542 2974 3554
rect 3004 3730 3062 3742
rect 3004 3554 3016 3730
rect 3050 3554 3062 3730
rect 3004 3542 3062 3554
<< pdiff >>
rect 36 4228 94 4240
rect 36 4052 48 4228
rect 82 4052 94 4228
rect 36 4040 94 4052
rect 124 4228 182 4240
rect 124 4052 136 4228
rect 170 4052 182 4228
rect 124 4040 182 4052
rect 356 4228 414 4240
rect 356 4052 368 4228
rect 402 4052 414 4228
rect 356 4040 414 4052
rect 444 4228 502 4240
rect 444 4052 456 4228
rect 490 4052 502 4228
rect 444 4040 502 4052
rect 676 4228 734 4240
rect 676 4052 688 4228
rect 722 4052 734 4228
rect 676 4040 734 4052
rect 764 4228 822 4240
rect 764 4052 776 4228
rect 810 4052 822 4228
rect 764 4040 822 4052
rect 996 4228 1054 4240
rect 996 4052 1008 4228
rect 1042 4052 1054 4228
rect 996 4040 1054 4052
rect 1084 4228 1142 4240
rect 1084 4052 1096 4228
rect 1130 4052 1142 4228
rect 1084 4040 1142 4052
rect 1316 4228 1374 4240
rect 1316 4052 1328 4228
rect 1362 4052 1374 4228
rect 1316 4040 1374 4052
rect 1404 4228 1462 4240
rect 1404 4052 1416 4228
rect 1450 4052 1462 4228
rect 1404 4040 1462 4052
rect 1636 4228 1694 4240
rect 1636 4052 1648 4228
rect 1682 4052 1694 4228
rect 1636 4040 1694 4052
rect 1724 4228 1782 4240
rect 1724 4052 1736 4228
rect 1770 4052 1782 4228
rect 1724 4040 1782 4052
rect 1956 4228 2014 4240
rect 1956 4052 1968 4228
rect 2002 4052 2014 4228
rect 1956 4040 2014 4052
rect 2044 4228 2102 4240
rect 2044 4052 2056 4228
rect 2090 4052 2102 4228
rect 2044 4040 2102 4052
rect 2276 4228 2334 4240
rect 2276 4052 2288 4228
rect 2322 4052 2334 4228
rect 2276 4040 2334 4052
rect 2364 4228 2422 4240
rect 2364 4052 2376 4228
rect 2410 4052 2422 4228
rect 2364 4040 2422 4052
rect 2596 4228 2654 4240
rect 2596 4052 2608 4228
rect 2642 4052 2654 4228
rect 2596 4040 2654 4052
rect 2684 4228 2742 4240
rect 2684 4052 2696 4228
rect 2730 4052 2742 4228
rect 2684 4040 2742 4052
rect 2916 4228 2974 4240
rect 2916 4052 2928 4228
rect 2962 4052 2974 4228
rect 2916 4040 2974 4052
rect 3004 4228 3062 4240
rect 3004 4052 3016 4228
rect 3050 4052 3062 4228
rect 3004 4040 3062 4052
<< ndiffc >>
rect 48 3554 82 3730
rect 136 3554 170 3730
rect 368 3554 402 3730
rect 456 3554 490 3730
rect 688 3554 722 3730
rect 776 3554 810 3730
rect 1008 3554 1042 3730
rect 1096 3554 1130 3730
rect 1328 3554 1362 3730
rect 1416 3554 1450 3730
rect 1648 3554 1682 3730
rect 1736 3554 1770 3730
rect 1968 3554 2002 3730
rect 2056 3554 2090 3730
rect 2288 3554 2322 3730
rect 2376 3554 2410 3730
rect 2608 3554 2642 3730
rect 2696 3554 2730 3730
rect 2928 3554 2962 3730
rect 3016 3554 3050 3730
<< pdiffc >>
rect 48 4052 82 4228
rect 136 4052 170 4228
rect 368 4052 402 4228
rect 456 4052 490 4228
rect 688 4052 722 4228
rect 776 4052 810 4228
rect 1008 4052 1042 4228
rect 1096 4052 1130 4228
rect 1328 4052 1362 4228
rect 1416 4052 1450 4228
rect 1648 4052 1682 4228
rect 1736 4052 1770 4228
rect 1968 4052 2002 4228
rect 2056 4052 2090 4228
rect 2288 4052 2322 4228
rect 2376 4052 2410 4228
rect 2608 4052 2642 4228
rect 2696 4052 2730 4228
rect 2928 4052 2962 4228
rect 3016 4052 3050 4228
<< psubdiff >>
rect -66 3820 3164 3854
rect -66 3402 -32 3820
rect 250 3402 288 3820
rect 570 3402 608 3820
rect 890 3402 928 3820
rect 1210 3402 1248 3820
rect 1530 3402 1568 3820
rect 1850 3402 1888 3820
rect 2170 3402 2208 3820
rect 2490 3402 2528 3820
rect 2810 3402 2848 3820
rect 3130 3402 3164 3820
rect -66 3368 30 3402
rect 188 3368 350 3402
rect 508 3368 670 3402
rect 828 3368 990 3402
rect 1148 3368 1310 3402
rect 1468 3368 1630 3402
rect 1788 3368 1950 3402
rect 2108 3368 2270 3402
rect 2428 3368 2590 3402
rect 2748 3368 2910 3402
rect 3068 3368 3164 3402
<< nsubdiff >>
rect -66 4390 30 4424
rect 188 4390 350 4424
rect 508 4390 670 4424
rect 828 4390 990 4424
rect 1148 4390 1310 4424
rect 1468 4390 1630 4424
rect 1788 4390 1950 4424
rect 2108 4390 2270 4424
rect 2428 4390 2590 4424
rect 2748 4390 2910 4424
rect 3068 4390 3164 4424
rect -66 3962 -32 4390
rect 250 3962 288 4390
rect 570 3962 608 4390
rect 890 3962 928 4390
rect 1210 3962 1248 4390
rect 1530 3962 1568 4390
rect 1850 3962 1888 4390
rect 2170 3962 2208 4390
rect 2490 3962 2528 4390
rect 2810 3962 2848 4390
rect 3130 3962 3164 4390
rect -66 3928 3164 3962
<< psubdiffcont >>
rect 30 3368 188 3402
rect 350 3368 508 3402
rect 670 3368 828 3402
rect 990 3368 1148 3402
rect 1310 3368 1468 3402
rect 1630 3368 1788 3402
rect 1950 3368 2108 3402
rect 2270 3368 2428 3402
rect 2590 3368 2748 3402
rect 2910 3368 3068 3402
<< nsubdiffcont >>
rect 30 4390 188 4424
rect 350 4390 508 4424
rect 670 4390 828 4424
rect 990 4390 1148 4424
rect 1310 4390 1468 4424
rect 1630 4390 1788 4424
rect 1950 4390 2108 4424
rect 2270 4390 2428 4424
rect 2590 4390 2748 4424
rect 2910 4390 3068 4424
<< poly >>
rect 76 4321 142 4337
rect 76 4287 92 4321
rect 126 4287 142 4321
rect 76 4271 142 4287
rect 94 4240 124 4271
rect 94 4014 124 4040
rect 396 4321 462 4337
rect 396 4287 412 4321
rect 446 4287 462 4321
rect 396 4271 462 4287
rect 414 4240 444 4271
rect 414 4014 444 4040
rect 716 4321 782 4337
rect 716 4287 732 4321
rect 766 4287 782 4321
rect 716 4271 782 4287
rect 734 4240 764 4271
rect 734 4014 764 4040
rect 1036 4321 1102 4337
rect 1036 4287 1052 4321
rect 1086 4287 1102 4321
rect 1036 4271 1102 4287
rect 1054 4240 1084 4271
rect 1054 4014 1084 4040
rect 1356 4321 1422 4337
rect 1356 4287 1372 4321
rect 1406 4287 1422 4321
rect 1356 4271 1422 4287
rect 1374 4240 1404 4271
rect 1374 4014 1404 4040
rect 1676 4321 1742 4337
rect 1676 4287 1692 4321
rect 1726 4287 1742 4321
rect 1676 4271 1742 4287
rect 1694 4240 1724 4271
rect 1694 4014 1724 4040
rect 1996 4321 2062 4337
rect 1996 4287 2012 4321
rect 2046 4287 2062 4321
rect 1996 4271 2062 4287
rect 2014 4240 2044 4271
rect 2014 4014 2044 4040
rect 2316 4321 2382 4337
rect 2316 4287 2332 4321
rect 2366 4287 2382 4321
rect 2316 4271 2382 4287
rect 2334 4240 2364 4271
rect 2334 4014 2364 4040
rect 2636 4321 2702 4337
rect 2636 4287 2652 4321
rect 2686 4287 2702 4321
rect 2636 4271 2702 4287
rect 2654 4240 2684 4271
rect 2654 4014 2684 4040
rect 2956 4321 3022 4337
rect 2956 4287 2972 4321
rect 3006 4287 3022 4321
rect 2956 4271 3022 4287
rect 2974 4240 3004 4271
rect 2974 4014 3004 4040
rect 94 3742 124 3768
rect 94 3520 124 3542
rect 76 3504 142 3520
rect 76 3470 92 3504
rect 126 3470 142 3504
rect 76 3454 142 3470
rect 414 3742 444 3768
rect 414 3520 444 3542
rect 396 3504 462 3520
rect 396 3470 412 3504
rect 446 3470 462 3504
rect 396 3454 462 3470
rect 734 3742 764 3768
rect 734 3520 764 3542
rect 716 3504 782 3520
rect 716 3470 732 3504
rect 766 3470 782 3504
rect 716 3454 782 3470
rect 1054 3742 1084 3768
rect 1054 3520 1084 3542
rect 1036 3504 1102 3520
rect 1036 3470 1052 3504
rect 1086 3470 1102 3504
rect 1036 3454 1102 3470
rect 1374 3742 1404 3768
rect 1374 3520 1404 3542
rect 1356 3504 1422 3520
rect 1356 3470 1372 3504
rect 1406 3470 1422 3504
rect 1356 3454 1422 3470
rect 1694 3742 1724 3768
rect 1694 3520 1724 3542
rect 1676 3504 1742 3520
rect 1676 3470 1692 3504
rect 1726 3470 1742 3504
rect 1676 3454 1742 3470
rect 2014 3742 2044 3768
rect 2014 3520 2044 3542
rect 1996 3504 2062 3520
rect 1996 3470 2012 3504
rect 2046 3470 2062 3504
rect 1996 3454 2062 3470
rect 2334 3742 2364 3768
rect 2334 3520 2364 3542
rect 2316 3504 2382 3520
rect 2316 3470 2332 3504
rect 2366 3470 2382 3504
rect 2316 3454 2382 3470
rect 2654 3742 2684 3768
rect 2654 3520 2684 3542
rect 2636 3504 2702 3520
rect 2636 3470 2652 3504
rect 2686 3470 2702 3504
rect 2636 3454 2702 3470
rect 2974 3742 3004 3768
rect 2974 3520 3004 3542
rect 2956 3504 3022 3520
rect 2956 3470 2972 3504
rect 3006 3470 3022 3504
rect 2956 3454 3022 3470
<< polycont >>
rect 92 4287 126 4321
rect 412 4287 446 4321
rect 732 4287 766 4321
rect 1052 4287 1086 4321
rect 1372 4287 1406 4321
rect 1692 4287 1726 4321
rect 2012 4287 2046 4321
rect 2332 4287 2366 4321
rect 2652 4287 2686 4321
rect 2972 4287 3006 4321
rect 92 3470 126 3504
rect 412 3470 446 3504
rect 732 3470 766 3504
rect 1052 3470 1086 3504
rect 1372 3470 1406 3504
rect 1692 3470 1726 3504
rect 2012 3470 2046 3504
rect 2332 3470 2366 3504
rect 2652 3470 2686 3504
rect 2972 3470 3006 3504
<< locali >>
rect -142 4452 3218 4472
rect -142 4412 -12 4452
rect 228 4412 308 4452
rect 548 4412 628 4452
rect 868 4412 948 4452
rect 1188 4412 1268 4452
rect 1508 4412 1588 4452
rect 1828 4412 1908 4452
rect 2148 4412 2228 4452
rect 2468 4412 2548 4452
rect 2788 4412 2868 4452
rect 3108 4412 3218 4452
rect -142 4390 30 4412
rect 188 4390 350 4412
rect 508 4390 670 4412
rect 828 4390 990 4412
rect 1148 4390 1310 4412
rect 1468 4390 1630 4412
rect 1788 4390 1950 4412
rect 2108 4390 2270 4412
rect 2428 4390 2590 4412
rect 2748 4390 2910 4412
rect 3068 4390 3218 4412
rect -142 4382 3218 4390
rect 76 4287 92 4321
rect 126 4287 142 4321
rect 396 4287 412 4321
rect 446 4287 462 4321
rect 716 4287 732 4321
rect 766 4287 782 4321
rect 1036 4287 1052 4321
rect 1086 4287 1102 4321
rect 1356 4287 1372 4321
rect 1406 4287 1422 4321
rect 1676 4287 1692 4321
rect 1726 4287 1742 4321
rect 1996 4287 2012 4321
rect 2046 4287 2062 4321
rect 2316 4287 2332 4321
rect 2366 4287 2382 4321
rect 2636 4287 2652 4321
rect 2686 4287 2702 4321
rect 2956 4287 2972 4321
rect 3006 4287 3022 4321
rect 48 4228 82 4244
rect 48 4036 82 4052
rect 136 4228 170 4244
rect 136 4036 170 4052
rect 368 4228 402 4244
rect 368 4036 402 4052
rect 456 4228 490 4244
rect 456 4036 490 4052
rect 688 4228 722 4244
rect 688 4036 722 4052
rect 776 4228 810 4244
rect 776 4036 810 4052
rect 1008 4228 1042 4244
rect 1008 4036 1042 4052
rect 1096 4228 1130 4244
rect 1096 4036 1130 4052
rect 1328 4228 1362 4244
rect 1328 4036 1362 4052
rect 1416 4228 1450 4244
rect 1416 4036 1450 4052
rect 1648 4228 1682 4244
rect 1648 4036 1682 4052
rect 1736 4228 1770 4244
rect 1736 4036 1770 4052
rect 1968 4228 2002 4244
rect 1968 4036 2002 4052
rect 2056 4228 2090 4244
rect 2056 4036 2090 4052
rect 2288 4228 2322 4244
rect 2288 4036 2322 4052
rect 2376 4228 2410 4244
rect 2376 4036 2410 4052
rect 2608 4228 2642 4244
rect 2608 4036 2642 4052
rect 2696 4228 2730 4244
rect 2696 4036 2730 4052
rect 2928 4228 2962 4244
rect 2928 4036 2962 4052
rect 3016 4228 3050 4244
rect 3016 4036 3050 4052
rect 48 3730 82 3746
rect 48 3538 82 3554
rect 136 3730 170 3746
rect 136 3538 170 3554
rect 368 3730 402 3746
rect 368 3538 402 3554
rect 456 3730 490 3746
rect 456 3538 490 3554
rect 688 3730 722 3746
rect 688 3538 722 3554
rect 776 3730 810 3746
rect 776 3538 810 3554
rect 1008 3730 1042 3746
rect 1008 3538 1042 3554
rect 1096 3730 1130 3746
rect 1096 3538 1130 3554
rect 1328 3730 1362 3746
rect 1328 3538 1362 3554
rect 1416 3730 1450 3746
rect 1416 3538 1450 3554
rect 1648 3730 1682 3746
rect 1648 3538 1682 3554
rect 1736 3730 1770 3746
rect 1736 3538 1770 3554
rect 1968 3730 2002 3746
rect 1968 3538 2002 3554
rect 2056 3730 2090 3746
rect 2056 3538 2090 3554
rect 2288 3730 2322 3746
rect 2288 3538 2322 3554
rect 2376 3730 2410 3746
rect 2376 3538 2410 3554
rect 2608 3730 2642 3746
rect 2608 3538 2642 3554
rect 2696 3730 2730 3746
rect 2696 3538 2730 3554
rect 2928 3730 2962 3746
rect 2928 3538 2962 3554
rect 3016 3730 3050 3746
rect 3016 3538 3050 3554
rect 76 3470 92 3504
rect 126 3470 142 3504
rect 396 3470 412 3504
rect 446 3470 462 3504
rect 716 3470 732 3504
rect 766 3470 782 3504
rect 1036 3470 1052 3504
rect 1086 3470 1102 3504
rect 1356 3470 1372 3504
rect 1406 3470 1422 3504
rect 1676 3470 1692 3504
rect 1726 3470 1742 3504
rect 1996 3470 2012 3504
rect 2046 3470 2062 3504
rect 2316 3470 2332 3504
rect 2366 3470 2382 3504
rect 2636 3470 2652 3504
rect 2686 3470 2702 3504
rect 2956 3470 2972 3504
rect 3006 3470 3022 3504
rect -142 3402 3168 3412
rect -142 3382 30 3402
rect 188 3382 350 3402
rect 508 3382 670 3402
rect 828 3382 990 3402
rect 1148 3382 1310 3402
rect 1468 3382 1630 3402
rect 1788 3382 1950 3402
rect 2108 3382 2270 3402
rect 2428 3382 2590 3402
rect 2748 3382 2910 3402
rect 3068 3382 3168 3402
rect -142 3342 -12 3382
rect 228 3342 308 3382
rect 548 3342 628 3382
rect 868 3342 948 3382
rect 1188 3342 1268 3382
rect 1508 3342 1588 3382
rect 1828 3342 1908 3382
rect 2148 3342 2228 3382
rect 2468 3342 2548 3382
rect 2788 3342 2868 3382
rect 3108 3342 3168 3382
rect -142 3322 3168 3342
<< viali >>
rect -12 4424 228 4452
rect -12 4412 30 4424
rect 30 4412 188 4424
rect 188 4412 228 4424
rect 308 4424 548 4452
rect 308 4412 350 4424
rect 350 4412 508 4424
rect 508 4412 548 4424
rect 628 4424 868 4452
rect 628 4412 670 4424
rect 670 4412 828 4424
rect 828 4412 868 4424
rect 948 4424 1188 4452
rect 948 4412 990 4424
rect 990 4412 1148 4424
rect 1148 4412 1188 4424
rect 1268 4424 1508 4452
rect 1268 4412 1310 4424
rect 1310 4412 1468 4424
rect 1468 4412 1508 4424
rect 1588 4424 1828 4452
rect 1588 4412 1630 4424
rect 1630 4412 1788 4424
rect 1788 4412 1828 4424
rect 1908 4424 2148 4452
rect 1908 4412 1950 4424
rect 1950 4412 2108 4424
rect 2108 4412 2148 4424
rect 2228 4424 2468 4452
rect 2228 4412 2270 4424
rect 2270 4412 2428 4424
rect 2428 4412 2468 4424
rect 2548 4424 2788 4452
rect 2548 4412 2590 4424
rect 2590 4412 2748 4424
rect 2748 4412 2788 4424
rect 2868 4424 3108 4452
rect 2868 4412 2910 4424
rect 2910 4412 3068 4424
rect 3068 4412 3108 4424
rect 92 4287 126 4321
rect 412 4287 446 4321
rect 732 4287 766 4321
rect 1052 4287 1086 4321
rect 1372 4287 1406 4321
rect 1692 4287 1726 4321
rect 2012 4287 2046 4321
rect 2332 4287 2366 4321
rect 2652 4287 2686 4321
rect 2972 4287 3006 4321
rect 48 4052 82 4228
rect 136 4052 170 4228
rect 368 4052 402 4228
rect 456 4052 490 4228
rect 688 4052 722 4228
rect 776 4052 810 4228
rect 1008 4052 1042 4228
rect 1096 4052 1130 4228
rect 1328 4052 1362 4228
rect 1416 4052 1450 4228
rect 1648 4052 1682 4228
rect 1736 4052 1770 4228
rect 1968 4052 2002 4228
rect 2056 4052 2090 4228
rect 2288 4052 2322 4228
rect 2376 4052 2410 4228
rect 2608 4052 2642 4228
rect 2696 4052 2730 4228
rect 2928 4052 2962 4228
rect 3016 4052 3050 4228
rect 48 3554 82 3730
rect 136 3554 170 3730
rect 368 3554 402 3730
rect 456 3554 490 3730
rect 688 3554 722 3730
rect 776 3554 810 3730
rect 1008 3554 1042 3730
rect 1096 3554 1130 3730
rect 1328 3554 1362 3730
rect 1416 3554 1450 3730
rect 1648 3554 1682 3730
rect 1736 3554 1770 3730
rect 1968 3554 2002 3730
rect 2056 3554 2090 3730
rect 2288 3554 2322 3730
rect 2376 3554 2410 3730
rect 2608 3554 2642 3730
rect 2696 3554 2730 3730
rect 2928 3554 2962 3730
rect 3016 3554 3050 3730
rect 92 3470 126 3504
rect 412 3470 446 3504
rect 732 3470 766 3504
rect 1052 3470 1086 3504
rect 1372 3470 1406 3504
rect 1692 3470 1726 3504
rect 2012 3470 2046 3504
rect 2332 3470 2366 3504
rect 2652 3470 2686 3504
rect 2972 3470 3006 3504
rect -12 3368 30 3382
rect 30 3368 188 3382
rect 188 3368 228 3382
rect -12 3342 228 3368
rect 308 3368 350 3382
rect 350 3368 508 3382
rect 508 3368 548 3382
rect 308 3342 548 3368
rect 628 3368 670 3382
rect 670 3368 828 3382
rect 828 3368 868 3382
rect 628 3342 868 3368
rect 948 3368 990 3382
rect 990 3368 1148 3382
rect 1148 3368 1188 3382
rect 948 3342 1188 3368
rect 1268 3368 1310 3382
rect 1310 3368 1468 3382
rect 1468 3368 1508 3382
rect 1268 3342 1508 3368
rect 1588 3368 1630 3382
rect 1630 3368 1788 3382
rect 1788 3368 1828 3382
rect 1588 3342 1828 3368
rect 1908 3368 1950 3382
rect 1950 3368 2108 3382
rect 2108 3368 2148 3382
rect 1908 3342 2148 3368
rect 2228 3368 2270 3382
rect 2270 3368 2428 3382
rect 2428 3368 2468 3382
rect 2228 3342 2468 3368
rect 2548 3368 2590 3382
rect 2590 3368 2748 3382
rect 2748 3368 2788 3382
rect 2548 3342 2788 3368
rect 2868 3368 2910 3382
rect 2910 3368 3068 3382
rect 3068 3368 3108 3382
rect 2868 3342 3108 3368
<< metal1 >>
rect -182 4452 3258 4472
rect -182 4412 -12 4452
rect 228 4412 308 4452
rect 548 4412 628 4452
rect 868 4412 948 4452
rect 1188 4412 1268 4452
rect 1508 4412 1588 4452
rect 1828 4412 1908 4452
rect 2148 4412 2228 4452
rect 2468 4412 2548 4452
rect 2788 4412 2868 4452
rect 3108 4412 3258 4452
rect -182 4402 3258 4412
rect 58 4282 78 4342
rect 138 4282 158 4342
rect 378 4282 398 4342
rect 458 4282 478 4342
rect 698 4282 718 4342
rect 778 4282 798 4342
rect 1018 4282 1038 4342
rect 1098 4282 1118 4342
rect 1338 4282 1358 4342
rect 1418 4282 1438 4342
rect 1658 4282 1678 4342
rect 1738 4282 1758 4342
rect 1978 4282 1998 4342
rect 2058 4282 2078 4342
rect 2298 4282 2318 4342
rect 2378 4282 2398 4342
rect 2618 4282 2638 4342
rect 2698 4282 2718 4342
rect 2938 4282 2958 4342
rect 3018 4282 3038 4342
rect 80 4281 138 4282
rect 400 4281 458 4282
rect 720 4281 778 4282
rect 1040 4281 1098 4282
rect 1360 4281 1418 4282
rect 1680 4281 1738 4282
rect 2000 4281 2058 4282
rect 2320 4281 2378 4282
rect 2640 4281 2698 4282
rect 2960 4281 3018 4282
rect 42 4228 88 4240
rect 42 4052 48 4228
rect 82 4052 88 4228
rect 42 4040 88 4052
rect 130 4228 176 4240
rect 130 4052 136 4228
rect 170 4052 176 4228
rect 130 4040 176 4052
rect 362 4228 408 4240
rect 362 4052 368 4228
rect 402 4052 408 4228
rect 362 4040 408 4052
rect 450 4228 496 4240
rect 450 4052 456 4228
rect 490 4052 496 4228
rect 450 4040 496 4052
rect 682 4228 728 4240
rect 682 4052 688 4228
rect 722 4052 728 4228
rect 682 4040 728 4052
rect 770 4228 816 4240
rect 770 4052 776 4228
rect 810 4052 816 4228
rect 770 4040 816 4052
rect 1002 4228 1048 4240
rect 1002 4052 1008 4228
rect 1042 4052 1048 4228
rect 1002 4040 1048 4052
rect 1090 4228 1136 4240
rect 1090 4052 1096 4228
rect 1130 4052 1136 4228
rect 1090 4040 1136 4052
rect 1322 4228 1368 4240
rect 1322 4052 1328 4228
rect 1362 4052 1368 4228
rect 1322 4040 1368 4052
rect 1410 4228 1456 4240
rect 1410 4052 1416 4228
rect 1450 4052 1456 4228
rect 1410 4040 1456 4052
rect 1642 4228 1688 4240
rect 1642 4052 1648 4228
rect 1682 4052 1688 4228
rect 1642 4040 1688 4052
rect 1730 4228 1776 4240
rect 1730 4052 1736 4228
rect 1770 4052 1776 4228
rect 1730 4040 1776 4052
rect 1962 4228 2008 4240
rect 1962 4052 1968 4228
rect 2002 4052 2008 4228
rect 1962 4040 2008 4052
rect 2050 4228 2096 4240
rect 2050 4052 2056 4228
rect 2090 4052 2096 4228
rect 2050 4040 2096 4052
rect 2282 4228 2328 4240
rect 2282 4052 2288 4228
rect 2322 4052 2328 4228
rect 2282 4040 2328 4052
rect 2370 4228 2416 4240
rect 2370 4052 2376 4228
rect 2410 4052 2416 4228
rect 2370 4040 2416 4052
rect 2602 4228 2648 4240
rect 2602 4052 2608 4228
rect 2642 4052 2648 4228
rect 2602 4040 2648 4052
rect 2690 4228 2736 4240
rect 2690 4052 2696 4228
rect 2730 4052 2736 4228
rect 2690 4040 2736 4052
rect 2922 4228 2968 4240
rect 2922 4052 2928 4228
rect 2962 4052 2968 4228
rect 2922 4040 2968 4052
rect 3010 4228 3056 4240
rect 3010 4052 3016 4228
rect 3050 4052 3056 4228
rect 3010 4040 3056 4052
rect 48 3932 78 4040
rect -2 3922 78 3932
rect -2 3862 8 3922
rect 68 3862 78 3922
rect -2 3852 78 3862
rect 48 3742 78 3852
rect 138 3932 168 4040
rect 368 3932 398 4040
rect 138 3920 248 3932
rect 138 3860 180 3920
rect 240 3860 248 3920
rect 138 3852 248 3860
rect 318 3922 398 3932
rect 318 3862 328 3922
rect 388 3862 398 3922
rect 318 3852 398 3862
rect 138 3742 168 3852
rect 368 3742 398 3852
rect 458 3932 488 4040
rect 688 3932 718 4040
rect 458 3852 568 3932
rect 638 3922 718 3932
rect 638 3862 648 3922
rect 708 3862 718 3922
rect 638 3852 718 3862
rect 458 3742 488 3852
rect 688 3742 718 3852
rect 778 3932 808 4040
rect 1008 3932 1038 4040
rect 778 3852 888 3932
rect 958 3922 1038 3932
rect 958 3862 968 3922
rect 1028 3862 1038 3922
rect 958 3852 1038 3862
rect 778 3742 808 3852
rect 1008 3742 1038 3852
rect 1098 3932 1128 4040
rect 1328 3932 1358 4040
rect 1098 3852 1208 3932
rect 1278 3922 1358 3932
rect 1278 3862 1288 3922
rect 1348 3862 1358 3922
rect 1278 3852 1358 3862
rect 1098 3742 1128 3852
rect 1328 3742 1358 3852
rect 1418 3932 1448 4040
rect 1648 3932 1678 4040
rect 1418 3852 1528 3932
rect 1598 3922 1678 3932
rect 1598 3862 1608 3922
rect 1668 3862 1678 3922
rect 1598 3852 1678 3862
rect 1418 3742 1448 3852
rect 1648 3742 1678 3852
rect 1738 3932 1768 4040
rect 1968 3932 1998 4040
rect 1738 3852 1848 3932
rect 1918 3922 1998 3932
rect 1918 3862 1928 3922
rect 1988 3862 1998 3922
rect 1918 3852 1998 3862
rect 1738 3742 1768 3852
rect 1968 3742 1998 3852
rect 2058 3932 2088 4040
rect 2288 3932 2318 4040
rect 2058 3852 2168 3932
rect 2238 3922 2318 3932
rect 2238 3862 2248 3922
rect 2308 3862 2318 3922
rect 2238 3852 2318 3862
rect 2058 3742 2088 3852
rect 2288 3742 2318 3852
rect 2378 3932 2408 4040
rect 2608 3932 2638 4040
rect 2378 3852 2488 3932
rect 2558 3922 2638 3932
rect 2558 3862 2568 3922
rect 2628 3862 2638 3922
rect 2558 3852 2638 3862
rect 2378 3742 2408 3852
rect 2608 3742 2638 3852
rect 2698 3932 2728 4040
rect 2928 3932 2958 4040
rect 2698 3852 2808 3932
rect 2878 3922 2958 3932
rect 2878 3862 2888 3922
rect 2948 3862 2958 3922
rect 2878 3852 2958 3862
rect 2698 3742 2728 3852
rect 2928 3742 2958 3852
rect 3018 3932 3048 4040
rect 3018 3852 3128 3932
rect 3018 3742 3048 3852
rect 42 3730 88 3742
rect 42 3554 48 3730
rect 82 3554 88 3730
rect 42 3542 88 3554
rect 130 3730 176 3742
rect 130 3554 136 3730
rect 170 3554 176 3730
rect 130 3542 176 3554
rect 362 3730 408 3742
rect 362 3554 368 3730
rect 402 3554 408 3730
rect 362 3542 408 3554
rect 450 3730 496 3742
rect 450 3554 456 3730
rect 490 3554 496 3730
rect 450 3542 496 3554
rect 682 3730 728 3742
rect 682 3554 688 3730
rect 722 3554 728 3730
rect 682 3542 728 3554
rect 770 3730 816 3742
rect 770 3554 776 3730
rect 810 3554 816 3730
rect 770 3542 816 3554
rect 1002 3730 1048 3742
rect 1002 3554 1008 3730
rect 1042 3554 1048 3730
rect 1002 3542 1048 3554
rect 1090 3730 1136 3742
rect 1090 3554 1096 3730
rect 1130 3554 1136 3730
rect 1090 3542 1136 3554
rect 1322 3730 1368 3742
rect 1322 3554 1328 3730
rect 1362 3554 1368 3730
rect 1322 3542 1368 3554
rect 1410 3730 1456 3742
rect 1410 3554 1416 3730
rect 1450 3554 1456 3730
rect 1410 3542 1456 3554
rect 1642 3730 1688 3742
rect 1642 3554 1648 3730
rect 1682 3554 1688 3730
rect 1642 3542 1688 3554
rect 1730 3730 1776 3742
rect 1730 3554 1736 3730
rect 1770 3554 1776 3730
rect 1730 3542 1776 3554
rect 1962 3730 2008 3742
rect 1962 3554 1968 3730
rect 2002 3554 2008 3730
rect 1962 3542 2008 3554
rect 2050 3730 2096 3742
rect 2050 3554 2056 3730
rect 2090 3554 2096 3730
rect 2050 3542 2096 3554
rect 2282 3730 2328 3742
rect 2282 3554 2288 3730
rect 2322 3554 2328 3730
rect 2282 3542 2328 3554
rect 2370 3730 2416 3742
rect 2370 3554 2376 3730
rect 2410 3554 2416 3730
rect 2370 3542 2416 3554
rect 2602 3730 2648 3742
rect 2602 3554 2608 3730
rect 2642 3554 2648 3730
rect 2602 3542 2648 3554
rect 2690 3730 2736 3742
rect 2690 3554 2696 3730
rect 2730 3554 2736 3730
rect 2690 3542 2736 3554
rect 2922 3730 2968 3742
rect 2922 3554 2928 3730
rect 2962 3554 2968 3730
rect 2922 3542 2968 3554
rect 3010 3730 3056 3742
rect 3010 3554 3016 3730
rect 3050 3554 3056 3730
rect 3010 3542 3056 3554
rect 58 3442 78 3512
rect 138 3442 158 3512
rect 58 3432 158 3442
rect 378 3442 398 3512
rect 458 3442 478 3512
rect 378 3432 478 3442
rect 698 3442 718 3512
rect 778 3442 798 3512
rect 698 3432 798 3442
rect 1018 3442 1038 3512
rect 1098 3442 1118 3512
rect 1018 3432 1118 3442
rect 1338 3442 1358 3512
rect 1418 3442 1438 3512
rect 1338 3432 1438 3442
rect 1658 3442 1678 3512
rect 1738 3442 1758 3512
rect 1658 3432 1758 3442
rect 1978 3442 1998 3512
rect 2058 3442 2078 3512
rect 1978 3432 2078 3442
rect 2298 3442 2318 3512
rect 2378 3442 2398 3512
rect 2298 3432 2398 3442
rect 2618 3442 2638 3512
rect 2698 3442 2718 3512
rect 2618 3432 2718 3442
rect 2938 3442 2958 3512
rect 3018 3442 3038 3512
rect 2938 3432 3038 3442
rect -182 3382 3208 3392
rect -182 3342 -12 3382
rect 228 3342 308 3382
rect 548 3342 628 3382
rect 868 3342 948 3382
rect 1188 3342 1268 3382
rect 1508 3342 1588 3382
rect 1828 3342 1908 3382
rect 2148 3342 2228 3382
rect 2468 3342 2548 3382
rect 2788 3342 2868 3382
rect 3108 3342 3208 3382
rect -182 3322 3208 3342
rect -142 3232 188 3262
rect 178 3202 188 3232
rect 248 3232 508 3262
rect 248 3202 258 3232
rect 498 3202 508 3232
rect 568 3232 828 3262
rect 568 3202 578 3232
rect 818 3202 828 3232
rect 888 3232 1148 3262
rect 888 3202 898 3232
rect 1138 3202 1148 3232
rect 1208 3232 1468 3262
rect 1208 3202 1218 3232
rect 1458 3202 1468 3232
rect 1528 3232 1788 3262
rect 1528 3202 1538 3232
rect 1778 3202 1788 3232
rect 1848 3232 2108 3262
rect 1848 3202 1858 3232
rect 2098 3202 2108 3232
rect 2168 3232 2428 3262
rect 2168 3202 2178 3232
rect 2418 3202 2428 3232
rect 2488 3232 2748 3262
rect 2488 3202 2498 3232
rect 2738 3202 2748 3232
rect 2808 3232 3068 3262
rect 2808 3202 2818 3232
rect 3058 3202 3068 3232
rect 3128 3232 3208 3262
rect 3128 3202 3138 3232
<< via1 >>
rect 78 4321 138 4342
rect 78 4287 92 4321
rect 92 4287 126 4321
rect 126 4287 138 4321
rect 78 4282 138 4287
rect 398 4321 458 4342
rect 398 4287 412 4321
rect 412 4287 446 4321
rect 446 4287 458 4321
rect 398 4282 458 4287
rect 718 4321 778 4342
rect 718 4287 732 4321
rect 732 4287 766 4321
rect 766 4287 778 4321
rect 718 4282 778 4287
rect 1038 4321 1098 4342
rect 1038 4287 1052 4321
rect 1052 4287 1086 4321
rect 1086 4287 1098 4321
rect 1038 4282 1098 4287
rect 1358 4321 1418 4342
rect 1358 4287 1372 4321
rect 1372 4287 1406 4321
rect 1406 4287 1418 4321
rect 1358 4282 1418 4287
rect 1678 4321 1738 4342
rect 1678 4287 1692 4321
rect 1692 4287 1726 4321
rect 1726 4287 1738 4321
rect 1678 4282 1738 4287
rect 1998 4321 2058 4342
rect 1998 4287 2012 4321
rect 2012 4287 2046 4321
rect 2046 4287 2058 4321
rect 1998 4282 2058 4287
rect 2318 4321 2378 4342
rect 2318 4287 2332 4321
rect 2332 4287 2366 4321
rect 2366 4287 2378 4321
rect 2318 4282 2378 4287
rect 2638 4321 2698 4342
rect 2638 4287 2652 4321
rect 2652 4287 2686 4321
rect 2686 4287 2698 4321
rect 2638 4282 2698 4287
rect 2958 4321 3018 4342
rect 2958 4287 2972 4321
rect 2972 4287 3006 4321
rect 3006 4287 3018 4321
rect 2958 4282 3018 4287
rect 8 3862 68 3922
rect 180 3860 240 3920
rect 328 3862 388 3922
rect 648 3862 708 3922
rect 968 3862 1028 3922
rect 1288 3862 1348 3922
rect 1608 3862 1668 3922
rect 1928 3862 1988 3922
rect 2248 3862 2308 3922
rect 2568 3862 2628 3922
rect 2888 3862 2948 3922
rect 78 3504 138 3512
rect 78 3470 92 3504
rect 92 3470 126 3504
rect 126 3470 138 3504
rect 78 3442 138 3470
rect 398 3504 458 3512
rect 398 3470 412 3504
rect 412 3470 446 3504
rect 446 3470 458 3504
rect 398 3442 458 3470
rect 718 3504 778 3512
rect 718 3470 732 3504
rect 732 3470 766 3504
rect 766 3470 778 3504
rect 718 3442 778 3470
rect 1038 3504 1098 3512
rect 1038 3470 1052 3504
rect 1052 3470 1086 3504
rect 1086 3470 1098 3504
rect 1038 3442 1098 3470
rect 1358 3504 1418 3512
rect 1358 3470 1372 3504
rect 1372 3470 1406 3504
rect 1406 3470 1418 3504
rect 1358 3442 1418 3470
rect 1678 3504 1738 3512
rect 1678 3470 1692 3504
rect 1692 3470 1726 3504
rect 1726 3470 1738 3504
rect 1678 3442 1738 3470
rect 1998 3504 2058 3512
rect 1998 3470 2012 3504
rect 2012 3470 2046 3504
rect 2046 3470 2058 3504
rect 1998 3442 2058 3470
rect 2318 3504 2378 3512
rect 2318 3470 2332 3504
rect 2332 3470 2366 3504
rect 2366 3470 2378 3504
rect 2318 3442 2378 3470
rect 2638 3504 2698 3512
rect 2638 3470 2652 3504
rect 2652 3470 2686 3504
rect 2686 3470 2698 3504
rect 2638 3442 2698 3470
rect 2958 3504 3018 3512
rect 2958 3470 2972 3504
rect 2972 3470 3006 3504
rect 3006 3470 3018 3504
rect 2958 3442 3018 3470
rect 188 3202 248 3262
rect 508 3202 568 3262
rect 828 3202 888 3262
rect 1148 3202 1208 3262
rect 1468 3202 1528 3262
rect 1788 3202 1848 3262
rect 2108 3202 2168 3262
rect 2428 3202 2488 3262
rect 2748 3202 2808 3262
rect 3068 3202 3128 3262
<< metal2 >>
rect -142 4502 3188 4532
rect -2 3932 28 4502
rect 68 4282 78 4342
rect 138 4282 148 4342
rect -2 3922 78 3932
rect -2 3862 8 3922
rect 68 3862 78 3922
rect -2 3852 78 3862
rect 108 3572 138 4282
rect 318 3932 348 4502
rect 388 4282 398 4342
rect 458 4282 468 4342
rect 168 3922 248 3932
rect 168 3862 178 3922
rect 238 3920 248 3922
rect 168 3860 180 3862
rect 240 3860 248 3920
rect 168 3852 248 3860
rect 318 3922 398 3932
rect 318 3862 328 3922
rect 388 3862 398 3922
rect 318 3852 398 3862
rect 428 3572 458 4282
rect 638 3932 668 4502
rect 708 4282 718 4342
rect 778 4282 788 4342
rect 488 3922 568 3932
rect 488 3862 498 3922
rect 558 3862 568 3922
rect 488 3852 568 3862
rect 638 3922 718 3932
rect 638 3862 648 3922
rect 708 3862 718 3922
rect 638 3852 718 3862
rect 748 3572 778 4282
rect 958 3932 988 4502
rect 1028 4282 1038 4342
rect 1098 4282 1108 4342
rect 808 3922 888 3932
rect 808 3862 818 3922
rect 878 3862 888 3922
rect 808 3852 888 3862
rect 958 3922 1038 3932
rect 958 3862 968 3922
rect 1028 3862 1038 3922
rect 958 3852 1038 3862
rect 1068 3572 1098 4282
rect 1278 3932 1308 4502
rect 1348 4282 1358 4342
rect 1418 4282 1428 4342
rect 1128 3922 1208 3932
rect 1128 3862 1138 3922
rect 1198 3862 1208 3922
rect 1128 3852 1208 3862
rect 1278 3922 1358 3932
rect 1278 3862 1288 3922
rect 1348 3862 1358 3922
rect 1278 3852 1358 3862
rect 1388 3572 1418 4282
rect 1598 3932 1628 4502
rect 1668 4282 1678 4342
rect 1738 4282 1748 4342
rect 1448 3922 1528 3932
rect 1448 3862 1458 3922
rect 1518 3862 1528 3922
rect 1448 3852 1528 3862
rect 1598 3922 1678 3932
rect 1598 3862 1608 3922
rect 1668 3862 1678 3922
rect 1598 3852 1678 3862
rect 1708 3572 1738 4282
rect 1918 3932 1948 4502
rect 1988 4282 1998 4342
rect 2058 4282 2068 4342
rect 1768 3922 1848 3932
rect 1768 3862 1778 3922
rect 1838 3862 1848 3922
rect 1768 3852 1848 3862
rect 1918 3922 1998 3932
rect 1918 3862 1928 3922
rect 1988 3862 1998 3922
rect 1918 3852 1998 3862
rect 2028 3572 2058 4282
rect 2238 3932 2268 4502
rect 2308 4282 2318 4342
rect 2378 4282 2388 4342
rect 2088 3922 2168 3932
rect 2088 3862 2098 3922
rect 2158 3862 2168 3922
rect 2088 3852 2168 3862
rect 2238 3922 2318 3932
rect 2238 3862 2248 3922
rect 2308 3862 2318 3922
rect 2238 3852 2318 3862
rect 2348 3572 2378 4282
rect 2558 3932 2588 4502
rect 2628 4282 2638 4342
rect 2698 4282 2708 4342
rect 2408 3922 2488 3932
rect 2408 3862 2418 3922
rect 2478 3862 2488 3922
rect 2408 3852 2488 3862
rect 2558 3922 2638 3932
rect 2558 3862 2568 3922
rect 2628 3862 2638 3922
rect 2558 3852 2638 3862
rect 2668 3572 2698 4282
rect 2878 3932 2908 4502
rect 2948 4282 2958 4342
rect 3018 4282 3028 4342
rect 2728 3922 2808 3932
rect 2728 3862 2738 3922
rect 2798 3862 2808 3922
rect 2728 3852 2808 3862
rect 2878 3922 2958 3932
rect 2878 3862 2888 3922
rect 2948 3862 2958 3922
rect 2878 3852 2958 3862
rect 2988 3572 3018 4282
rect 3048 3922 3128 3932
rect 3048 3862 3058 3922
rect 3118 3862 3128 3922
rect 3048 3852 3128 3862
rect 108 3542 208 3572
rect 428 3542 528 3572
rect 748 3542 848 3572
rect 1068 3542 1168 3572
rect 1388 3542 1488 3572
rect 1708 3542 1808 3572
rect 2028 3542 2128 3572
rect 2348 3542 2448 3572
rect 2668 3542 2768 3572
rect 2988 3542 3088 3572
rect 68 3442 78 3512
rect 138 3442 148 3512
rect 68 3432 148 3442
rect 98 3262 128 3432
rect 48 3252 128 3262
rect 48 3192 58 3252
rect 118 3192 128 3252
rect 178 3262 208 3542
rect 388 3442 398 3512
rect 458 3442 468 3512
rect 388 3432 468 3442
rect 418 3262 448 3432
rect 178 3202 188 3262
rect 248 3202 258 3262
rect 368 3252 448 3262
rect 48 3182 128 3192
rect 368 3192 378 3252
rect 438 3192 448 3252
rect 498 3262 528 3542
rect 708 3442 718 3512
rect 778 3442 788 3512
rect 708 3432 788 3442
rect 738 3262 768 3432
rect 498 3202 508 3262
rect 568 3202 578 3262
rect 688 3252 768 3262
rect 368 3182 448 3192
rect 688 3192 698 3252
rect 758 3192 768 3252
rect 818 3262 848 3542
rect 1028 3442 1038 3512
rect 1098 3442 1108 3512
rect 1028 3432 1108 3442
rect 1058 3262 1088 3432
rect 818 3202 828 3262
rect 888 3202 898 3262
rect 1008 3252 1088 3262
rect 688 3182 768 3192
rect 1008 3192 1018 3252
rect 1078 3192 1088 3252
rect 1138 3262 1168 3542
rect 1348 3442 1358 3512
rect 1418 3442 1428 3512
rect 1348 3432 1428 3442
rect 1378 3262 1408 3432
rect 1138 3202 1148 3262
rect 1208 3202 1218 3262
rect 1328 3252 1408 3262
rect 1008 3182 1088 3192
rect 1328 3192 1338 3252
rect 1398 3192 1408 3252
rect 1458 3262 1488 3542
rect 1668 3442 1678 3512
rect 1738 3442 1748 3512
rect 1668 3432 1748 3442
rect 1698 3262 1728 3432
rect 1458 3202 1468 3262
rect 1528 3202 1538 3262
rect 1648 3252 1728 3262
rect 1328 3182 1408 3192
rect 1648 3192 1658 3252
rect 1718 3192 1728 3252
rect 1778 3262 1808 3542
rect 1988 3442 1998 3512
rect 2058 3442 2068 3512
rect 1988 3432 2068 3442
rect 2018 3262 2048 3432
rect 1778 3202 1788 3262
rect 1848 3202 1858 3262
rect 1968 3252 2048 3262
rect 1648 3182 1728 3192
rect 1968 3192 1978 3252
rect 2038 3192 2048 3252
rect 2098 3262 2128 3542
rect 2308 3442 2318 3512
rect 2378 3442 2388 3512
rect 2308 3432 2388 3442
rect 2338 3262 2368 3432
rect 2098 3202 2108 3262
rect 2168 3202 2178 3262
rect 2288 3252 2368 3262
rect 1968 3182 2048 3192
rect 2288 3192 2298 3252
rect 2358 3192 2368 3252
rect 2418 3262 2448 3542
rect 2628 3442 2638 3512
rect 2698 3442 2708 3512
rect 2628 3432 2708 3442
rect 2658 3262 2688 3432
rect 2418 3202 2428 3262
rect 2488 3202 2498 3262
rect 2608 3252 2688 3262
rect 2288 3182 2368 3192
rect 2608 3192 2618 3252
rect 2678 3192 2688 3252
rect 2738 3262 2768 3542
rect 2948 3442 2958 3512
rect 3018 3442 3028 3512
rect 2948 3432 3028 3442
rect 2978 3262 3008 3432
rect 2738 3202 2748 3262
rect 2808 3202 2818 3262
rect 2928 3252 3008 3262
rect 2608 3182 2688 3192
rect 2928 3192 2938 3252
rect 2998 3192 3008 3252
rect 3058 3262 3088 3542
rect 3058 3202 3068 3262
rect 3128 3202 3138 3262
rect 2928 3182 3008 3192
<< via2 >>
rect 178 3920 238 3922
rect 178 3862 180 3920
rect 180 3862 238 3920
rect 498 3862 558 3922
rect 818 3862 878 3922
rect 1138 3862 1198 3922
rect 1458 3862 1518 3922
rect 1778 3862 1838 3922
rect 2098 3862 2158 3922
rect 2418 3862 2478 3922
rect 2738 3862 2798 3922
rect 3058 3862 3118 3922
rect 58 3192 118 3252
rect 378 3192 438 3252
rect 698 3192 758 3252
rect 1018 3192 1078 3252
rect 1338 3192 1398 3252
rect 1658 3192 1718 3252
rect 1978 3192 2038 3252
rect 2298 3192 2358 3252
rect 2618 3192 2678 3252
rect 2938 3192 2998 3252
<< metal3 >>
rect 168 3932 288 3942
rect 168 3862 178 3932
rect 248 3862 288 3932
rect 168 3852 288 3862
rect 488 3932 608 3942
rect 488 3862 498 3932
rect 568 3862 608 3932
rect 488 3852 608 3862
rect 808 3932 928 3942
rect 808 3862 818 3932
rect 888 3862 928 3932
rect 808 3852 928 3862
rect 1128 3932 1248 3942
rect 1128 3862 1138 3932
rect 1208 3862 1248 3932
rect 1128 3852 1248 3862
rect 1448 3932 1568 3942
rect 1448 3862 1458 3932
rect 1528 3862 1568 3932
rect 1448 3852 1568 3862
rect 1768 3932 1888 3942
rect 1768 3862 1778 3932
rect 1848 3862 1888 3932
rect 1768 3852 1888 3862
rect 2088 3932 2208 3942
rect 2088 3862 2098 3932
rect 2168 3862 2208 3932
rect 2088 3852 2208 3862
rect 2408 3932 2528 3942
rect 2408 3862 2418 3932
rect 2488 3862 2528 3932
rect 2408 3852 2528 3862
rect 2728 3932 2848 3942
rect 2728 3862 2738 3932
rect 2808 3862 2848 3932
rect 2728 3852 2848 3862
rect 3048 3932 3168 3942
rect 3048 3862 3058 3932
rect 3128 3862 3168 3932
rect 3048 3852 3168 3862
rect -142 3252 3208 3262
rect -142 3202 58 3252
rect 48 3192 58 3202
rect 118 3202 378 3252
rect 118 3192 128 3202
rect 48 3182 128 3192
rect 368 3192 378 3202
rect 438 3202 698 3252
rect 438 3192 448 3202
rect 368 3182 448 3192
rect 688 3192 698 3202
rect 758 3202 1018 3252
rect 758 3192 768 3202
rect 688 3182 768 3192
rect 1008 3192 1018 3202
rect 1078 3202 1338 3252
rect 1078 3192 1088 3202
rect 1008 3182 1088 3192
rect 1328 3192 1338 3202
rect 1398 3202 1658 3252
rect 1398 3192 1408 3202
rect 1328 3182 1408 3192
rect 1648 3192 1658 3202
rect 1718 3202 1978 3252
rect 1718 3192 1728 3202
rect 1648 3182 1728 3192
rect 1968 3192 1978 3202
rect 2038 3202 2298 3252
rect 2038 3192 2048 3202
rect 1968 3182 2048 3192
rect 2288 3192 2298 3202
rect 2358 3202 2618 3252
rect 2358 3192 2368 3202
rect 2288 3182 2368 3192
rect 2608 3192 2618 3202
rect 2678 3202 2938 3252
rect 2678 3192 2688 3202
rect 2608 3182 2688 3192
rect 2928 3192 2938 3202
rect 2998 3232 3208 3252
rect 2998 3202 3198 3232
rect 2998 3192 3008 3202
rect 2928 3182 3008 3192
<< via3 >>
rect 178 3922 248 3932
rect 178 3862 238 3922
rect 238 3862 248 3922
rect 498 3922 568 3932
rect 498 3862 558 3922
rect 558 3862 568 3922
rect 818 3922 888 3932
rect 818 3862 878 3922
rect 878 3862 888 3922
rect 1138 3922 1208 3932
rect 1138 3862 1198 3922
rect 1198 3862 1208 3922
rect 1458 3922 1528 3932
rect 1458 3862 1518 3922
rect 1518 3862 1528 3922
rect 1778 3922 1848 3932
rect 1778 3862 1838 3922
rect 1838 3862 1848 3922
rect 2098 3922 2168 3932
rect 2098 3862 2158 3922
rect 2158 3862 2168 3922
rect 2418 3922 2488 3932
rect 2418 3862 2478 3922
rect 2478 3862 2488 3922
rect 2738 3922 2808 3932
rect 2738 3862 2798 3922
rect 2798 3862 2808 3922
rect 3058 3922 3128 3932
rect 3058 3862 3118 3922
rect 3118 3862 3128 3922
<< metal4 >>
rect 168 3932 288 3942
rect 488 3932 608 3942
rect 808 3932 928 3942
rect 1128 3932 1248 3942
rect 1448 3932 1568 3942
rect 1768 3932 1888 3942
rect 2088 3932 2208 3942
rect 2408 3932 2528 3942
rect 2728 3932 2848 3942
rect 3048 3932 3168 3942
rect 168 3862 178 3932
rect 248 3872 498 3932
rect 248 3862 288 3872
rect 168 3852 288 3862
rect 488 3862 498 3872
rect 568 3872 818 3932
rect 568 3862 608 3872
rect 488 3852 608 3862
rect 808 3862 818 3872
rect 888 3872 1138 3932
rect 888 3862 928 3872
rect 808 3852 928 3862
rect 1128 3862 1138 3872
rect 1208 3872 1458 3932
rect 1208 3862 1248 3872
rect 1128 3852 1248 3862
rect 1448 3862 1458 3872
rect 1528 3872 1778 3932
rect 1528 3862 1568 3872
rect 1448 3852 1568 3862
rect 1768 3862 1778 3872
rect 1848 3872 2098 3932
rect 1848 3862 1888 3872
rect 1768 3852 1888 3862
rect 2088 3862 2098 3872
rect 2168 3872 2418 3932
rect 2168 3862 2208 3872
rect 2088 3852 2208 3862
rect 2408 3862 2418 3872
rect 2488 3872 2738 3932
rect 2488 3862 2528 3872
rect 2408 3852 2528 3862
rect 2728 3862 2738 3872
rect 2808 3872 3058 3932
rect 2808 3862 2848 3872
rect 2728 3852 2848 3862
rect 3048 3862 3058 3872
rect 3128 3872 3258 3932
rect 3128 3862 3168 3872
rect 3048 3852 3168 3862
<< labels >>
flabel metal1 -82 4402 -22 4462 0 FreeSans 256 0 0 0 Vdd
port 3 nsew
flabel metal1 10 3864 70 3924 0 FreeSans 256 0 0 0 Vin
port 5 nsew
flabel metal1 -82 3332 -22 3392 0 FreeSans 256 0 0 0 sub
port 6 nsew
rlabel metal1 58 3432 68 3512 1 clk
port 7 n
rlabel metal1 148 4282 158 4342 1 clk_b
port 8 n
rlabel metal1 138 3862 168 3892 1 Vout
port 9 n
flabel metal1 238 4402 298 4462 0 FreeSans 256 0 0 0 Vdd
port 3 nsew
flabel metal1 330 3864 390 3924 0 FreeSans 256 0 0 0 Vin
port 5 nsew
flabel metal1 238 3332 298 3392 0 FreeSans 256 0 0 0 sub
port 6 nsew
rlabel metal1 378 3432 388 3512 1 clk
port 7 n
rlabel metal1 468 4282 478 4342 1 clk_b
port 8 n
rlabel metal1 458 3862 488 3892 1 Vout
port 9 n
flabel metal1 558 4402 618 4462 0 FreeSans 256 0 0 0 Vdd
port 3 nsew
flabel metal1 650 3864 710 3924 0 FreeSans 256 0 0 0 Vin
port 5 nsew
flabel metal1 558 3332 618 3392 0 FreeSans 256 0 0 0 sub
port 6 nsew
rlabel metal1 698 3432 708 3512 1 clk
port 7 n
rlabel metal1 788 4282 798 4342 1 clk_b
port 8 n
rlabel metal1 778 3862 808 3892 1 Vout
port 9 n
flabel metal1 878 4402 938 4462 0 FreeSans 256 0 0 0 Vdd
port 3 nsew
flabel metal1 970 3864 1030 3924 0 FreeSans 256 0 0 0 Vin
port 5 nsew
flabel metal1 878 3332 938 3392 0 FreeSans 256 0 0 0 sub
port 6 nsew
rlabel metal1 1018 3432 1028 3512 1 clk
port 7 n
rlabel metal1 1108 4282 1118 4342 1 clk_b
port 8 n
rlabel metal1 1098 3862 1128 3892 1 Vout
port 9 n
flabel metal1 1198 4402 1258 4462 0 FreeSans 256 0 0 0 Vdd
port 3 nsew
flabel metal1 1290 3864 1350 3924 0 FreeSans 256 0 0 0 Vin
port 5 nsew
flabel metal1 1198 3332 1258 3392 0 FreeSans 256 0 0 0 sub
port 6 nsew
rlabel metal1 1338 3432 1348 3512 1 clk
port 7 n
rlabel metal1 1428 4282 1438 4342 1 clk_b
port 8 n
rlabel metal1 1418 3862 1448 3892 1 Vout
port 9 n
flabel metal1 1838 4402 1898 4462 0 FreeSans 256 0 0 0 Vdd
port 3 nsew
flabel metal1 1930 3864 1990 3924 0 FreeSans 256 0 0 0 Vin
port 5 nsew
flabel metal1 1838 3332 1898 3392 0 FreeSans 256 0 0 0 sub
port 6 nsew
rlabel metal1 1978 3432 1988 3512 1 clk
port 7 n
rlabel metal1 2068 4282 2078 4342 1 clk_b
port 8 n
rlabel metal1 2058 3862 2088 3892 1 Vout
port 9 n
flabel metal1 1518 4402 1578 4462 0 FreeSans 256 0 0 0 Vdd
port 3 nsew
flabel metal1 1610 3864 1670 3924 0 FreeSans 256 0 0 0 Vin
port 5 nsew
flabel metal1 1518 3332 1578 3392 0 FreeSans 256 0 0 0 sub
port 6 nsew
rlabel metal1 1658 3432 1668 3512 1 clk
port 7 n
rlabel metal1 1748 4282 1758 4342 1 clk_b
port 8 n
rlabel metal1 1738 3862 1768 3892 1 Vout
port 9 n
flabel metal1 2158 4402 2218 4462 0 FreeSans 256 0 0 0 Vdd
port 3 nsew
flabel metal1 2250 3864 2310 3924 0 FreeSans 256 0 0 0 Vin
port 5 nsew
flabel metal1 2158 3332 2218 3392 0 FreeSans 256 0 0 0 sub
port 6 nsew
rlabel metal1 2298 3432 2308 3512 1 clk
port 7 n
rlabel metal1 2388 4282 2398 4342 1 clk_b
port 8 n
rlabel metal1 2378 3862 2408 3892 1 Vout
port 9 n
flabel metal1 2478 4402 2538 4462 0 FreeSans 256 0 0 0 Vdd
port 3 nsew
flabel metal1 2570 3864 2630 3924 0 FreeSans 256 0 0 0 Vin
port 5 nsew
flabel metal1 2478 3332 2538 3392 0 FreeSans 256 0 0 0 sub
port 6 nsew
rlabel metal1 2618 3432 2628 3512 1 clk
port 7 n
rlabel metal1 2708 4282 2718 4342 1 clk_b
port 8 n
rlabel metal1 2698 3862 2728 3892 1 Vout
port 9 n
flabel metal1 2798 4402 2858 4462 0 FreeSans 256 0 0 0 Vdd
port 3 nsew
flabel metal1 2890 3864 2950 3924 0 FreeSans 256 0 0 0 Vin
port 5 nsew
flabel metal1 2798 3332 2858 3392 0 FreeSans 256 0 0 0 sub
port 6 nsew
rlabel metal1 2938 3432 2948 3512 1 clk
port 7 n
rlabel metal1 3028 4282 3038 4342 1 clk_b
port 8 n
rlabel metal1 3018 3862 3048 3892 1 Vout
port 9 n
<< end >>
