magic
tech sky130A
magscale 1 2
timestamp 1728662986
<< pwell >>
rect 1326 -1043 1408 -1037
rect 1326 -1111 1408 -1049
<< locali >>
rect 1029 -56 1737 -34
rect 1029 -91 1183 -56
rect 1559 -91 1737 -56
rect 1029 -178 1737 -91
rect 1029 -422 1240 -178
rect 1505 -425 1737 -178
rect 1029 -1139 1241 -931
rect 1501 -1139 1742 -929
rect 1029 -1216 1742 -1139
rect 1029 -1252 1155 -1216
rect 1561 -1252 1742 -1216
rect 1029 -1276 1742 -1252
<< viali >>
rect 1183 -91 1559 -56
rect 1155 -1252 1561 -1216
<< metal1 >>
rect 1278 81 1478 222
rect 1278 28 1338 81
rect 1400 28 1478 81
rect 1278 22 1478 28
rect 978 -46 1178 -44
rect 978 -56 1682 -46
rect 978 -91 1183 -56
rect 1559 -91 1682 -56
rect 978 -107 1682 -91
rect 978 -244 1178 -107
rect 1327 -219 1411 -213
rect 1327 -272 1336 -219
rect 1402 -272 1411 -219
rect 1327 -282 1411 -272
rect 1300 -569 1345 -504
rect 1145 -769 1345 -569
rect 1387 -570 1432 -504
rect 1300 -830 1345 -769
rect 1386 -770 1586 -570
rect 1387 -830 1432 -770
rect 1328 -1049 1407 -1045
rect 977 -1208 1177 -1054
rect 1328 -1102 1335 -1049
rect 1401 -1102 1407 -1049
rect 1328 -1103 1407 -1102
rect 977 -1216 1666 -1208
rect 977 -1252 1155 -1216
rect 1561 -1252 1666 -1216
rect 977 -1254 1666 -1252
rect 1142 -1258 1666 -1254
rect 1280 -1324 1480 -1316
rect 1280 -1381 1335 -1324
rect 1398 -1381 1480 -1324
rect 1280 -1516 1480 -1381
<< via1 >>
rect 1338 28 1400 81
rect 1336 -272 1402 -219
rect 1335 -1102 1401 -1049
rect 1335 -1381 1398 -1324
<< metal2 >>
rect 1328 81 1408 87
rect 1328 28 1338 81
rect 1400 28 1408 81
rect 1328 22 1408 28
rect 1332 -216 1404 22
rect 1329 -219 1409 -216
rect 1329 -272 1336 -219
rect 1402 -272 1409 -219
rect 1329 -279 1409 -272
rect 1324 -1049 1410 -1042
rect 1324 -1102 1335 -1049
rect 1401 -1102 1410 -1049
rect 1324 -1108 1410 -1102
rect 1330 -1324 1402 -1108
rect 1330 -1381 1335 -1324
rect 1398 -1381 1402 -1324
rect 1330 -1407 1402 -1381
use sky130_fd_pr__pfet_01v8_NKK3FE  XM1 ~/saf
timestamp 1728654492
transform 1 0 1369 0 1 -380
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_5WP7M2  XM2 ~/saf
timestamp 1728654492
transform -1 0 1366 0 1 -948
box -211 -279 211 279
<< labels >>
flabel metal1 978 -244 1178 -44 0 FreeSans 256 0 0 0 vdd
port 4 nsew
flabel metal1 1145 -769 1345 -569 0 FreeSans 256 0 0 0 vin
port 3 nsew
flabel metal1 1386 -770 1586 -570 0 FreeSans 256 0 0 0 vout
port 2 nsew
flabel metal1 1280 -1516 1480 -1316 0 FreeSans 256 0 0 0 clk
port 0 nsew
flabel metal1 1278 22 1478 222 0 FreeSans 256 0 0 0 clk_b
port 5 nsew
flabel metal1 977 -1254 1177 -1054 0 FreeSans 256 0 0 0 sub
port 1 nsew
<< end >>
