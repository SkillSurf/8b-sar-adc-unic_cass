magic
tech sky130A
magscale 1 2
timestamp 1730665161
<< pwell >>
rect 1140 -930 1160 -890
rect 1520 -950 1980 -880
<< locali >>
rect 710 180 1520 200
rect 710 140 840 180
rect 1080 140 1160 180
rect 1400 140 1520 180
rect 710 110 1520 140
rect 710 -890 1520 -860
rect 710 -930 840 -890
rect 1080 -930 1140 -890
rect 1400 -930 1520 -890
rect 710 -950 1520 -930
<< viali >>
rect 840 140 1080 180
rect 1160 140 1400 180
rect 840 -930 1080 -890
rect 1140 -930 1400 -890
<< metal1 >>
rect 270 1100 1980 1130
rect 270 980 1980 1010
rect 270 860 1980 890
rect 270 740 1980 770
rect 270 620 1980 650
rect 270 500 1980 530
rect 270 380 1980 410
rect 270 320 1980 350
rect 800 260 810 290
rect 270 230 810 260
rect 870 260 880 290
rect 950 260 960 290
rect 870 230 960 260
rect 1020 260 1030 290
rect 1210 260 1220 290
rect 1020 230 1220 260
rect 1280 260 1290 290
rect 1350 260 1360 290
rect 1280 230 1360 260
rect 1420 260 1430 290
rect 1420 230 1980 260
rect 270 140 750 200
rect 810 180 1430 200
rect 810 140 840 180
rect 1080 140 1160 180
rect 1400 140 1430 180
rect 1490 140 1980 200
rect 270 130 1980 140
rect 910 70 1010 80
rect 910 10 930 70
rect 990 10 1010 70
rect 910 0 1010 10
rect 1220 70 1320 80
rect 1220 10 1240 70
rect 1300 10 1320 70
rect 1220 0 1320 10
rect 900 -340 930 -220
rect 850 -350 930 -340
rect 850 -410 860 -350
rect 920 -410 930 -350
rect 850 -420 930 -410
rect 900 -540 930 -420
rect 990 -340 1020 -220
rect 1210 -340 1240 -220
rect 990 -350 1240 -340
rect 990 -410 1030 -350
rect 1090 -410 1140 -350
rect 1200 -410 1240 -350
rect 990 -420 1240 -410
rect 990 -540 1020 -420
rect 1210 -540 1240 -420
rect 1300 -340 1330 -220
rect 1300 -350 1380 -340
rect 1300 -410 1310 -350
rect 1370 -410 1380 -350
rect 1300 -420 1380 -410
rect 1300 -540 1330 -420
rect 910 -770 1010 -760
rect 910 -830 930 -770
rect 990 -830 1010 -770
rect 910 -840 1010 -830
rect 1220 -770 1320 -760
rect 1220 -830 1240 -770
rect 1300 -830 1320 -770
rect 1220 -840 1320 -830
rect 270 -890 1980 -880
rect 270 -930 840 -890
rect 1080 -930 1140 -890
rect 1400 -930 1980 -890
rect 270 -950 1980 -930
rect 270 -1010 1980 -980
rect 270 -1130 1980 -1100
rect 270 -1250 1980 -1220
rect 270 -1370 1980 -1340
rect 270 -1490 1980 -1460
rect 270 -1610 1980 -1580
rect 270 -1730 1980 -1700
<< via1 >>
rect 810 230 870 290
rect 960 230 1020 290
rect 1220 230 1280 290
rect 1360 230 1420 290
rect 750 140 810 200
rect 1430 140 1490 200
rect 930 10 990 70
rect 1240 10 1300 70
rect 860 -410 920 -350
rect 1030 -410 1090 -350
rect 1140 -410 1200 -350
rect 1310 -410 1370 -350
rect 930 -830 990 -770
rect 1240 -830 1300 -770
<< metal2 >>
rect 270 1100 1980 1130
rect 270 980 1980 1010
rect 270 860 1980 890
rect 270 740 1980 770
rect 270 620 1980 650
rect 270 500 1980 530
rect 270 380 1980 410
rect 800 230 810 290
rect 870 230 880 290
rect 740 140 750 200
rect 810 140 820 200
rect 790 -920 820 140
rect 850 -340 880 230
rect 950 230 960 290
rect 1020 230 1030 290
rect 1210 230 1220 290
rect 1280 230 1290 290
rect 950 80 980 230
rect 1260 80 1290 230
rect 1350 230 1360 290
rect 1420 230 1430 290
rect 920 70 1000 80
rect 920 10 930 70
rect 990 10 1000 70
rect 920 0 1000 10
rect 1230 70 1310 80
rect 1230 10 1240 70
rect 1300 10 1310 70
rect 1230 0 1310 10
rect 1010 -340 1220 -330
rect 1350 -340 1380 230
rect 850 -350 930 -340
rect 850 -410 860 -350
rect 920 -410 930 -350
rect 850 -420 930 -410
rect 1010 -410 1030 -340
rect 1100 -410 1140 -340
rect 1210 -410 1220 -340
rect 1010 -430 1220 -410
rect 1300 -350 1380 -340
rect 1300 -410 1310 -350
rect 1370 -410 1380 -350
rect 1300 -420 1380 -410
rect 1420 140 1430 200
rect 1490 140 1500 200
rect 920 -770 1000 -760
rect 920 -830 930 -770
rect 990 -830 1000 -770
rect 920 -840 1000 -830
rect 1230 -770 1310 -760
rect 1230 -830 1240 -770
rect 1300 -830 1310 -770
rect 1230 -840 1310 -830
rect 950 -920 980 -840
rect 790 -950 980 -920
rect 1260 -920 1290 -840
rect 1420 -920 1450 140
rect 1260 -950 1450 -920
rect 270 -1010 1980 -980
rect 270 -1130 1980 -1100
rect 270 -1250 1980 -1220
rect 270 -1370 1980 -1340
rect 270 -1490 1980 -1460
rect 270 -1610 1980 -1580
rect 270 -1730 1980 -1700
<< via2 >>
rect 1030 -350 1100 -340
rect 1030 -410 1090 -350
rect 1090 -410 1100 -350
rect 1140 -350 1210 -340
rect 1140 -410 1200 -350
rect 1200 -410 1210 -350
<< metal3 >>
rect 990 -340 1240 -310
rect 990 -420 1030 -340
rect 1100 -420 1140 -340
rect 1210 -420 1240 -340
rect 990 -450 1240 -420
rect 380 -1830 440 -1820
<< via3 >>
rect 1030 -410 1100 -340
rect 1030 -420 1100 -410
rect 1140 -410 1210 -340
rect 1140 -420 1210 -410
<< metal4 >>
rect 990 -340 1240 -310
rect 990 -420 1030 -340
rect 1100 -420 1140 -340
rect 1210 -420 1240 -340
rect 990 -450 1240 -420
rect 460 -1920 520 -1840
rect 1090 -1900 1150 -450
rect 380 -2250 510 -2190
rect 480 -3490 550 -3420
use sky130_fd_pr__cap_mim_m3_1_BZXSER  sky130_fd_pr__cap_mim_m3_1_BZXSER_0
timestamp 1728835232
transform 0 1 1120 1 0 -2704
box -886 -740 886 740
use sky130_fd_pr__nfet_01v8_5WU4M2  sky130_fd_pr__nfet_01v8_5WU4M2_0 ~/final
timestamp 1728804544
transform -1 0 1271 0 -1 -661
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_QKK3FL  sky130_fd_pr__pfet_01v8_QKK3FL_0 ~/final
timestamp 1728804544
transform -1 0 1271 0 -1 -96
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_NKK3FE  XM1 ~/final
timestamp 1728804544
transform 1 0 961 0 1 -96
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_5WP7M2  XM2 ~/final
timestamp 1730665161
transform 1 0 961 0 1 -661
box -211 -279 211 279
<< labels >>
flabel via1 860 -410 900 -360 0 FreeSans 320 0 0 0 Vin
flabel metal2 920 -830 980 -780 0 FreeSans 320 0 0 0 phi1
flabel metal1 1260 -840 1320 -790 0 FreeSans 240 0 0 0 phi2
flabel metal2 1330 -420 1380 -370 0 FreeSans 240 0 0 0 GND
flabel metal2 1260 200 1290 230 0 FreeSans 160 0 0 0 phi2_n
flabel metal2 950 200 980 230 0 FreeSans 160 0 0 0 phi1_n
flabel metal1 1080 130 1110 160 0 FreeSans 160 0 0 0 Vdd
flabel metal4 480 -3490 550 -3420 0 FreeSans 160 0 0 0 com_x
flabel metal1 740 -940 780 -900 0 FreeSans 160 0 0 0 sub
<< end >>
