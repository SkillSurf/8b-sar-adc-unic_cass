magic
tech sky130A
timestamp 1730665161
<< metal1 >>
rect -65 2230 6775 2245
rect -65 2170 6775 2185
rect -65 2110 6775 2125
rect -65 2050 6775 2065
rect -65 1990 6775 2005
rect -65 1930 6775 1945
rect -5 1870 705 1885
rect 875 1870 1485 1885
rect 1850 1870 2390 1885
rect 2695 1870 3235 1885
rect 3540 1870 4105 1885
rect 4410 1870 4965 1885
rect 5270 1870 5835 1885
rect 6140 1870 6615 1885
rect -5 1840 705 1855
rect 875 1840 1485 1855
rect 1850 1840 2390 1855
rect 2695 1840 3235 1855
rect 3540 1840 4105 1855
rect 4410 1840 4965 1855
rect 5270 1840 5835 1855
rect 6140 1840 6615 1855
rect -5 1795 705 1810
rect 875 1795 1485 1810
rect 1850 1795 2390 1810
rect 2695 1795 3235 1810
rect 3540 1795 4105 1810
rect 4410 1795 4965 1810
rect 5270 1795 5835 1810
rect 6140 1795 6615 1810
rect -5 1745 705 1780
rect 875 1745 1485 1780
rect 1850 1745 2390 1780
rect 2695 1745 3235 1780
rect 3540 1745 4105 1780
rect 4410 1745 4965 1780
rect 5270 1745 5835 1780
rect 6140 1745 6615 1780
rect -5 1205 705 1240
rect 875 1205 1485 1240
rect 1850 1205 2390 1240
rect 2695 1205 3235 1240
rect 3540 1205 4105 1240
rect 4410 1205 4965 1240
rect 5270 1205 5835 1240
rect 6140 1205 6615 1240
rect -5 1175 705 1190
rect 875 1175 1485 1190
rect 1850 1175 2390 1190
rect 2695 1175 3235 1190
rect 3540 1175 4105 1190
rect 4410 1175 4965 1190
rect 5270 1175 5835 1190
rect 6140 1175 6615 1190
rect -65 1115 6775 1130
rect -65 1055 6775 1070
rect -65 995 6775 1010
rect -65 935 6775 950
rect -65 875 6775 890
rect -65 815 6775 830
<< metal4 >>
rect -65 -75 6775 -45
use cap_final  cap_final_0 ~/dac_lay
timestamp 1730665161
transform 1 0 -200 0 1 1680
box 135 -1795 990 205
use cap_final  cap_final_1
timestamp 1730665161
transform 1 0 5785 0 1 1680
box 135 -1795 990 205
use cap_final  cap_final_2
timestamp 1730665161
transform 1 0 655 0 1 1680
box 135 -1795 990 205
use cap_final  cap_final_3
timestamp 1730665161
transform 1 0 1510 0 1 1680
box 135 -1795 990 205
use cap_final  cap_final_4
timestamp 1730665161
transform 1 0 2365 0 1 1680
box 135 -1795 990 205
use cap_final  cap_final_5
timestamp 1730665161
transform 1 0 3220 0 1 1680
box 135 -1795 990 205
use cap_final  cap_final_6
timestamp 1730665161
transform 1 0 4075 0 1 1680
box 135 -1795 990 205
use cap_final  cap_final_7
timestamp 1730665161
transform 1 0 4930 0 1 1680
box 135 -1795 990 205
<< end >>
