magic
tech sky130A
timestamp 1730665161
<< metal1 >>
rect 6470 2300 6475 2315
rect 0 2285 6475 2300
rect 6505 2300 6510 2315
rect 7325 2300 7330 2315
rect 6505 2285 7330 2300
rect 7360 2300 7365 2315
rect 7360 2285 13680 2300
rect 5615 2240 5620 2255
rect 0 2225 5620 2240
rect 5650 2240 5655 2255
rect 8180 2240 8185 2255
rect 5650 2225 8185 2240
rect 8215 2240 8220 2255
rect 8215 2225 13680 2240
rect 4760 2180 4765 2195
rect 0 2165 4765 2180
rect 4795 2180 4800 2195
rect 9035 2180 9040 2195
rect 4795 2165 9040 2180
rect 9070 2180 9075 2195
rect 9070 2165 13680 2180
rect 3905 2120 3910 2135
rect 0 2105 3910 2120
rect 3940 2120 3945 2135
rect 9890 2120 9895 2135
rect 3940 2105 9895 2120
rect 9925 2120 9930 2135
rect 9925 2105 13680 2120
rect 2195 2060 2200 2075
rect 0 2045 2200 2060
rect 2230 2060 2235 2075
rect 3050 2060 3055 2075
rect 2230 2045 3055 2060
rect 3085 2060 3090 2075
rect 10745 2060 10750 2075
rect 3085 2045 10750 2060
rect 10780 2060 10785 2075
rect 11600 2060 11605 2075
rect 10780 2045 11605 2060
rect 11635 2060 11640 2075
rect 11635 2045 13680 2060
rect 485 2000 490 2015
rect 0 1985 490 2000
rect 520 2000 525 2015
rect 1340 2000 1345 2015
rect 520 1985 1345 2000
rect 1375 2000 1380 2015
rect 12455 2000 12460 2015
rect 1375 1985 12460 2000
rect 12490 2000 12495 2015
rect 13310 2000 13315 2015
rect 12490 1985 13315 2000
rect 13345 2000 13350 2015
rect 13345 1985 13680 2000
rect 485 1275 490 1305
rect 520 1275 525 1305
rect 1180 1290 1345 1305
rect 1340 1275 1345 1290
rect 1375 1275 1380 1305
rect 12295 1290 12460 1305
rect 12455 1275 12460 1290
rect 12490 1275 12495 1305
rect 13150 1290 13315 1305
rect 13310 1275 13315 1290
rect 13345 1275 13350 1305
rect 2035 1230 2200 1245
rect 2195 1215 2200 1230
rect 2230 1215 2235 1245
rect 2890 1230 3055 1245
rect 3050 1215 3055 1230
rect 3085 1215 3090 1245
rect 10585 1230 10750 1245
rect 10745 1215 10750 1230
rect 10780 1215 10785 1245
rect 11440 1230 11605 1245
rect 11600 1215 11605 1230
rect 11635 1230 13680 1245
rect 11635 1215 11640 1230
rect 0 1170 2035 1185
rect 3745 1170 3910 1185
rect 3905 1155 3910 1170
rect 3940 1155 3945 1185
rect 9730 1170 9895 1185
rect 9890 1155 9895 1170
rect 9925 1170 13680 1185
rect 9925 1155 9930 1170
rect 0 1110 4070 1125
rect 4600 1110 4765 1125
rect 4760 1095 4765 1110
rect 4795 1095 4800 1125
rect 8875 1110 9040 1125
rect 9035 1095 9040 1110
rect 9070 1110 13680 1125
rect 9070 1095 9075 1110
rect 0 1050 4070 1065
rect 5455 1050 5620 1065
rect 5615 1035 5620 1050
rect 5650 1035 5655 1065
rect 8020 1050 8185 1065
rect 8180 1035 8185 1050
rect 8215 1050 13680 1065
rect 8215 1035 8220 1050
rect 0 990 4070 1005
rect 6310 990 6475 1005
rect 6470 975 6475 990
rect 6505 975 6510 1005
rect 7165 990 7330 1005
rect 7325 975 7330 990
rect 7360 990 7465 1005
rect 9705 990 13680 1005
rect 7360 975 7365 990
<< via1 >>
rect 6475 2285 6505 2315
rect 7330 2285 7360 2315
rect 5620 2225 5650 2255
rect 8185 2225 8215 2255
rect 4765 2165 4795 2195
rect 9040 2165 9070 2195
rect 3910 2105 3940 2135
rect 9895 2105 9925 2135
rect 2200 2045 2230 2075
rect 3055 2045 3085 2075
rect 10750 2045 10780 2075
rect 11605 2045 11635 2075
rect 490 1985 520 2015
rect 1345 1985 1375 2015
rect 12460 1985 12490 2015
rect 13315 1985 13345 2015
rect 490 1275 520 1305
rect 1345 1275 1375 1305
rect 12460 1275 12490 1305
rect 13315 1275 13345 1305
rect 2200 1215 2230 1245
rect 3055 1215 3085 1245
rect 10750 1215 10780 1245
rect 11605 1215 11635 1245
rect 3910 1155 3940 1185
rect 9895 1155 9925 1185
rect 4765 1095 4795 1125
rect 9040 1095 9070 1125
rect 5620 1035 5650 1065
rect 8185 1035 8215 1065
rect 6475 975 6505 1005
rect 7330 975 7360 1005
<< metal2 >>
rect 6310 2320 6350 2325
rect 6310 2300 6315 2320
rect 0 2290 6315 2300
rect 6345 2290 6350 2320
rect 7165 2320 7205 2325
rect 0 2285 6350 2290
rect 6470 2285 6475 2315
rect 6505 2285 6510 2315
rect 7165 2290 7170 2320
rect 7200 2290 7205 2320
rect 7425 2320 7465 2325
rect 7165 2285 7205 2290
rect 7325 2285 7330 2315
rect 7360 2285 7365 2315
rect 7425 2290 7430 2320
rect 7460 2300 7465 2320
rect 7460 2290 13680 2300
rect 7425 2285 13680 2290
rect 5455 2260 5495 2265
rect 5455 2240 5460 2260
rect 0 2230 5460 2240
rect 5490 2230 5495 2260
rect 0 2225 5495 2230
rect 5615 2225 5620 2255
rect 5650 2225 5655 2255
rect 4600 2200 4640 2205
rect 4600 2180 4605 2200
rect 0 2170 4605 2180
rect 4635 2170 4640 2200
rect 0 2165 4640 2170
rect 4760 2165 4765 2195
rect 4795 2165 4800 2195
rect 3745 2140 3785 2145
rect 3745 2120 3750 2140
rect 0 2110 3750 2120
rect 3780 2110 3785 2140
rect 0 2105 3785 2110
rect 3905 2105 3910 2135
rect 3940 2105 3945 2135
rect 2035 2080 2075 2085
rect 2035 2060 2040 2080
rect 0 2050 2040 2060
rect 2070 2050 2075 2080
rect 2890 2080 2930 2085
rect 0 2045 2075 2050
rect 2195 2045 2200 2075
rect 2230 2045 2235 2075
rect 2890 2050 2895 2080
rect 2925 2050 2930 2080
rect 2890 2045 2930 2050
rect 3050 2045 3055 2075
rect 3085 2045 3090 2075
rect 325 2020 365 2025
rect 325 2000 330 2020
rect 0 1990 330 2000
rect 360 1990 365 2020
rect 1180 2020 1220 2025
rect 0 1985 365 1990
rect 485 1985 490 2015
rect 520 1985 525 2015
rect 1180 1990 1185 2020
rect 1215 1990 1220 2020
rect 1180 1985 1220 1990
rect 1340 1985 1345 2015
rect 1375 1985 1380 2015
rect 340 1970 355 1985
rect 495 1970 510 1985
rect 1195 1970 1210 1985
rect 1350 1970 1365 1985
rect 2050 1970 2065 2045
rect 2205 1970 2220 2045
rect 2905 1970 2920 2045
rect 3060 1970 3075 2045
rect 3760 1970 3775 2105
rect 3915 1970 3930 2105
rect 4615 1970 4630 2165
rect 4770 1970 4785 2165
rect 5470 1970 5485 2225
rect 5625 1970 5640 2225
rect 6325 1970 6340 2285
rect 6480 1970 6495 2285
rect 7180 1970 7195 2285
rect 7335 1970 7350 2285
rect 8020 2260 8060 2265
rect 8020 2230 8025 2260
rect 8055 2230 8060 2260
rect 8280 2260 8320 2265
rect 8020 2225 8060 2230
rect 8180 2225 8185 2255
rect 8215 2225 8220 2255
rect 8280 2230 8285 2260
rect 8315 2240 8320 2260
rect 8315 2230 13680 2240
rect 8280 2225 13680 2230
rect 8035 1970 8050 2225
rect 8190 1970 8205 2225
rect 8875 2200 8915 2205
rect 8875 2170 8880 2200
rect 8910 2170 8915 2200
rect 9135 2200 9175 2205
rect 8875 2165 8915 2170
rect 9035 2165 9040 2195
rect 9070 2165 9075 2195
rect 9135 2170 9140 2200
rect 9170 2180 9175 2200
rect 9170 2170 13680 2180
rect 9135 2165 13680 2170
rect 8890 1970 8905 2165
rect 9045 1970 9060 2165
rect 9730 2140 9770 2145
rect 9730 2110 9735 2140
rect 9765 2110 9770 2140
rect 9990 2140 10030 2145
rect 9730 2105 9770 2110
rect 9890 2105 9895 2135
rect 9925 2105 9930 2135
rect 9990 2110 9995 2140
rect 10025 2120 10030 2140
rect 10025 2110 13680 2120
rect 9990 2105 13680 2110
rect 9745 1970 9760 2105
rect 9900 1970 9915 2105
rect 10585 2080 10625 2085
rect 10585 2050 10590 2080
rect 10620 2050 10625 2080
rect 11440 2080 11480 2085
rect 10585 2045 10625 2050
rect 10745 2045 10750 2075
rect 10780 2045 10785 2075
rect 11440 2050 11445 2080
rect 11475 2050 11480 2080
rect 11700 2080 11740 2085
rect 11440 2045 11480 2050
rect 11600 2045 11605 2075
rect 11635 2045 11640 2075
rect 11700 2050 11705 2080
rect 11735 2060 11740 2080
rect 11735 2050 13680 2060
rect 11700 2045 13680 2050
rect 10600 1970 10615 2045
rect 10755 1970 10770 2045
rect 11455 1970 11470 2045
rect 11610 1970 11625 2045
rect 12295 2020 12335 2025
rect 12295 1990 12300 2020
rect 12330 1990 12335 2020
rect 13150 2020 13190 2025
rect 12295 1985 12335 1990
rect 12455 1985 12460 2015
rect 12490 1985 12495 2015
rect 13150 1990 13155 2020
rect 13185 1990 13190 2020
rect 13410 2020 13450 2025
rect 13150 1985 13190 1990
rect 13310 1985 13315 2015
rect 13345 1985 13350 2015
rect 13410 1990 13415 2020
rect 13445 2000 13450 2020
rect 13445 1990 13680 2000
rect 13410 1985 13680 1990
rect 12310 1970 12325 1985
rect 12465 1970 12480 1985
rect 13165 1970 13180 1985
rect 13320 1970 13335 1985
rect 340 1305 355 1310
rect 495 1305 510 1310
rect 1195 1305 1210 1310
rect 1350 1305 1365 1310
rect 0 1300 365 1305
rect 0 1290 330 1300
rect 325 1270 330 1290
rect 360 1270 365 1300
rect 485 1275 490 1305
rect 520 1275 525 1305
rect 1180 1300 1220 1305
rect 325 1265 365 1270
rect 1180 1270 1185 1300
rect 1215 1270 1220 1300
rect 1340 1275 1345 1305
rect 1375 1275 1380 1305
rect 1180 1265 1220 1270
rect 2050 1245 2065 1310
rect 2205 1245 2220 1310
rect 2905 1245 2920 1310
rect 3060 1245 3075 1310
rect 0 1240 2075 1245
rect 0 1230 2040 1240
rect 2035 1210 2040 1230
rect 2070 1210 2075 1240
rect 2195 1215 2200 1245
rect 2230 1215 2235 1245
rect 2890 1240 2930 1245
rect 2035 1205 2075 1210
rect 2890 1210 2895 1240
rect 2925 1210 2930 1240
rect 3050 1215 3055 1245
rect 3085 1215 3090 1245
rect 2890 1205 2930 1210
rect 3760 1185 3775 1310
rect 3915 1185 3930 1310
rect 0 1180 3785 1185
rect 0 1170 3750 1180
rect 3745 1150 3750 1170
rect 3780 1150 3785 1180
rect 3905 1155 3910 1185
rect 3940 1155 3945 1185
rect 3745 1145 3785 1150
rect 4615 1125 4630 1310
rect 4770 1125 4785 1310
rect 0 1120 4640 1125
rect 0 1110 4605 1120
rect 4600 1090 4605 1110
rect 4635 1090 4640 1120
rect 4760 1095 4765 1125
rect 4795 1095 4800 1125
rect 4600 1085 4640 1090
rect 5470 1065 5485 1310
rect 5625 1065 5640 1310
rect 0 1060 5495 1065
rect 0 1050 5460 1060
rect 5455 1030 5460 1050
rect 5490 1030 5495 1060
rect 5615 1035 5620 1065
rect 5650 1035 5655 1065
rect 5455 1025 5495 1030
rect 6325 1005 6340 1310
rect 6480 1005 6495 1310
rect 7180 1005 7195 1310
rect 7335 1005 7350 1310
rect 8035 1065 8050 1310
rect 8190 1065 8205 1310
rect 8890 1125 8905 1310
rect 9045 1125 9060 1310
rect 9745 1185 9760 1310
rect 9900 1185 9915 1310
rect 10600 1245 10615 1310
rect 10755 1245 10770 1310
rect 11455 1245 11470 1310
rect 11610 1245 11625 1310
rect 12310 1305 12325 1310
rect 12465 1305 12480 1310
rect 13165 1305 13180 1310
rect 13320 1305 13335 1310
rect 12295 1300 12335 1305
rect 12295 1270 12300 1300
rect 12330 1270 12335 1300
rect 12455 1275 12460 1305
rect 12490 1275 12495 1305
rect 13150 1300 13190 1305
rect 12295 1265 12335 1270
rect 13150 1270 13155 1300
rect 13185 1270 13190 1300
rect 13310 1275 13315 1305
rect 13345 1275 13350 1305
rect 13410 1300 13680 1305
rect 13150 1265 13190 1270
rect 13410 1270 13415 1300
rect 13445 1290 13680 1300
rect 13445 1270 13450 1290
rect 13410 1265 13450 1270
rect 10585 1240 10625 1245
rect 10585 1210 10590 1240
rect 10620 1210 10625 1240
rect 10745 1215 10750 1245
rect 10780 1215 10785 1245
rect 11440 1240 11480 1245
rect 10585 1205 10625 1210
rect 11440 1210 11445 1240
rect 11475 1210 11480 1240
rect 11600 1215 11605 1245
rect 11635 1215 11640 1245
rect 11700 1240 13680 1245
rect 11440 1205 11480 1210
rect 11700 1210 11705 1240
rect 11735 1230 13680 1240
rect 11735 1210 11740 1230
rect 11700 1205 11740 1210
rect 9730 1180 9770 1185
rect 9730 1150 9735 1180
rect 9765 1150 9770 1180
rect 9890 1155 9895 1185
rect 9925 1155 9930 1185
rect 9990 1180 13680 1185
rect 9730 1145 9770 1150
rect 9990 1150 9995 1180
rect 10025 1170 13680 1180
rect 10025 1150 10030 1170
rect 9990 1145 10030 1150
rect 8875 1120 8915 1125
rect 8875 1090 8880 1120
rect 8910 1090 8915 1120
rect 9035 1095 9040 1125
rect 9070 1095 9075 1125
rect 9135 1120 13680 1125
rect 8875 1085 8915 1090
rect 9135 1090 9140 1120
rect 9170 1110 13680 1120
rect 9170 1090 9175 1110
rect 9135 1085 9175 1090
rect 8020 1060 8060 1065
rect 8020 1030 8025 1060
rect 8055 1030 8060 1060
rect 8180 1035 8185 1065
rect 8215 1035 8220 1065
rect 8280 1060 13680 1065
rect 8020 1025 8060 1030
rect 8280 1030 8285 1060
rect 8315 1050 13680 1060
rect 8315 1030 8320 1050
rect 8280 1025 8320 1030
rect 0 1000 6350 1005
rect 0 990 6315 1000
rect 6310 970 6315 990
rect 6345 970 6350 1000
rect 6470 975 6475 1005
rect 6505 975 6510 1005
rect 7165 1000 7205 1005
rect 6310 965 6350 970
rect 7165 970 7170 1000
rect 7200 970 7205 1000
rect 7325 975 7330 1005
rect 7360 975 7365 1005
rect 7425 1000 13680 1005
rect 7165 965 7205 970
rect 7425 970 7430 1000
rect 7460 990 13680 1000
rect 7460 970 7465 990
rect 7425 965 7465 970
<< via2 >>
rect 6315 2290 6345 2320
rect 7170 2290 7200 2320
rect 7430 2290 7460 2320
rect 5460 2230 5490 2260
rect 4605 2170 4635 2200
rect 3750 2110 3780 2140
rect 2040 2050 2070 2080
rect 2895 2050 2925 2080
rect 330 1990 360 2020
rect 1185 1990 1215 2020
rect 8025 2230 8055 2260
rect 8285 2230 8315 2260
rect 8880 2170 8910 2200
rect 9140 2170 9170 2200
rect 9735 2110 9765 2140
rect 9995 2110 10025 2140
rect 10590 2050 10620 2080
rect 11445 2050 11475 2080
rect 11705 2050 11735 2080
rect 12300 1990 12330 2020
rect 13155 1990 13185 2020
rect 13415 1990 13445 2020
rect 330 1270 360 1300
rect 1185 1270 1215 1300
rect 2040 1210 2070 1240
rect 2895 1210 2925 1240
rect 3750 1150 3780 1180
rect 4605 1090 4635 1120
rect 5460 1030 5490 1060
rect 12300 1270 12330 1300
rect 13155 1270 13185 1300
rect 13415 1270 13445 1300
rect 10590 1210 10620 1240
rect 11445 1210 11475 1240
rect 11705 1210 11735 1240
rect 9735 1150 9765 1180
rect 9995 1150 10025 1180
rect 8880 1090 8910 1120
rect 9140 1090 9170 1120
rect 8025 1030 8055 1060
rect 8285 1030 8315 1060
rect 6315 970 6345 1000
rect 7170 970 7200 1000
rect 7430 970 7460 1000
<< metal3 >>
rect 6310 2320 6350 2325
rect 6310 2290 6315 2320
rect 6345 2315 6350 2320
rect 7165 2320 7205 2325
rect 7165 2315 7170 2320
rect 6345 2290 7170 2315
rect 7200 2315 7205 2320
rect 7425 2320 7465 2325
rect 7425 2315 7430 2320
rect 7200 2290 7430 2315
rect 7460 2290 7465 2320
rect 6310 2285 7465 2290
rect 5455 2260 5495 2265
rect 5455 2230 5460 2260
rect 5490 2255 5495 2260
rect 8020 2260 8060 2265
rect 8020 2255 8025 2260
rect 5490 2230 8025 2255
rect 8055 2255 8060 2260
rect 8280 2260 8320 2265
rect 8280 2255 8285 2260
rect 8055 2230 8285 2255
rect 8315 2230 8320 2260
rect 5455 2225 8320 2230
rect 4600 2200 4640 2205
rect 4600 2170 4605 2200
rect 4635 2195 4640 2200
rect 8875 2200 8915 2205
rect 8875 2195 8880 2200
rect 4635 2170 8880 2195
rect 8910 2195 8915 2200
rect 9135 2200 9175 2205
rect 9135 2195 9140 2200
rect 8910 2170 9140 2195
rect 9170 2170 9175 2200
rect 4600 2165 9175 2170
rect 3745 2140 3785 2145
rect 3745 2110 3750 2140
rect 3780 2135 3785 2140
rect 9730 2140 9770 2145
rect 9730 2135 9735 2140
rect 3780 2110 9735 2135
rect 9765 2135 9770 2140
rect 9990 2140 10030 2145
rect 9990 2135 9995 2140
rect 9765 2110 9995 2135
rect 10025 2110 10030 2140
rect 3745 2105 10030 2110
rect 2035 2080 2075 2085
rect 2035 2050 2040 2080
rect 2070 2075 2075 2080
rect 2890 2080 2930 2085
rect 2890 2075 2895 2080
rect 2070 2050 2895 2075
rect 2925 2075 2930 2080
rect 10585 2080 10625 2085
rect 10585 2075 10590 2080
rect 2925 2050 10590 2075
rect 10620 2075 10625 2080
rect 11440 2080 11480 2085
rect 11440 2075 11445 2080
rect 10620 2050 11445 2075
rect 11475 2075 11480 2080
rect 11700 2080 11740 2085
rect 11700 2075 11705 2080
rect 11475 2050 11705 2075
rect 11735 2050 11740 2080
rect 2035 2045 11740 2050
rect 325 2020 365 2025
rect 325 1990 330 2020
rect 360 2015 365 2020
rect 1180 2020 1220 2025
rect 1180 2015 1185 2020
rect 360 1990 1185 2015
rect 1215 2015 1220 2020
rect 12295 2020 12335 2025
rect 12295 2015 12300 2020
rect 1215 1990 12300 2015
rect 12330 2015 12335 2020
rect 13150 2020 13190 2025
rect 13150 2015 13155 2020
rect 12330 1990 13155 2015
rect 13185 2015 13190 2020
rect 13410 2020 13450 2025
rect 13410 2015 13415 2020
rect 13185 1990 13415 2015
rect 13445 1990 13450 2020
rect 325 1985 13450 1990
rect 325 1300 13450 1305
rect 325 1270 330 1300
rect 360 1275 1185 1300
rect 360 1270 365 1275
rect 325 1265 365 1270
rect 1180 1270 1185 1275
rect 1215 1275 12300 1300
rect 1215 1270 1220 1275
rect 1180 1265 1220 1270
rect 12295 1270 12300 1275
rect 12330 1275 13155 1300
rect 12330 1270 12335 1275
rect 12295 1265 12335 1270
rect 13150 1270 13155 1275
rect 13185 1275 13415 1300
rect 13185 1270 13190 1275
rect 13150 1265 13190 1270
rect 13410 1270 13415 1275
rect 13445 1270 13450 1300
rect 13410 1265 13450 1270
rect 2035 1240 11740 1245
rect 2035 1210 2040 1240
rect 2070 1215 2895 1240
rect 2070 1210 2075 1215
rect 2035 1205 2075 1210
rect 2890 1210 2895 1215
rect 2925 1215 10590 1240
rect 2925 1210 2930 1215
rect 2890 1205 2930 1210
rect 10585 1210 10590 1215
rect 10620 1215 11445 1240
rect 10620 1210 10625 1215
rect 10585 1205 10625 1210
rect 11440 1210 11445 1215
rect 11475 1215 11705 1240
rect 11475 1210 11480 1215
rect 11440 1205 11480 1210
rect 11700 1210 11705 1215
rect 11735 1210 11740 1240
rect 11700 1205 11740 1210
rect 3745 1180 10030 1185
rect 3745 1150 3750 1180
rect 3780 1155 9735 1180
rect 3780 1150 3785 1155
rect 3745 1145 3785 1150
rect 9730 1150 9735 1155
rect 9765 1155 9995 1180
rect 9765 1150 9770 1155
rect 9730 1145 9770 1150
rect 9990 1150 9995 1155
rect 10025 1150 10030 1180
rect 9990 1145 10030 1150
rect 4600 1120 9175 1125
rect 4600 1090 4605 1120
rect 4635 1095 8880 1120
rect 4635 1090 4640 1095
rect 4600 1085 4640 1090
rect 8875 1090 8880 1095
rect 8910 1095 9140 1120
rect 8910 1090 8915 1095
rect 8875 1085 8915 1090
rect 9135 1090 9140 1095
rect 9170 1090 9175 1120
rect 9135 1085 9175 1090
rect 5455 1060 8320 1065
rect 5455 1030 5460 1060
rect 5490 1035 8025 1060
rect 5490 1030 5495 1035
rect 5455 1025 5495 1030
rect 8020 1030 8025 1035
rect 8055 1035 8285 1060
rect 8055 1030 8060 1035
rect 8020 1025 8060 1030
rect 8280 1030 8285 1035
rect 8315 1030 8320 1060
rect 8280 1025 8320 1030
rect 6310 1000 7465 1005
rect 6310 970 6315 1000
rect 6345 975 7170 1000
rect 6345 970 6350 975
rect 6310 965 6350 970
rect 7165 970 7170 975
rect 7200 975 7430 1000
rect 7200 970 7205 975
rect 7165 965 7205 970
rect 7425 970 7430 975
rect 7460 970 7465 1000
rect 7425 965 7465 970
<< metal4 >>
rect 410 1985 440 2330
rect 1265 1985 1295 2330
rect 2120 1985 2150 2330
rect 2975 1985 3005 2330
rect 3830 1985 3860 2330
rect 4685 1985 4715 2330
rect 5540 1985 5570 2330
rect 6395 1985 6425 2330
rect 7250 1985 7280 2330
rect 8105 1985 8135 2330
rect 8960 1985 8990 2330
rect 9815 1985 9845 2330
rect 10670 1985 10700 2330
rect 11525 1985 11555 2330
rect 12380 1985 12410 2330
rect 13235 1985 13265 2330
use 8_cap_array_final  8_cap_array_final_0
timestamp 1730665161
transform 1 0 65 0 1 115
box -65 -115 6775 2245
use 8_cap_array_final  8_cap_array_final_1
timestamp 1730665161
transform 1 0 6905 0 1 115
box -65 -115 6775 2245
<< end >>
