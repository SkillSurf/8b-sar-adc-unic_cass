magic
tech sky130A
magscale 1 2
timestamp 1728835232
<< metal3 >>
rect -886 712 886 740
rect -886 -712 802 712
rect 866 -712 886 712
rect -886 -740 886 -712
<< via3 >>
rect 802 -712 866 712
<< mimcap >>
rect -846 660 554 700
rect -846 -660 -806 660
rect 514 -660 554 660
rect -846 -700 554 -660
<< mimcapcontact >>
rect -806 -660 514 660
<< metal4 >>
rect 786 712 882 728
rect -807 660 515 661
rect -807 -660 -806 660
rect 514 -660 515 660
rect -807 -661 515 -660
rect 786 -712 802 712
rect 866 -712 882 712
rect 786 -728 882 -712
<< properties >>
string FIXED_BBOX -886 -740 594 740
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 7.00 l 7.00 val 103.32 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
