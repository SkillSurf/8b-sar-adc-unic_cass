magic
tech sky130A
timestamp 1730665161
<< metal1 >>
rect 930 -465 945 0
rect 2345 -355 2360 -225
rect 915 -485 945 -480
rect 915 -520 945 -515
rect 2345 -485 2375 -480
rect 2345 -520 2375 -515
rect 930 -6840 945 -550
rect 2345 -590 2360 -535
rect 990 -6840 1005 -625
rect 1050 -1265 1065 -1185
rect 1050 -1340 1065 -1295
rect 1035 -1345 1065 -1340
rect 1035 -1380 1065 -1375
rect 2225 -1340 2240 -1185
rect 2225 -1345 2255 -1340
rect 2225 -1380 2255 -1375
rect 1050 -6840 1065 -1380
rect 1110 -2120 1125 -2040
rect 1110 -2195 1125 -2150
rect 1095 -2200 1125 -2195
rect 1095 -2235 1125 -2230
rect 1110 -2340 1125 -2235
rect 2165 -2195 2180 -2040
rect 2165 -2200 2195 -2195
rect 2165 -2235 2195 -2230
rect 2165 -2340 2180 -2235
rect 1170 -2975 1185 -2895
rect 1170 -3050 1185 -3005
rect 1155 -3055 1185 -3050
rect 1155 -3090 1185 -3085
rect 1170 -3195 1185 -3090
rect 2105 -3050 2120 -2895
rect 2105 -3055 2135 -3050
rect 2105 -3090 2135 -3085
rect 2105 -3195 2120 -3090
rect 1110 -6840 1125 -3195
rect 1230 -3830 1245 -3750
rect 1230 -3905 1245 -3860
rect 1215 -3910 1245 -3905
rect 1215 -3945 1245 -3940
rect 2045 -3905 2060 -3750
rect 2045 -3910 2075 -3905
rect 2045 -3945 2075 -3940
rect 1230 -4760 1245 -4605
rect 1215 -4765 1245 -4760
rect 1215 -4800 1245 -4795
rect 1230 -4905 1245 -4800
rect 2045 -4760 2060 -4605
rect 2045 -4765 2075 -4760
rect 2045 -4800 2075 -4795
rect 2045 -4905 2060 -4800
rect 1170 -6840 1185 -4905
rect 1290 -5540 1305 -5460
rect 1290 -5615 1305 -5570
rect 1275 -5620 1305 -5615
rect 1275 -5655 1305 -5650
rect 1985 -5615 2000 -5460
rect 1985 -5620 2015 -5615
rect 1985 -5655 2015 -5650
rect 1290 -6470 1305 -6315
rect 1275 -6475 1305 -6470
rect 1275 -6510 1305 -6505
rect 1290 -6615 1305 -6510
rect 1985 -6470 2000 -6315
rect 1985 -6475 2015 -6470
rect 1985 -6510 2015 -6505
rect 1985 -6615 2000 -6510
rect 1230 -6840 1245 -6615
rect 2105 -6840 2120 -4905
rect 2165 -6840 2180 -3195
rect 2225 -6840 2240 -2340
rect 2285 -6840 2300 -1485
rect 2345 -6840 2360 -1485
<< via1 >>
rect 915 -515 945 -485
rect 2345 -515 2375 -485
rect 1035 -1375 1065 -1345
rect 2225 -1375 2255 -1345
rect 1095 -2230 1125 -2200
rect 2165 -2230 2195 -2200
rect 1155 -3085 1185 -3055
rect 2105 -3085 2135 -3055
rect 1215 -3940 1245 -3910
rect 2045 -3940 2075 -3910
rect 1215 -4795 1245 -4765
rect 2045 -4795 2075 -4765
rect 1275 -5650 1305 -5620
rect 1985 -5650 2015 -5620
rect 1275 -6505 1305 -6475
rect 1985 -6505 2015 -6475
<< metal2 >>
rect 930 -340 945 0
rect 2345 -340 2360 0
rect 930 -355 1310 -340
rect 1980 -355 2360 -340
rect 930 -450 945 -355
rect 885 -465 945 -450
rect 2345 -450 2360 -355
rect 2345 -465 2405 -450
rect 885 -535 900 -465
rect 915 -485 945 -480
rect 2345 -485 2375 -480
rect 945 -510 1310 -495
rect 1980 -510 2345 -495
rect 915 -520 945 -515
rect 2345 -520 2375 -515
rect 2390 -535 2405 -465
rect 885 -550 945 -535
rect 930 -6840 945 -550
rect 2345 -550 2405 -535
rect 965 -590 1005 -585
rect 965 -620 970 -590
rect 1000 -620 1005 -590
rect 965 -625 1005 -620
rect 990 -6840 1005 -625
rect 2285 -615 2325 -610
rect 2285 -645 2290 -615
rect 2320 -645 2325 -615
rect 2285 -650 2325 -645
rect 1025 -1190 1065 -1185
rect 1025 -1220 1030 -1190
rect 1060 -1195 1065 -1190
rect 2225 -1190 2265 -1185
rect 2225 -1195 2230 -1190
rect 1060 -1210 1310 -1195
rect 1980 -1210 2230 -1195
rect 1060 -1220 1065 -1210
rect 1025 -1225 1065 -1220
rect 2225 -1220 2230 -1210
rect 2260 -1220 2265 -1190
rect 2225 -1225 2265 -1220
rect 1035 -1345 1065 -1340
rect 2225 -1345 2255 -1340
rect 1065 -1365 1310 -1350
rect 1980 -1365 2225 -1350
rect 1035 -1380 1065 -1375
rect 2225 -1380 2255 -1375
rect 1025 -1450 1065 -1445
rect 1025 -1480 1030 -1450
rect 1060 -1480 1065 -1450
rect 1025 -1485 1065 -1480
rect 1050 -6840 1065 -1485
rect 2225 -1450 2265 -1445
rect 2225 -1480 2230 -1450
rect 2260 -1480 2265 -1450
rect 2225 -1485 2265 -1480
rect 1085 -2045 1125 -2040
rect 1085 -2075 1090 -2045
rect 1120 -2050 1125 -2045
rect 2165 -2045 2205 -2040
rect 2165 -2050 2170 -2045
rect 1120 -2065 1315 -2050
rect 1980 -2065 2170 -2050
rect 1120 -2075 1125 -2065
rect 1085 -2080 1125 -2075
rect 2165 -2075 2170 -2065
rect 2200 -2075 2205 -2045
rect 2165 -2080 2205 -2075
rect 1095 -2200 1125 -2195
rect 2165 -2200 2195 -2195
rect 1125 -2220 1315 -2205
rect 1980 -2220 2165 -2205
rect 1095 -2235 1125 -2230
rect 2165 -2235 2195 -2230
rect 1085 -2305 1125 -2300
rect 1085 -2335 1090 -2305
rect 1120 -2335 1125 -2305
rect 1085 -2340 1125 -2335
rect 1110 -6840 1125 -2340
rect 2165 -2305 2205 -2300
rect 2165 -2335 2170 -2305
rect 2200 -2335 2205 -2305
rect 2165 -2340 2205 -2335
rect 1145 -2900 1185 -2895
rect 1145 -2930 1150 -2900
rect 1180 -2905 1185 -2900
rect 2105 -2900 2145 -2895
rect 2105 -2905 2110 -2900
rect 1180 -2920 1310 -2905
rect 1980 -2920 2110 -2905
rect 1180 -2930 1185 -2920
rect 1145 -2935 1185 -2930
rect 2105 -2930 2110 -2920
rect 2140 -2930 2145 -2900
rect 2105 -2935 2145 -2930
rect 1155 -3055 1185 -3050
rect 2105 -3055 2135 -3050
rect 1185 -3075 1310 -3060
rect 1980 -3075 2105 -3060
rect 1155 -3090 1185 -3085
rect 2105 -3090 2135 -3085
rect 1145 -3160 1185 -3155
rect 1145 -3190 1150 -3160
rect 1180 -3190 1185 -3160
rect 1145 -3195 1185 -3190
rect 1170 -6840 1185 -3195
rect 2105 -3160 2145 -3155
rect 2105 -3190 2110 -3160
rect 2140 -3190 2145 -3160
rect 2105 -3195 2145 -3190
rect 1205 -3755 1245 -3750
rect 1205 -3785 1210 -3755
rect 1240 -3760 1245 -3755
rect 2045 -3755 2085 -3750
rect 2045 -3760 2050 -3755
rect 1240 -3775 1310 -3760
rect 1980 -3775 2050 -3760
rect 1240 -3785 1245 -3775
rect 1205 -3790 1245 -3785
rect 2045 -3785 2050 -3775
rect 2080 -3785 2085 -3755
rect 2045 -3790 2085 -3785
rect 1215 -3910 1245 -3905
rect 2045 -3910 2075 -3905
rect 1245 -3930 1310 -3915
rect 1980 -3930 2045 -3915
rect 1215 -3945 1245 -3940
rect 2045 -3945 2075 -3940
rect 1205 -4610 1245 -4605
rect 1205 -4640 1210 -4610
rect 1240 -4615 1245 -4610
rect 2045 -4610 2085 -4605
rect 2045 -4615 2050 -4610
rect 1240 -4630 1310 -4615
rect 1980 -4630 2050 -4615
rect 1240 -4640 1245 -4630
rect 1205 -4645 1245 -4640
rect 2045 -4640 2050 -4630
rect 2080 -4640 2085 -4610
rect 2045 -4645 2085 -4640
rect 1215 -4765 1245 -4760
rect 2045 -4765 2075 -4760
rect 1245 -4785 1310 -4770
rect 1980 -4785 2045 -4770
rect 1215 -4800 1245 -4795
rect 2045 -4800 2075 -4795
rect 1205 -4870 1245 -4865
rect 1205 -4900 1210 -4870
rect 1240 -4900 1245 -4870
rect 1205 -4905 1245 -4900
rect 1230 -6840 1245 -4905
rect 2045 -4870 2085 -4865
rect 2045 -4900 2050 -4870
rect 2080 -4900 2085 -4870
rect 2045 -4905 2085 -4900
rect 1265 -5465 1305 -5460
rect 1265 -5495 1270 -5465
rect 1300 -5470 1305 -5465
rect 1985 -5465 2025 -5460
rect 1985 -5470 1990 -5465
rect 1300 -5485 1310 -5470
rect 1980 -5485 1990 -5470
rect 1300 -5495 1305 -5485
rect 1265 -5500 1305 -5495
rect 1985 -5495 1990 -5485
rect 2020 -5495 2025 -5465
rect 1985 -5500 2025 -5495
rect 1275 -5620 1305 -5615
rect 1985 -5620 2015 -5615
rect 1305 -5640 1310 -5625
rect 1980 -5640 1985 -5625
rect 1275 -5655 1305 -5650
rect 1985 -5655 2015 -5650
rect 1265 -6320 1305 -6315
rect 1265 -6350 1270 -6320
rect 1300 -6325 1305 -6320
rect 1985 -6320 2025 -6315
rect 1985 -6325 1990 -6320
rect 1300 -6340 1310 -6325
rect 1980 -6340 1990 -6325
rect 1300 -6350 1305 -6340
rect 1265 -6355 1305 -6350
rect 1985 -6350 1990 -6340
rect 2020 -6350 2025 -6320
rect 1985 -6355 2025 -6350
rect 1275 -6475 1305 -6470
rect 1985 -6475 2015 -6470
rect 1305 -6495 1310 -6480
rect 1980 -6495 1985 -6480
rect 1275 -6510 1305 -6505
rect 1985 -6510 2015 -6505
rect 1265 -6580 1305 -6575
rect 1265 -6610 1270 -6580
rect 1300 -6610 1305 -6580
rect 1265 -6615 1305 -6610
rect 1290 -6840 1305 -6615
rect 1985 -6580 2025 -6575
rect 1985 -6610 1990 -6580
rect 2020 -6610 2025 -6580
rect 1985 -6615 2025 -6610
rect 1985 -6840 2000 -6615
rect 2045 -6840 2060 -4905
rect 2105 -6840 2120 -3195
rect 2165 -6840 2180 -2340
rect 2225 -6840 2240 -1485
rect 2285 -6840 2300 -650
rect 2345 -6840 2360 -550
<< via2 >>
rect 970 -620 1000 -590
rect 2290 -645 2320 -615
rect 1030 -1220 1060 -1190
rect 2230 -1220 2260 -1190
rect 1030 -1480 1060 -1450
rect 2230 -1480 2260 -1450
rect 1090 -2075 1120 -2045
rect 2170 -2075 2200 -2045
rect 1090 -2335 1120 -2305
rect 2170 -2335 2200 -2305
rect 1150 -2930 1180 -2900
rect 2110 -2930 2140 -2900
rect 1150 -3190 1180 -3160
rect 2110 -3190 2140 -3160
rect 1210 -3785 1240 -3755
rect 2050 -3785 2080 -3755
rect 1210 -4640 1240 -4610
rect 2050 -4640 2080 -4610
rect 1210 -4900 1240 -4870
rect 2050 -4900 2080 -4870
rect 1270 -5495 1300 -5465
rect 1990 -5495 2020 -5465
rect 1270 -6350 1300 -6320
rect 1990 -6350 2020 -6320
rect 1270 -6610 1300 -6580
rect 1990 -6610 2020 -6580
<< metal3 >>
rect 975 -585 1005 0
rect 965 -590 1005 -585
rect 965 -620 970 -590
rect 1000 -620 1005 -590
rect 965 -625 1005 -620
rect 1035 -1185 1065 0
rect 1025 -1190 1065 -1185
rect 1025 -1220 1030 -1190
rect 1060 -1220 1065 -1190
rect 1025 -1225 1065 -1220
rect 1035 -1445 1065 -1225
rect 1025 -1450 1065 -1445
rect 1025 -1480 1030 -1450
rect 1060 -1480 1065 -1450
rect 1025 -1485 1065 -1480
rect 1095 -2040 1125 0
rect 1085 -2045 1125 -2040
rect 1085 -2075 1090 -2045
rect 1120 -2075 1125 -2045
rect 1085 -2080 1125 -2075
rect 1095 -2300 1125 -2080
rect 1085 -2305 1125 -2300
rect 1085 -2335 1090 -2305
rect 1120 -2335 1125 -2305
rect 1085 -2340 1125 -2335
rect 1155 -2895 1185 0
rect 1145 -2900 1185 -2895
rect 1145 -2930 1150 -2900
rect 1180 -2930 1185 -2900
rect 1145 -2935 1185 -2930
rect 1155 -3155 1185 -2935
rect 1145 -3160 1185 -3155
rect 1145 -3190 1150 -3160
rect 1180 -3190 1185 -3160
rect 1145 -3195 1185 -3190
rect 1215 -3750 1245 0
rect 1205 -3755 1245 -3750
rect 1205 -3785 1210 -3755
rect 1240 -3785 1245 -3755
rect 1205 -3790 1245 -3785
rect 1215 -4605 1245 -3790
rect 1205 -4610 1245 -4605
rect 1205 -4640 1210 -4610
rect 1240 -4640 1245 -4610
rect 1205 -4645 1245 -4640
rect 1215 -4865 1245 -4645
rect 1205 -4870 1245 -4865
rect 1205 -4900 1210 -4870
rect 1240 -4900 1245 -4870
rect 1205 -4905 1245 -4900
rect 1275 -5460 1305 0
rect 1265 -5465 1305 -5460
rect 1265 -5495 1270 -5465
rect 1300 -5495 1305 -5465
rect 1265 -5500 1305 -5495
rect 1275 -6315 1305 -5500
rect 1265 -6320 1305 -6315
rect 1265 -6350 1270 -6320
rect 1300 -6350 1305 -6320
rect 1265 -6355 1305 -6350
rect 1275 -6575 1305 -6355
rect 1265 -6580 1305 -6575
rect 1265 -6610 1270 -6580
rect 1300 -6610 1305 -6580
rect 1265 -6615 1305 -6610
rect 1985 -5460 2015 0
rect 2045 -3750 2075 0
rect 2105 -2895 2135 0
rect 2165 -2040 2195 0
rect 2225 -1185 2255 0
rect 2285 -610 2315 0
rect 2285 -615 2325 -610
rect 2285 -645 2290 -615
rect 2320 -645 2325 -615
rect 2285 -650 2325 -645
rect 2225 -1190 2265 -1185
rect 2225 -1220 2230 -1190
rect 2260 -1220 2265 -1190
rect 2225 -1225 2265 -1220
rect 2225 -1445 2255 -1225
rect 2225 -1450 2265 -1445
rect 2225 -1480 2230 -1450
rect 2260 -1480 2265 -1450
rect 2225 -1485 2265 -1480
rect 2165 -2045 2205 -2040
rect 2165 -2075 2170 -2045
rect 2200 -2075 2205 -2045
rect 2165 -2080 2205 -2075
rect 2165 -2300 2195 -2080
rect 2165 -2305 2205 -2300
rect 2165 -2335 2170 -2305
rect 2200 -2335 2205 -2305
rect 2165 -2340 2205 -2335
rect 2105 -2900 2145 -2895
rect 2105 -2930 2110 -2900
rect 2140 -2930 2145 -2900
rect 2105 -2935 2145 -2930
rect 2105 -3155 2135 -2935
rect 2105 -3160 2145 -3155
rect 2105 -3190 2110 -3160
rect 2140 -3190 2145 -3160
rect 2105 -3195 2145 -3190
rect 2045 -3755 2085 -3750
rect 2045 -3785 2050 -3755
rect 2080 -3785 2085 -3755
rect 2045 -3790 2085 -3785
rect 2045 -4605 2075 -3790
rect 2045 -4610 2085 -4605
rect 2045 -4640 2050 -4610
rect 2080 -4640 2085 -4610
rect 2045 -4645 2085 -4640
rect 2045 -4865 2075 -4645
rect 2045 -4870 2085 -4865
rect 2045 -4900 2050 -4870
rect 2080 -4900 2085 -4870
rect 2045 -4905 2085 -4900
rect 1985 -5465 2025 -5460
rect 1985 -5495 1990 -5465
rect 2020 -5495 2025 -5465
rect 1985 -5500 2025 -5495
rect 1985 -6315 2015 -5500
rect 1985 -6320 2025 -6315
rect 1985 -6350 1990 -6320
rect 2020 -6350 2025 -6320
rect 1985 -6355 2025 -6350
rect 1985 -6575 2015 -6355
rect 1985 -6580 2025 -6575
rect 1985 -6610 1990 -6580
rect 2020 -6610 2025 -6580
rect 1985 -6615 2025 -6610
<< metal4 >>
rect 1205 -4715 1245 -4685
use 8_cap_array_final  8_cap_array_final_0
timestamp 1730665161
transform 0 1 115 -1 0 -65
box -65 -115 6775 2245
use mid_2_low  mid_2_low_0
timestamp 1730665161
transform 1 0 2495 0 1 0
box 0 -6840 2405 0
use mid_2_up_left  mid_2_up_left_0
timestamp 1730665161
transform 1 0 110 0 1 60
box -110 -60 2250 6780
use mid_2_up_left  mid_2_up_left_1
timestamp 1730665161
transform 1 0 2605 0 1 60
box -110 -60 2250 6780
<< end >>
