magic
tech sky130A
timestamp 1730665161
<< metal1 >>
rect 820 -60 835 6780
rect 880 2285 895 6780
rect 940 3135 955 6780
rect 1000 3135 1015 6780
rect 1060 4850 1075 6780
rect 1180 6450 1195 6555
rect 1875 6295 1890 6450
rect 1165 6290 1195 6295
rect 1165 6255 1195 6260
rect 1875 6290 1905 6295
rect 1875 6255 1905 6260
rect 1180 5515 1195 5595
rect 1180 5440 1195 5485
rect 1165 5435 1195 5440
rect 1875 5445 1890 5600
rect 1875 5440 1905 5445
rect 1875 5405 1905 5410
rect 1165 5400 1195 5405
rect 1180 5300 1195 5400
rect 1120 4660 1135 5070
rect 1120 4585 1135 4630
rect 1105 4580 1135 4585
rect 1935 4590 1950 4850
rect 1935 4585 1965 4590
rect 1935 4550 1965 4555
rect 1105 4545 1135 4550
rect 1120 3805 1135 4545
rect 1120 3730 1135 3775
rect 1105 3725 1135 3730
rect 1105 3690 1135 3695
rect 1935 3730 1950 3885
rect 1935 3725 1965 3730
rect 1935 3690 1965 3695
rect 1120 3590 1135 3690
rect 1060 2950 1075 3135
rect 1060 2875 1075 2920
rect 1045 2870 1075 2875
rect 1045 2835 1075 2840
rect 1995 2875 2010 3135
rect 1995 2870 2025 2875
rect 1995 2835 2025 2840
rect 1060 2735 1075 2835
rect 1000 2095 1015 2280
rect 1000 2020 1015 2065
rect 985 2015 1015 2020
rect 985 1980 1015 1985
rect 2055 2020 2070 2280
rect 2055 2015 2085 2020
rect 2055 1980 2085 1985
rect 1000 1880 1015 1980
rect 940 1240 955 1425
rect 940 1165 955 1210
rect 925 1160 955 1165
rect 925 1125 955 1130
rect 2115 1165 2130 1425
rect 2115 1160 2145 1165
rect 2115 1125 2145 1130
rect 940 1025 955 1125
rect 880 385 895 570
rect 880 310 895 355
rect 865 305 895 310
rect 865 270 895 275
rect 2175 310 2190 570
rect 2175 305 2205 310
rect 2175 270 2205 275
rect 880 170 895 270
rect 2235 -60 2250 -20
<< via1 >>
rect 1165 6260 1195 6290
rect 1875 6260 1905 6290
rect 1165 5405 1195 5435
rect 1875 5410 1905 5440
rect 1105 4550 1135 4580
rect 1935 4555 1965 4585
rect 1105 3695 1135 3725
rect 1935 3695 1965 3725
rect 1045 2840 1075 2870
rect 1995 2840 2025 2870
rect 985 1985 1015 2015
rect 2055 1985 2085 2015
rect 925 1130 955 1160
rect 2115 1130 2145 1160
rect 865 275 895 305
rect 2175 275 2205 305
<< metal2 >>
rect 820 -60 835 6780
rect 880 465 895 6780
rect 940 1320 955 6780
rect 1000 2175 1015 6780
rect 1060 3030 1075 6780
rect 1120 4740 1135 6780
rect 1180 6450 1195 6780
rect 1875 6555 1890 6780
rect 1875 6550 1915 6555
rect 1875 6520 1880 6550
rect 1910 6520 1915 6550
rect 1875 6515 1915 6520
rect 1155 6445 1195 6450
rect 1155 6415 1160 6445
rect 1190 6440 1195 6445
rect 1875 6445 1915 6450
rect 1875 6440 1880 6445
rect 1190 6425 1200 6440
rect 1870 6425 1880 6440
rect 1190 6415 1195 6425
rect 1155 6410 1195 6415
rect 1875 6415 1880 6425
rect 1910 6415 1915 6445
rect 1875 6410 1915 6415
rect 1165 6290 1195 6295
rect 1875 6290 1905 6295
rect 1195 6270 1200 6285
rect 1860 6270 1875 6285
rect 1165 6255 1195 6260
rect 1875 6255 1905 6260
rect 1875 5595 1915 5600
rect 1155 5590 1195 5595
rect 1155 5560 1160 5590
rect 1190 5585 1195 5590
rect 1875 5585 1880 5595
rect 1190 5570 1200 5585
rect 1870 5570 1880 5585
rect 1190 5560 1195 5570
rect 1875 5565 1880 5570
rect 1910 5565 1915 5595
rect 1875 5560 1915 5565
rect 1155 5555 1195 5560
rect 1875 5440 1905 5445
rect 1165 5435 1195 5440
rect 1195 5415 1200 5430
rect 1870 5415 1875 5430
rect 1875 5405 1905 5410
rect 1165 5400 1195 5405
rect 1095 4735 1135 4740
rect 1095 4705 1100 4735
rect 1130 4730 1135 4735
rect 1935 4745 1950 6780
rect 1935 4740 1975 4745
rect 1935 4730 1940 4740
rect 1130 4715 1200 4730
rect 1865 4715 1940 4730
rect 1130 4705 1135 4715
rect 1935 4710 1940 4715
rect 1970 4710 1975 4740
rect 1935 4705 1975 4710
rect 1095 4700 1135 4705
rect 1935 4585 1965 4590
rect 1105 4580 1135 4585
rect 1135 4560 1200 4575
rect 1870 4560 1935 4575
rect 1935 4550 1965 4555
rect 1105 4545 1135 4550
rect 1095 3880 1135 3885
rect 1095 3850 1100 3880
rect 1130 3875 1135 3880
rect 1935 3880 1975 3885
rect 1935 3875 1940 3880
rect 1130 3860 1200 3875
rect 1870 3860 1940 3875
rect 1130 3850 1135 3860
rect 1095 3845 1135 3850
rect 1935 3850 1940 3860
rect 1970 3850 1975 3880
rect 1935 3845 1975 3850
rect 1105 3725 1135 3730
rect 1935 3725 1965 3730
rect 1135 3705 1200 3720
rect 1870 3705 1935 3720
rect 1105 3690 1135 3695
rect 1935 3690 1965 3695
rect 1035 3025 1075 3030
rect 1035 2995 1040 3025
rect 1070 3020 1075 3025
rect 1995 3030 2010 6780
rect 1995 3025 2035 3030
rect 1995 3020 2000 3025
rect 1070 3005 1200 3020
rect 1870 3005 2000 3020
rect 1070 2995 1075 3005
rect 1035 2990 1075 2995
rect 1995 2995 2000 3005
rect 2030 2995 2035 3025
rect 1995 2990 2035 2995
rect 1045 2870 1075 2875
rect 1995 2870 2025 2875
rect 1075 2850 1200 2865
rect 1870 2850 1995 2865
rect 1045 2835 1075 2840
rect 1995 2835 2025 2840
rect 975 2170 1015 2175
rect 975 2140 980 2170
rect 1010 2165 1015 2170
rect 2055 2175 2070 6780
rect 2055 2170 2095 2175
rect 2055 2165 2060 2170
rect 1010 2150 1200 2165
rect 1870 2150 2060 2165
rect 1010 2140 1015 2150
rect 975 2135 1015 2140
rect 2055 2140 2060 2150
rect 2090 2140 2095 2170
rect 2055 2135 2095 2140
rect 985 2015 1015 2020
rect 2055 2015 2085 2020
rect 1015 1995 1200 2010
rect 1870 1995 2055 2010
rect 985 1980 1015 1985
rect 2055 1980 2085 1985
rect 915 1315 955 1320
rect 915 1285 920 1315
rect 950 1310 955 1315
rect 2115 1320 2130 6780
rect 2115 1315 2155 1320
rect 2115 1310 2120 1315
rect 950 1295 1200 1310
rect 1870 1295 2120 1310
rect 950 1285 955 1295
rect 915 1280 955 1285
rect 2115 1285 2120 1295
rect 2150 1285 2155 1315
rect 2115 1280 2155 1285
rect 925 1160 955 1165
rect 2115 1160 2145 1165
rect 955 1140 1200 1155
rect 1870 1140 2115 1155
rect 925 1125 955 1130
rect 2115 1125 2145 1130
rect 855 460 895 465
rect 855 430 860 460
rect 890 455 895 460
rect 2175 465 2190 6780
rect 2175 460 2215 465
rect 2175 455 2180 460
rect 890 440 1200 455
rect 1870 440 2180 455
rect 890 430 895 440
rect 855 425 895 430
rect 2175 430 2180 440
rect 2210 430 2215 460
rect 2175 425 2215 430
rect 865 305 895 310
rect 2175 305 2205 310
rect 895 285 1200 300
rect 1870 285 2175 300
rect 865 270 895 275
rect 2175 270 2205 275
rect 2235 -60 2250 6780
<< via2 >>
rect 1880 6520 1910 6550
rect 1160 6415 1190 6445
rect 1880 6415 1910 6445
rect 1160 5560 1190 5590
rect 1880 5565 1910 5595
rect 1100 4705 1130 4735
rect 1940 4710 1970 4740
rect 1100 3850 1130 3880
rect 1940 3850 1970 3880
rect 1040 2995 1070 3025
rect 2000 2995 2030 3025
rect 980 2140 1010 2170
rect 2060 2140 2090 2170
rect 920 1285 950 1315
rect 2120 1285 2150 1315
rect 860 430 890 460
rect 2180 430 2210 460
<< metal3 >>
rect 1875 6550 1915 6555
rect 1875 6520 1880 6550
rect 1910 6520 1915 6550
rect 1875 6515 1915 6520
rect 1875 6450 1905 6515
rect 1155 6445 1195 6450
rect 1155 6415 1160 6445
rect 1190 6415 1195 6445
rect 1155 6410 1195 6415
rect 1165 5595 1195 6410
rect 1155 5590 1195 5595
rect 1155 5560 1160 5590
rect 1190 5560 1195 5590
rect 1155 5555 1195 5560
rect 1095 4735 1135 4740
rect 1095 4705 1100 4735
rect 1130 4705 1135 4735
rect 1095 4700 1135 4705
rect 1105 3885 1135 4700
rect 1095 3880 1135 3885
rect 1095 3850 1100 3880
rect 1130 3850 1135 3880
rect 1095 3845 1135 3850
rect 1035 3025 1075 3030
rect 1035 2995 1040 3025
rect 1070 2995 1075 3025
rect 1035 2990 1075 2995
rect 975 2170 1015 2175
rect 975 2140 980 2170
rect 1010 2140 1015 2170
rect 975 2135 1015 2140
rect 915 1315 955 1320
rect 915 1285 920 1315
rect 950 1285 955 1315
rect 915 1280 955 1285
rect 855 460 895 465
rect 855 430 860 460
rect 890 430 895 460
rect 855 425 895 430
rect 865 -60 895 425
rect 925 -60 955 1280
rect 985 -60 1015 2135
rect 1045 -60 1075 2990
rect 1105 -60 1135 3845
rect 1165 -60 1195 5555
rect 1875 6445 1915 6450
rect 1875 6415 1880 6445
rect 1910 6415 1915 6445
rect 1875 6410 1915 6415
rect 1875 5600 1905 6410
rect 1875 5595 1915 5600
rect 1875 5565 1880 5595
rect 1910 5565 1915 5595
rect 1875 5560 1915 5565
rect 1875 -60 1905 5560
rect 1935 4740 1975 4745
rect 1935 4710 1940 4740
rect 1970 4710 1975 4740
rect 1935 4705 1975 4710
rect 1935 3885 1965 4705
rect 1935 3880 1975 3885
rect 1935 3850 1940 3880
rect 1970 3850 1975 3880
rect 1935 3845 1975 3850
rect 1935 -60 1965 3845
rect 1995 3025 2035 3030
rect 1995 2995 2000 3025
rect 2030 2995 2035 3025
rect 1995 2990 2035 2995
rect 1995 -60 2025 2990
rect 2055 2170 2095 2175
rect 2055 2140 2060 2170
rect 2090 2140 2095 2170
rect 2055 2135 2095 2140
rect 2055 -60 2085 2135
rect 2115 1315 2155 1320
rect 2115 1285 2120 1315
rect 2150 1285 2155 1315
rect 2115 1280 2155 1285
rect 2115 -60 2145 1280
rect 2175 460 2215 465
rect 2175 430 2180 460
rect 2210 430 2215 460
rect 2175 425 2215 430
rect 2175 -60 2205 425
use 8_cap_array_final  8_cap_array_final_1
timestamp 1730665161
transform 0 1 5 -1 0 6715
box -65 -115 6775 2245
<< end >>
