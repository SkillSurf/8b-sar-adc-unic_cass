magic
tech sky130A
magscale 1 2
timestamp 1728842282
<< pwell >>
rect 1140 -930 1160 -890
rect 1520 -950 1850 -880
<< locali >>
rect 710 180 1520 200
rect 710 140 840 180
rect 1080 140 1160 180
rect 1400 140 1520 180
rect 710 110 1520 140
rect 710 -890 1520 -860
rect 710 -930 840 -890
rect 1080 -930 1140 -890
rect 1400 -930 1520 -890
rect 710 -950 1520 -930
<< viali >>
rect 840 140 1080 180
rect 1160 140 1400 180
rect 840 -930 1080 -890
rect 1140 -930 1400 -890
<< metal1 >>
rect 370 530 1850 540
rect 370 510 840 530
rect 830 470 840 510
rect 900 510 1850 530
rect 900 470 910 510
rect 830 460 910 470
rect 1330 470 1410 480
rect 1330 430 1340 470
rect 370 410 1340 430
rect 1400 430 1410 470
rect 1400 410 1850 430
rect 370 400 1850 410
rect 370 360 1850 370
rect 370 340 1250 360
rect 920 300 1000 310
rect 920 260 930 300
rect 370 240 930 260
rect 990 260 1000 300
rect 1240 300 1250 340
rect 1310 340 1850 360
rect 1310 300 1320 340
rect 1240 290 1320 300
rect 990 240 1850 260
rect 370 230 1850 240
rect 370 180 1850 200
rect 370 140 840 180
rect 1080 140 1160 180
rect 1400 140 1850 180
rect 370 130 1850 140
rect 910 70 1010 80
rect 910 10 930 70
rect 990 10 1010 70
rect 910 0 1010 10
rect 1220 70 1320 80
rect 1220 10 1240 70
rect 1300 10 1320 70
rect 1220 0 1320 10
rect 900 -340 930 -220
rect 850 -350 930 -340
rect 850 -410 860 -350
rect 920 -410 930 -350
rect 850 -420 930 -410
rect 900 -540 930 -420
rect 990 -340 1020 -220
rect 1210 -340 1240 -220
rect 990 -350 1240 -340
rect 990 -410 1030 -350
rect 1090 -410 1140 -350
rect 1200 -410 1240 -350
rect 990 -420 1240 -410
rect 990 -540 1020 -420
rect 1210 -540 1240 -420
rect 1300 -340 1330 -220
rect 1300 -350 1380 -340
rect 1300 -410 1310 -350
rect 1370 -410 1380 -350
rect 1300 -420 1380 -410
rect 1300 -540 1330 -420
rect 910 -770 1010 -760
rect 910 -830 930 -770
rect 990 -830 1010 -770
rect 910 -840 1010 -830
rect 1220 -770 1320 -760
rect 1220 -830 1240 -770
rect 1300 -830 1320 -770
rect 1220 -840 1320 -830
rect 370 -890 1850 -880
rect 370 -930 840 -890
rect 1080 -930 1140 -890
rect 1400 -930 1850 -890
rect 370 -950 1850 -930
rect 370 -990 1850 -980
rect 370 -1010 940 -990
rect 930 -1050 940 -1010
rect 1000 -1010 1850 -990
rect 1000 -1050 1010 -1010
rect 1240 -1090 1250 -1060
rect 370 -1120 1250 -1090
rect 1310 -1090 1320 -1060
rect 1310 -1120 1850 -1090
rect 370 -3170 1850 -3150
rect 370 -3190 470 -3170
rect 450 -3230 470 -3190
rect 530 -3190 1850 -3170
rect 530 -3230 550 -3190
rect 450 -3250 550 -3230
<< via1 >>
rect 840 470 900 530
rect 1340 410 1400 470
rect 930 240 990 300
rect 1250 300 1310 360
rect 930 10 990 70
rect 1240 10 1300 70
rect 860 -410 920 -350
rect 1030 -410 1090 -350
rect 1140 -410 1200 -350
rect 1310 -410 1370 -350
rect 930 -830 990 -770
rect 1240 -830 1300 -770
rect 940 -1050 1000 -990
rect 1250 -1120 1310 -1060
rect 470 -3230 530 -3170
<< metal2 >>
rect 830 530 910 540
rect 830 470 840 530
rect 900 470 910 530
rect 830 460 910 470
rect 1330 470 1410 480
rect 850 -340 880 460
rect 1330 410 1340 470
rect 1400 410 1410 470
rect 1330 400 1410 410
rect 1240 360 1320 370
rect 920 300 1000 310
rect 920 240 930 300
rect 990 240 1000 300
rect 1240 300 1250 360
rect 1310 300 1320 360
rect 1240 290 1320 300
rect 920 230 1000 240
rect 950 80 980 230
rect 1260 80 1290 290
rect 920 70 1000 80
rect 920 10 930 70
rect 990 10 1000 70
rect 920 0 1000 10
rect 1230 70 1310 80
rect 1230 10 1240 70
rect 1300 10 1310 70
rect 1230 0 1310 10
rect 1350 -340 1380 400
rect 850 -350 930 -340
rect 850 -410 860 -350
rect 920 -410 930 -350
rect 850 -420 930 -410
rect 1020 -350 1210 -340
rect 1020 -410 1030 -350
rect 1090 -410 1140 -350
rect 1200 -410 1210 -350
rect 1020 -420 1210 -410
rect 1300 -350 1380 -340
rect 1300 -410 1310 -350
rect 1370 -410 1380 -350
rect 1300 -420 1380 -410
rect 920 -770 1000 -760
rect 920 -830 930 -770
rect 990 -830 1000 -770
rect 920 -840 1000 -830
rect 950 -980 980 -840
rect 1100 -960 1130 -420
rect 1230 -770 1310 -760
rect 1230 -830 1240 -770
rect 1300 -830 1310 -770
rect 1230 -840 1310 -830
rect 1060 -970 1170 -960
rect 930 -990 1010 -980
rect 930 -1050 940 -990
rect 1000 -1050 1010 -990
rect 1060 -1050 1070 -970
rect 1160 -1050 1170 -970
rect 1060 -1060 1170 -1050
rect 1260 -1060 1290 -840
rect 1240 -1120 1250 -1060
rect 1310 -1120 1320 -1060
rect 450 -3170 550 -3150
rect 450 -3230 470 -3170
rect 530 -3230 550 -3170
rect 450 -3250 550 -3230
<< via2 >>
rect 1070 -1050 1160 -970
rect 470 -3230 530 -3170
<< metal3 >>
rect 1060 -970 1170 -960
rect 1060 -1050 1070 -970
rect 1160 -1050 1170 -970
rect 1060 -1060 1170 -1050
rect 450 -3160 550 -3150
rect 450 -3240 460 -3160
rect 540 -3240 550 -3160
rect 450 -3250 550 -3240
<< via3 >>
rect 1070 -1050 1160 -970
rect 460 -3170 540 -3160
rect 460 -3230 470 -3170
rect 470 -3230 530 -3170
rect 530 -3230 540 -3170
rect 460 -3240 540 -3230
<< metal4 >>
rect 1060 -970 1170 -960
rect 1060 -1050 1070 -970
rect 1160 -1050 1170 -970
rect 1060 -1160 1170 -1050
rect 450 -3160 550 -2840
rect 450 -3240 460 -3160
rect 540 -3240 550 -3160
rect 450 -3250 550 -3240
use sky130_fd_pr__cap_mim_m3_1_BZXSER  sky130_fd_pr__cap_mim_m3_1_BZXSER_0
timestamp 1728836072
transform 0 -1 1110 1 0 -2034
box -886 -740 886 740
use sky130_fd_pr__nfet_01v8_5WU4M2  sky130_fd_pr__nfet_01v8_5WU4M2_0
timestamp 1728804544
transform -1 0 1271 0 -1 -661
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_QKK3FL  sky130_fd_pr__pfet_01v8_QKK3FL_0
timestamp 1728804544
transform -1 0 1271 0 -1 -96
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_NKK3FE  XM1
timestamp 1728804544
transform 1 0 961 0 1 -96
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_5WP7M2  XM2
timestamp 1728804544
transform 1 0 961 0 1 -661
box -211 -279 211 279
<< labels >>
flabel metal1 770 -940 830 -880 0 FreeSans 256 0 0 0 sub
port 6 nsew
flabel metal1 1080 -940 1140 -880 0 FreeSans 256 0 0 0 sub
port 1 nsew
flabel via1 840 470 900 530 0 FreeSans 256 0 0 0 Vin
port 5 nsew
flabel via1 1340 410 1400 470 0 FreeSans 256 0 0 0 GND
port 9 nsew
flabel via1 930 240 990 300 0 FreeSans 256 0 0 0 phi1_n
port 4 nsew
flabel via1 1250 300 1310 360 0 FreeSans 256 0 0 0 phi2_n
port 10 nsew
flabel via1 1250 -1120 1310 -1060 0 FreeSans 256 0 0 0 phi2
port 8 nsew
flabel via1 940 -1050 1000 -990 0 FreeSans 256 0 0 0 phi1
port 2 nsew
flabel metal1 770 130 830 190 0 FreeSans 256 0 0 0 Vdd
port 3 nsew
flabel metal1 1100 130 1150 190 0 FreeSans 256 0 0 0 Vdd
port 7 nsew
flabel via1 470 -3230 530 -3170 0 FreeSans 256 0 0 0 com_x
port 0 nsew
<< end >>
