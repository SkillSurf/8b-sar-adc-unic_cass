magic
tech sky130A
timestamp 1730649634
<< pwell >>
rect -3185 14950 -3150 14995
<< metal1 >>
rect 2075 16310 2080 16325
rect -2570 16295 2080 16310
rect 2110 16310 2115 16325
rect 4570 16310 4575 16325
rect 2110 16295 4575 16310
rect 4605 16310 4610 16325
rect 7065 16310 7070 16325
rect 4605 16295 7070 16310
rect 7100 16310 7105 16325
rect 9560 16310 9565 16325
rect 7100 16295 9565 16310
rect 9595 16310 9600 16325
rect 12055 16310 12060 16325
rect 9595 16295 12060 16310
rect 12090 16310 12095 16325
rect 14550 16310 14555 16325
rect 12090 16295 14555 16310
rect 14585 16310 14590 16325
rect 17045 16310 17050 16325
rect 14585 16295 17050 16310
rect 17080 16310 17085 16325
rect 19540 16310 19545 16325
rect 17080 16295 19545 16310
rect 19575 16310 19580 16325
rect 22035 16310 22040 16325
rect 19575 16295 22040 16310
rect 22070 16310 22075 16325
rect 24530 16310 24535 16325
rect 22070 16295 24535 16310
rect 24565 16310 24570 16325
rect 27025 16310 27030 16325
rect 24565 16295 27030 16310
rect 27060 16310 27065 16325
rect 29520 16310 29525 16325
rect 27060 16295 29525 16310
rect 29555 16310 29560 16325
rect 32015 16310 32020 16325
rect 29555 16295 32020 16310
rect 32050 16310 32055 16325
rect 34510 16310 34515 16325
rect 32050 16295 34515 16310
rect 34545 16310 34550 16325
rect 37005 16310 37010 16325
rect 34545 16295 37010 16310
rect 37040 16310 37045 16325
rect 39500 16310 39505 16325
rect 37040 16295 39505 16310
rect 39535 16310 39540 16325
rect 39535 16295 42325 16310
rect 1210 16240 1240 16260
rect 2045 16240 2050 16255
rect -2570 16225 2050 16240
rect 2080 16240 2085 16255
rect 3705 16240 3735 16260
rect 4540 16240 4545 16255
rect 2080 16225 4545 16240
rect 4575 16240 4580 16255
rect 6200 16240 6230 16260
rect 7035 16240 7040 16255
rect 4575 16225 7040 16240
rect 7070 16240 7075 16255
rect 8695 16240 8725 16260
rect 9530 16240 9535 16255
rect 7070 16225 9535 16240
rect 9565 16240 9570 16255
rect 11190 16240 11220 16260
rect 12025 16240 12030 16255
rect 9565 16225 12030 16240
rect 12060 16240 12065 16255
rect 13685 16240 13715 16260
rect 14520 16240 14525 16255
rect 12060 16225 14525 16240
rect 14555 16240 14560 16255
rect 16180 16240 16210 16260
rect 17015 16240 17020 16255
rect 14555 16225 17020 16240
rect 17050 16240 17055 16255
rect 18675 16240 18705 16260
rect 19510 16240 19515 16255
rect 17050 16225 19515 16240
rect 19545 16240 19550 16255
rect 21170 16240 21200 16260
rect 22005 16240 22010 16255
rect 19545 16225 22010 16240
rect 22040 16240 22045 16255
rect 23665 16240 23695 16260
rect 24500 16240 24505 16255
rect 22040 16225 24505 16240
rect 24535 16240 24540 16255
rect 26160 16240 26190 16260
rect 26995 16240 27000 16255
rect 24535 16225 27000 16240
rect 27030 16240 27035 16255
rect 28655 16240 28685 16260
rect 29490 16240 29495 16255
rect 27030 16225 29495 16240
rect 29525 16240 29530 16255
rect 31150 16240 31180 16260
rect 31985 16240 31990 16255
rect 29525 16225 31990 16240
rect 32020 16240 32025 16255
rect 33645 16240 33675 16260
rect 34480 16240 34485 16255
rect 32020 16225 34485 16240
rect 34515 16240 34520 16255
rect 36140 16240 36170 16260
rect 36975 16240 36980 16255
rect 34515 16225 36980 16240
rect 37010 16240 37015 16255
rect 38635 16240 38665 16260
rect 39470 16240 39475 16255
rect 37010 16225 39475 16240
rect 39505 16240 39510 16255
rect 39505 16225 42325 16240
rect 7155 16170 7160 16185
rect -2570 16155 7160 16170
rect 7190 16170 7195 16185
rect 9650 16170 9655 16185
rect 7190 16155 9655 16170
rect 9685 16170 9690 16185
rect 12145 16170 12150 16185
rect 9685 16155 12150 16170
rect 12180 16170 12185 16185
rect 14640 16170 14645 16185
rect 12180 16155 14645 16170
rect 14675 16170 14680 16185
rect 17135 16170 17140 16185
rect 14675 16155 17140 16170
rect 17170 16170 17175 16185
rect 19630 16170 19635 16185
rect 17170 16155 19635 16170
rect 19665 16170 19670 16185
rect 22125 16170 22130 16185
rect 19665 16155 22130 16170
rect 22160 16170 22165 16185
rect 24620 16170 24625 16185
rect 22160 16155 24625 16170
rect 24655 16170 24660 16185
rect 27115 16170 27120 16185
rect 24655 16155 27120 16170
rect 27150 16170 27155 16185
rect 29610 16170 29615 16185
rect 27150 16155 29615 16170
rect 29645 16170 29650 16185
rect 32105 16170 32110 16185
rect 29645 16155 32110 16170
rect 32140 16170 32145 16185
rect 34600 16170 34605 16185
rect 32140 16155 34605 16170
rect 34635 16170 34640 16185
rect 34635 16155 42325 16170
rect 6110 16100 6140 16120
rect 7125 16100 7130 16115
rect -2570 16085 7130 16100
rect 7160 16100 7165 16115
rect 8605 16100 8635 16120
rect 9620 16100 9625 16115
rect 7160 16085 9625 16100
rect 9655 16100 9660 16115
rect 11100 16100 11130 16120
rect 12115 16100 12120 16115
rect 9655 16085 12120 16100
rect 12150 16100 12155 16115
rect 13595 16100 13625 16120
rect 14610 16100 14615 16115
rect 12150 16085 14615 16100
rect 14645 16100 14650 16115
rect 16090 16100 16120 16120
rect 17105 16100 17110 16115
rect 14645 16085 17110 16100
rect 17140 16100 17145 16115
rect 18585 16100 18615 16120
rect 19600 16100 19605 16115
rect 17140 16085 19605 16100
rect 19635 16100 19640 16115
rect 21080 16100 21110 16120
rect 22095 16100 22100 16115
rect 19635 16085 22100 16100
rect 22130 16100 22135 16115
rect 23575 16100 23605 16120
rect 24590 16100 24595 16115
rect 22130 16085 24595 16100
rect 24625 16100 24630 16115
rect 26070 16100 26100 16120
rect 27085 16100 27090 16115
rect 24625 16085 27090 16100
rect 27120 16100 27125 16115
rect 28565 16100 28595 16120
rect 29580 16100 29585 16115
rect 27120 16085 29585 16100
rect 29615 16100 29620 16115
rect 31060 16100 31090 16120
rect 32075 16100 32080 16115
rect 29615 16085 32080 16100
rect 32110 16100 32115 16115
rect 33555 16100 33585 16120
rect 34570 16100 34575 16115
rect 32110 16085 34575 16100
rect 34605 16100 34610 16115
rect 34605 16085 42325 16100
rect 12325 16030 12330 16045
rect -2570 16015 12330 16030
rect 12360 16030 12365 16045
rect 14820 16030 14825 16045
rect 12360 16015 14825 16030
rect 14855 16030 14860 16045
rect 17225 16030 17230 16045
rect 14855 16015 17230 16030
rect 17260 16030 17265 16045
rect 19720 16030 19725 16045
rect 17260 16015 19725 16030
rect 19755 16030 19760 16045
rect 22215 16030 22220 16045
rect 19755 16015 22220 16030
rect 22250 16030 22255 16045
rect 24710 16030 24715 16045
rect 22250 16015 24715 16030
rect 24745 16030 24750 16045
rect 27295 16030 27300 16045
rect 24745 16015 27300 16030
rect 27330 16030 27335 16045
rect 29790 16030 29795 16045
rect 27330 16015 29795 16030
rect 29825 16030 29830 16045
rect 29825 16015 42325 16030
rect 10920 15960 10950 15980
rect 12295 15960 12300 15975
rect -2570 15945 12300 15960
rect 12330 15960 12335 15975
rect 13415 15960 13445 15980
rect 14790 15960 14795 15975
rect 12330 15945 14795 15960
rect 14825 15960 14830 15975
rect 16000 15960 16030 15980
rect 17195 15960 17200 15975
rect 14825 15945 17200 15960
rect 17230 15960 17235 15975
rect 18495 15960 18525 15980
rect 19690 15960 19695 15975
rect 17230 15945 19695 15960
rect 19725 15960 19730 15975
rect 20990 15960 21020 15980
rect 22185 15960 22190 15975
rect 19725 15945 22190 15960
rect 22220 15960 22225 15975
rect 23485 15960 23515 15980
rect 24680 15960 24685 15975
rect 22220 15945 24685 15960
rect 24715 15960 24720 15975
rect 25890 15960 25920 15980
rect 27265 15960 27270 15975
rect 24715 15945 27270 15960
rect 27300 15960 27305 15975
rect 28385 15960 28415 15980
rect 29760 15960 29765 15975
rect 27300 15945 29765 15960
rect 29795 15960 29800 15975
rect 29795 15945 42325 15960
rect 12235 15890 12240 15905
rect -2570 15875 12240 15890
rect 12270 15890 12275 15905
rect 14730 15890 14735 15905
rect 12270 15875 14735 15890
rect 14765 15890 14770 15905
rect 17315 15890 17320 15905
rect 14765 15875 17320 15890
rect 17350 15890 17355 15905
rect 19810 15890 19815 15905
rect 17350 15875 19815 15890
rect 19845 15890 19850 15905
rect 22305 15890 22310 15905
rect 19845 15875 22310 15890
rect 22340 15890 22345 15905
rect 24800 15890 24805 15905
rect 22340 15875 24805 15890
rect 24835 15890 24840 15905
rect 27205 15890 27210 15905
rect 24835 15875 27210 15890
rect 27240 15890 27245 15905
rect 29700 15890 29705 15905
rect 27240 15875 29705 15890
rect 29735 15890 29740 15905
rect 29735 15875 42325 15890
rect 11010 15820 11040 15840
rect 12205 15820 12210 15835
rect -2570 15805 12210 15820
rect 12240 15820 12245 15835
rect 13505 15820 13535 15840
rect 14700 15820 14705 15835
rect 12240 15805 14705 15820
rect 14735 15820 14740 15835
rect 15910 15820 15940 15840
rect 17285 15820 17290 15835
rect 14735 15805 17290 15820
rect 17320 15820 17325 15835
rect 18405 15820 18435 15840
rect 19780 15820 19785 15835
rect 17320 15805 19785 15820
rect 19815 15820 19820 15835
rect 20900 15820 20930 15840
rect 22275 15820 22280 15835
rect 19815 15805 22280 15820
rect 22310 15820 22315 15835
rect 23395 15820 23425 15840
rect 24770 15820 24775 15835
rect 22310 15805 24775 15820
rect 24805 15820 24810 15835
rect 25980 15820 26010 15840
rect 27175 15820 27180 15835
rect 24805 15805 27180 15820
rect 27210 15820 27215 15835
rect 28475 15820 28505 15840
rect 29670 15820 29675 15835
rect 27210 15805 29675 15820
rect 29705 15820 29710 15835
rect 29705 15805 42325 15820
rect 17495 15750 17500 15765
rect -2570 15735 17500 15750
rect 17530 15750 17535 15765
rect 19900 15750 19905 15765
rect 17530 15735 19905 15750
rect 19935 15750 19940 15765
rect 22395 15750 22400 15765
rect 19935 15735 22400 15750
rect 22430 15750 22435 15765
rect 24980 15750 24985 15765
rect 22430 15735 24985 15750
rect 25015 15750 25020 15765
rect 25015 15735 42325 15750
rect 15730 15680 15760 15700
rect 17465 15680 17470 15695
rect -2570 15665 17470 15680
rect 17500 15680 17505 15695
rect 18315 15680 18345 15700
rect 19870 15680 19875 15695
rect 17500 15665 19875 15680
rect 19905 15680 19910 15695
rect 20810 15680 20840 15700
rect 22365 15680 22370 15695
rect 19905 15665 22370 15680
rect 22400 15680 22405 15695
rect 23215 15680 23245 15700
rect 24950 15680 24955 15695
rect 22400 15665 24955 15680
rect 24985 15680 24990 15695
rect 24985 15665 42325 15680
rect 17405 15610 17410 15625
rect -2570 15595 17410 15610
rect 17440 15610 17445 15625
rect 24890 15610 24895 15625
rect 17440 15595 24895 15610
rect 24925 15610 24930 15625
rect 24925 15595 42325 15610
rect 15820 15540 15850 15560
rect 17375 15540 17380 15555
rect -2570 15525 17380 15540
rect 17410 15540 17415 15555
rect 23305 15540 23335 15560
rect 24860 15540 24865 15555
rect 17410 15525 24865 15540
rect 24895 15540 24900 15555
rect 24895 15525 42325 15540
rect 19990 15470 19995 15485
rect -2570 15455 19995 15470
rect 20025 15470 20030 15485
rect 22575 15470 22580 15485
rect 20025 15455 22580 15470
rect 22610 15470 22615 15485
rect 22610 15455 42325 15470
rect 18225 15400 18255 15420
rect 19960 15400 19965 15415
rect -2570 15385 19965 15400
rect 19995 15400 20000 15415
rect 22545 15400 22550 15415
rect 19995 15385 22550 15400
rect 22580 15400 22585 15415
rect 22580 15385 42325 15400
rect 22500 15330 22505 15345
rect -2570 15315 22505 15330
rect 22535 15330 22540 15345
rect 22535 15315 42325 15330
rect 22455 15260 22460 15275
rect -2570 15245 22460 15260
rect 22490 15260 22495 15275
rect 22490 15245 42325 15260
rect 18105 15190 18135 15210
rect 20080 15190 20085 15205
rect -2590 15185 20085 15190
rect -2790 15175 20085 15185
rect 20115 15190 20120 15205
rect 20115 15175 42325 15190
rect -2790 15170 -2570 15175
rect 18135 15120 18165 15140
rect 20045 15120 20050 15135
rect -2585 15115 20050 15120
rect -2790 15105 20050 15115
rect 20080 15120 20085 15135
rect 20080 15105 42325 15120
rect -2790 15100 -2570 15105
rect -2795 14975 -2780 15070
rect -2765 15060 -2715 15070
rect -2555 15060 -2550 15090
rect -2520 15075 42325 15090
rect -2520 15060 -2515 15075
rect -2765 15030 -2755 15060
rect -2725 15045 -2715 15060
rect -430 15045 -425 15060
rect -2725 15030 -425 15045
rect -395 15045 -390 15060
rect 1930 15045 1935 15060
rect -395 15030 1935 15045
rect 1965 15045 1970 15060
rect 4425 15045 4430 15060
rect 1965 15030 4430 15045
rect 4460 15045 4465 15060
rect 6920 15045 6925 15060
rect 4460 15030 6925 15045
rect 6955 15045 6960 15060
rect 9415 15045 9420 15060
rect 6955 15030 9420 15045
rect 9450 15045 9455 15060
rect 11910 15045 11915 15060
rect 9450 15030 11915 15045
rect 11945 15045 11950 15060
rect 14405 15045 14410 15060
rect 11945 15030 14410 15045
rect 14440 15045 14445 15060
rect 16900 15045 16905 15060
rect 14440 15030 16905 15045
rect 16935 15045 16940 15060
rect 19395 15045 19400 15060
rect 16935 15030 19400 15045
rect 19430 15045 19435 15060
rect 21890 15045 21895 15060
rect 19430 15030 21895 15045
rect 21925 15045 21930 15060
rect 24385 15045 24390 15060
rect 21925 15030 24390 15045
rect 24420 15045 24425 15060
rect 26880 15045 26885 15060
rect 24420 15030 26885 15045
rect 26915 15045 26920 15060
rect 29375 15045 29380 15060
rect 26915 15030 29380 15045
rect 29410 15045 29415 15060
rect 31870 15045 31875 15060
rect 29410 15030 31875 15045
rect 31905 15045 31910 15060
rect 34365 15045 34370 15060
rect 31905 15030 34370 15045
rect 34400 15045 34405 15060
rect 36860 15045 36865 15060
rect 34400 15030 36865 15045
rect 36895 15045 36900 15060
rect 39355 15045 39360 15060
rect 36895 15030 39360 15045
rect 39390 15045 39395 15060
rect 41715 15045 41720 15060
rect 39390 15030 41720 15045
rect 41750 15045 41755 15060
rect 41750 15030 42325 15045
rect -2765 15020 -2715 15030
rect -2625 14995 -2585 15000
rect -2625 14975 -2620 14995
rect -2795 14965 -2620 14975
rect -2590 14965 -2585 14995
rect -2795 14960 -2585 14965
rect -2570 14960 42325 14975
rect -2685 14925 -2645 14930
rect -2685 14895 -2680 14925
rect -2650 14895 -2645 14925
rect -2685 14890 -2645 14895
rect -2685 14525 -2655 14890
rect -450 14615 -435 14960
rect 1175 14795 1205 14800
rect 1205 14765 1305 14775
rect 1175 14760 1305 14765
rect -605 14600 -435 14615
rect -1040 14540 -1035 14570
rect -1005 14540 -1000 14570
rect -605 14540 -590 14600
rect -505 14570 -465 14575
rect -505 14540 -500 14570
rect -470 14540 -465 14570
rect -1040 14535 -1000 14540
rect -635 14535 -585 14540
rect -505 14535 -465 14540
rect -450 14535 -435 14600
rect -420 14570 -390 14575
rect -420 14535 -390 14540
rect 1290 14535 1305 14760
rect 1855 14570 1895 14575
rect 1320 14540 1325 14570
rect 1355 14540 1360 14570
rect 1320 14535 1360 14540
rect 1855 14540 1860 14570
rect 1890 14540 1895 14570
rect 1855 14535 1895 14540
rect 1910 14535 1925 14960
rect 2085 14795 2115 14800
rect 1985 14765 2085 14775
rect 1985 14760 2115 14765
rect 3670 14795 3700 14800
rect 3700 14765 3800 14775
rect 3670 14760 3800 14765
rect 1940 14570 1970 14575
rect 1940 14535 1970 14540
rect 1985 14535 2000 14760
rect 3785 14535 3800 14760
rect 4350 14570 4390 14575
rect 3815 14540 3820 14570
rect 3850 14540 3855 14570
rect 3815 14535 3855 14540
rect 4350 14540 4355 14570
rect 4385 14540 4390 14570
rect 4350 14535 4390 14540
rect 4405 14535 4420 14960
rect 4580 14795 4610 14800
rect 4480 14765 4580 14775
rect 6165 14795 6195 14800
rect 4480 14760 4610 14765
rect 6075 14765 6105 14770
rect 4435 14570 4465 14575
rect 4435 14535 4465 14540
rect 4480 14535 4495 14760
rect 6195 14765 6295 14775
rect 6165 14760 6295 14765
rect 6105 14735 6235 14745
rect 6075 14730 6235 14735
rect 6220 14535 6235 14730
rect 6280 14535 6295 14760
rect 6845 14570 6885 14575
rect 6310 14540 6315 14570
rect 6345 14540 6350 14570
rect 6310 14535 6350 14540
rect 6845 14540 6850 14570
rect 6880 14540 6885 14570
rect 6845 14535 6885 14540
rect 6900 14535 6915 14960
rect 7075 14795 7105 14800
rect 6975 14765 7075 14775
rect 8660 14795 8690 14800
rect 6975 14760 7105 14765
rect 7165 14765 7195 14770
rect 6930 14570 6960 14575
rect 6930 14535 6960 14540
rect 6975 14535 6990 14760
rect 7035 14735 7165 14745
rect 7035 14730 7195 14735
rect 8570 14765 8600 14770
rect 8690 14765 8790 14775
rect 8660 14760 8790 14765
rect 8600 14735 8730 14745
rect 8570 14730 8730 14735
rect 7035 14535 7050 14730
rect 8715 14535 8730 14730
rect 8775 14535 8790 14760
rect 9340 14570 9380 14575
rect 8805 14540 8810 14570
rect 8840 14540 8845 14570
rect 8805 14535 8845 14540
rect 9340 14540 9345 14570
rect 9375 14540 9380 14570
rect 9340 14535 9380 14540
rect 9395 14535 9410 14960
rect 9570 14795 9600 14800
rect 9470 14765 9570 14775
rect 11155 14795 11185 14800
rect 9470 14760 9600 14765
rect 9660 14765 9690 14770
rect 9425 14570 9455 14575
rect 9425 14535 9455 14540
rect 9470 14535 9485 14760
rect 9530 14735 9660 14745
rect 11065 14765 11095 14770
rect 9530 14730 9690 14735
rect 10975 14735 11005 14740
rect 9530 14535 9545 14730
rect 10885 14705 10915 14710
rect 11185 14765 11285 14775
rect 11155 14760 11285 14765
rect 11095 14735 11225 14745
rect 11065 14730 11225 14735
rect 11005 14705 11165 14715
rect 10975 14700 11165 14705
rect 10915 14675 11105 14685
rect 10885 14670 11105 14675
rect 11090 14535 11105 14670
rect 11150 14535 11165 14700
rect 11210 14535 11225 14730
rect 11270 14535 11285 14760
rect 11835 14570 11875 14575
rect 11300 14540 11305 14570
rect 11335 14540 11340 14570
rect 11300 14535 11340 14540
rect 11835 14540 11840 14570
rect 11870 14540 11875 14570
rect 11835 14535 11875 14540
rect 11890 14535 11905 14960
rect 12065 14795 12095 14800
rect 11965 14765 12065 14775
rect 13650 14795 13680 14800
rect 11965 14760 12095 14765
rect 12155 14765 12185 14770
rect 11920 14570 11950 14575
rect 11920 14535 11950 14540
rect 11965 14535 11980 14760
rect 12025 14735 12155 14745
rect 13560 14765 13590 14770
rect 12025 14730 12185 14735
rect 12245 14735 12275 14740
rect 12025 14535 12040 14730
rect 12085 14705 12245 14715
rect 13470 14735 13500 14740
rect 12085 14700 12275 14705
rect 12335 14705 12365 14710
rect 12085 14535 12100 14700
rect 12145 14675 12335 14685
rect 12145 14670 12365 14675
rect 13380 14705 13410 14710
rect 13680 14765 13780 14775
rect 13650 14760 13780 14765
rect 13590 14735 13720 14745
rect 13560 14730 13720 14735
rect 13500 14705 13660 14715
rect 13470 14700 13660 14705
rect 13410 14675 13600 14685
rect 13380 14670 13600 14675
rect 12145 14535 12160 14670
rect 13585 14535 13600 14670
rect 13645 14535 13660 14700
rect 13705 14535 13720 14730
rect 13765 14535 13780 14760
rect 14330 14570 14370 14575
rect 13795 14540 13800 14570
rect 13830 14540 13835 14570
rect 13795 14535 13835 14540
rect 14330 14540 14335 14570
rect 14365 14540 14370 14570
rect 14330 14535 14370 14540
rect 14385 14535 14400 14960
rect 14560 14795 14590 14800
rect 14460 14765 14560 14775
rect 16145 14795 16175 14800
rect 14460 14760 14590 14765
rect 14650 14765 14680 14770
rect 14415 14570 14445 14575
rect 14415 14535 14445 14540
rect 14460 14535 14475 14760
rect 14520 14735 14650 14745
rect 16055 14765 16085 14770
rect 14520 14730 14680 14735
rect 14740 14735 14770 14740
rect 14520 14535 14535 14730
rect 14580 14705 14740 14715
rect 15965 14735 15995 14740
rect 14580 14700 14770 14705
rect 14830 14705 14860 14710
rect 14580 14535 14595 14700
rect 14640 14675 14830 14685
rect 15875 14705 15905 14710
rect 14640 14670 14860 14675
rect 15785 14675 15815 14680
rect 14640 14535 14655 14670
rect 15695 14645 15725 14650
rect 16175 14765 16275 14775
rect 16145 14760 16275 14765
rect 16085 14735 16215 14745
rect 16055 14730 16215 14735
rect 15995 14705 16155 14715
rect 15965 14700 16155 14705
rect 15905 14675 16095 14685
rect 15875 14670 16095 14675
rect 15815 14645 16035 14655
rect 15785 14640 16035 14645
rect 15725 14615 15975 14625
rect 15695 14610 15975 14615
rect 15960 14535 15975 14610
rect 16020 14535 16035 14640
rect 16080 14535 16095 14670
rect 16140 14535 16155 14700
rect 16200 14535 16215 14730
rect 16260 14535 16275 14760
rect 16825 14570 16865 14575
rect 16290 14540 16295 14570
rect 16325 14540 16330 14570
rect 16290 14535 16330 14540
rect 16825 14540 16830 14570
rect 16860 14540 16865 14570
rect 16825 14535 16865 14540
rect 16880 14535 16895 14960
rect 17055 14795 17085 14800
rect 16955 14765 17055 14775
rect 18640 14795 18670 14800
rect 16955 14760 17085 14765
rect 17145 14765 17175 14770
rect 16910 14570 16940 14575
rect 16910 14535 16940 14540
rect 16955 14535 16970 14760
rect 17015 14735 17145 14745
rect 18550 14765 18580 14770
rect 17015 14730 17175 14735
rect 17235 14735 17265 14740
rect 17015 14535 17030 14730
rect 17075 14705 17235 14715
rect 18460 14735 18490 14740
rect 17075 14700 17265 14705
rect 17325 14705 17355 14710
rect 17075 14535 17090 14700
rect 17135 14675 17325 14685
rect 18370 14705 18400 14710
rect 17135 14670 17355 14675
rect 17415 14675 17445 14680
rect 17135 14535 17150 14670
rect 17195 14645 17415 14655
rect 18280 14675 18310 14680
rect 17195 14640 17445 14645
rect 17505 14645 17535 14650
rect 17195 14535 17210 14640
rect 17255 14615 17505 14625
rect 18190 14645 18220 14650
rect 17255 14610 17535 14615
rect 18100 14615 18130 14620
rect 17255 14535 17270 14610
rect 18670 14765 18770 14775
rect 18640 14760 18770 14765
rect 18580 14735 18710 14745
rect 18550 14730 18710 14735
rect 18490 14705 18650 14715
rect 18460 14700 18650 14705
rect 18400 14675 18590 14685
rect 18370 14670 18590 14675
rect 18310 14645 18530 14655
rect 18280 14640 18530 14645
rect 18220 14615 18470 14625
rect 18190 14610 18470 14615
rect 18130 14585 18410 14595
rect 18100 14580 18410 14585
rect 18395 14535 18410 14580
rect 18455 14535 18470 14610
rect 18515 14535 18530 14640
rect 18575 14535 18590 14670
rect 18635 14535 18650 14700
rect 18695 14535 18710 14730
rect 18755 14535 18770 14760
rect 19320 14570 19360 14575
rect 18785 14540 18790 14570
rect 18820 14540 18825 14570
rect 18785 14535 18825 14540
rect 19320 14540 19325 14570
rect 19355 14540 19360 14570
rect 19320 14535 19360 14540
rect 19375 14535 19390 14960
rect 19550 14795 19580 14800
rect 19450 14765 19550 14775
rect 21135 14795 21165 14800
rect 19450 14760 19580 14765
rect 19640 14765 19670 14770
rect 19405 14570 19435 14575
rect 19405 14535 19435 14540
rect 19450 14535 19465 14760
rect 19510 14735 19640 14745
rect 21045 14765 21075 14770
rect 19510 14730 19670 14735
rect 19730 14735 19760 14740
rect 19510 14535 19525 14730
rect 19570 14705 19730 14715
rect 20955 14735 20985 14740
rect 19570 14700 19760 14705
rect 19820 14705 19850 14710
rect 19570 14535 19585 14700
rect 19630 14675 19820 14685
rect 20865 14705 20895 14710
rect 19630 14670 19850 14675
rect 19910 14675 19940 14680
rect 19630 14535 19645 14670
rect 19690 14645 19910 14655
rect 20775 14675 20805 14680
rect 19690 14640 19940 14645
rect 20000 14645 20030 14650
rect 19690 14535 19705 14640
rect 19750 14615 20000 14625
rect 20685 14645 20715 14650
rect 19750 14610 20030 14615
rect 20090 14615 20120 14620
rect 19750 14535 19765 14610
rect 19810 14585 20090 14595
rect 19810 14580 20120 14585
rect 20595 14615 20625 14620
rect 21165 14765 21265 14775
rect 21135 14760 21265 14765
rect 21075 14735 21205 14745
rect 21045 14730 21205 14735
rect 20985 14705 21145 14715
rect 20955 14700 21145 14705
rect 20895 14675 21085 14685
rect 20865 14670 21085 14675
rect 20805 14645 21025 14655
rect 20775 14640 21025 14645
rect 20715 14615 20965 14625
rect 20685 14610 20965 14615
rect 20625 14585 20905 14595
rect 20595 14580 20905 14585
rect 19810 14535 19825 14580
rect 20890 14535 20905 14580
rect 20950 14535 20965 14610
rect 21010 14535 21025 14640
rect 21070 14535 21085 14670
rect 21130 14535 21145 14700
rect 21190 14535 21205 14730
rect 21250 14535 21265 14760
rect 21815 14570 21855 14575
rect 21280 14540 21285 14570
rect 21315 14540 21320 14570
rect 21280 14535 21320 14540
rect 21815 14540 21820 14570
rect 21850 14540 21855 14570
rect 21815 14535 21855 14540
rect 21870 14535 21885 14960
rect 22045 14795 22075 14800
rect 21945 14765 22045 14775
rect 23630 14795 23660 14800
rect 21945 14760 22075 14765
rect 22135 14765 22165 14770
rect 21900 14570 21930 14575
rect 21900 14535 21930 14540
rect 21945 14535 21960 14760
rect 22005 14735 22135 14745
rect 23540 14765 23570 14770
rect 22005 14730 22165 14735
rect 22225 14735 22255 14740
rect 22005 14535 22020 14730
rect 22065 14705 22225 14715
rect 23450 14735 23480 14740
rect 22065 14700 22255 14705
rect 22315 14705 22345 14710
rect 22065 14535 22080 14700
rect 22125 14675 22315 14685
rect 23360 14705 23390 14710
rect 22125 14670 22345 14675
rect 22405 14675 22435 14680
rect 22125 14535 22140 14670
rect 22185 14645 22405 14655
rect 23270 14675 23300 14680
rect 22185 14640 22435 14645
rect 22495 14645 22525 14650
rect 22185 14535 22200 14640
rect 22245 14615 22495 14625
rect 23180 14645 23210 14650
rect 22245 14610 22525 14615
rect 22585 14615 22615 14620
rect 22245 14535 22260 14610
rect 22305 14585 22585 14595
rect 23660 14765 23760 14775
rect 23630 14760 23760 14765
rect 23570 14735 23700 14745
rect 23540 14730 23700 14735
rect 23480 14705 23640 14715
rect 23450 14700 23640 14705
rect 23390 14675 23580 14685
rect 23360 14670 23580 14675
rect 23300 14645 23520 14655
rect 23270 14640 23520 14645
rect 23210 14615 23460 14625
rect 23180 14610 23460 14615
rect 22305 14580 22615 14585
rect 22305 14535 22320 14580
rect 23445 14535 23460 14610
rect 23505 14535 23520 14640
rect 23565 14535 23580 14670
rect 23625 14535 23640 14700
rect 23685 14535 23700 14730
rect 23745 14535 23760 14760
rect 24310 14570 24350 14575
rect 23775 14540 23780 14570
rect 23810 14540 23815 14570
rect 23775 14535 23815 14540
rect 24310 14540 24315 14570
rect 24345 14540 24350 14570
rect 24310 14535 24350 14540
rect 24365 14535 24380 14960
rect 24540 14795 24570 14800
rect 24440 14765 24540 14775
rect 26125 14795 26155 14800
rect 24440 14760 24570 14765
rect 24630 14765 24660 14770
rect 24395 14570 24425 14575
rect 24395 14535 24425 14540
rect 24440 14535 24455 14760
rect 24500 14735 24630 14745
rect 26035 14765 26065 14770
rect 24500 14730 24660 14735
rect 24720 14735 24750 14740
rect 24500 14535 24515 14730
rect 24560 14705 24720 14715
rect 25945 14735 25975 14740
rect 24560 14700 24750 14705
rect 24810 14705 24840 14710
rect 24560 14535 24575 14700
rect 24620 14675 24810 14685
rect 25855 14705 25885 14710
rect 24620 14670 24840 14675
rect 24900 14675 24930 14680
rect 24620 14535 24635 14670
rect 24680 14645 24900 14655
rect 26155 14765 26255 14775
rect 26125 14760 26255 14765
rect 26065 14735 26195 14745
rect 26035 14730 26195 14735
rect 25975 14705 26135 14715
rect 25945 14700 26135 14705
rect 25885 14675 26075 14685
rect 25855 14670 26075 14675
rect 24680 14640 24930 14645
rect 24990 14645 25020 14650
rect 24680 14535 24695 14640
rect 24740 14615 24990 14625
rect 24740 14610 25020 14615
rect 24740 14535 24755 14610
rect 26060 14535 26075 14670
rect 26120 14535 26135 14700
rect 26180 14535 26195 14730
rect 26240 14535 26255 14760
rect 26805 14570 26845 14575
rect 26270 14540 26275 14570
rect 26305 14540 26310 14570
rect 26270 14535 26310 14540
rect 26805 14540 26810 14570
rect 26840 14540 26845 14570
rect 26805 14535 26845 14540
rect 26860 14535 26875 14960
rect 27035 14795 27065 14800
rect 26935 14765 27035 14775
rect 28620 14795 28650 14800
rect 26935 14760 27065 14765
rect 27125 14765 27155 14770
rect 26890 14570 26920 14575
rect 26890 14535 26920 14540
rect 26935 14535 26950 14760
rect 26995 14735 27125 14745
rect 28530 14765 28560 14770
rect 26995 14730 27155 14735
rect 27215 14735 27245 14740
rect 26995 14535 27010 14730
rect 27055 14705 27215 14715
rect 28440 14735 28470 14740
rect 27055 14700 27245 14705
rect 27305 14705 27335 14710
rect 27055 14535 27070 14700
rect 27115 14675 27305 14685
rect 27115 14670 27335 14675
rect 28350 14705 28380 14710
rect 28650 14765 28750 14775
rect 28620 14760 28750 14765
rect 28560 14735 28690 14745
rect 28530 14730 28690 14735
rect 28470 14705 28630 14715
rect 28440 14700 28630 14705
rect 28380 14675 28570 14685
rect 28350 14670 28570 14675
rect 27115 14535 27130 14670
rect 28555 14535 28570 14670
rect 28615 14535 28630 14700
rect 28675 14535 28690 14730
rect 28735 14535 28750 14760
rect 29300 14570 29340 14575
rect 28765 14540 28770 14570
rect 28800 14540 28805 14570
rect 28765 14535 28805 14540
rect 29300 14540 29305 14570
rect 29335 14540 29340 14570
rect 29300 14535 29340 14540
rect 29355 14535 29370 14960
rect 29530 14795 29560 14800
rect 29430 14765 29530 14775
rect 31115 14795 31145 14800
rect 29430 14760 29560 14765
rect 29620 14765 29650 14770
rect 29385 14570 29415 14575
rect 29385 14535 29415 14540
rect 29430 14535 29445 14760
rect 29490 14735 29620 14745
rect 31025 14765 31055 14770
rect 29490 14730 29650 14735
rect 29710 14735 29740 14740
rect 29490 14535 29505 14730
rect 29550 14705 29710 14715
rect 31145 14765 31245 14775
rect 31115 14760 31245 14765
rect 31055 14735 31185 14745
rect 31025 14730 31185 14735
rect 29550 14700 29740 14705
rect 29800 14705 29830 14710
rect 29550 14535 29565 14700
rect 29610 14675 29800 14685
rect 29610 14670 29830 14675
rect 29610 14535 29625 14670
rect 31170 14535 31185 14730
rect 31230 14535 31245 14760
rect 31795 14570 31835 14575
rect 31260 14540 31265 14570
rect 31295 14540 31300 14570
rect 31260 14535 31300 14540
rect 31795 14540 31800 14570
rect 31830 14540 31835 14570
rect 31795 14535 31835 14540
rect 31850 14535 31865 14960
rect 32025 14795 32055 14800
rect 31925 14765 32025 14775
rect 33610 14795 33640 14800
rect 31925 14760 32055 14765
rect 32115 14765 32145 14770
rect 31880 14570 31910 14575
rect 31880 14535 31910 14540
rect 31925 14535 31940 14760
rect 31985 14735 32115 14745
rect 31985 14730 32145 14735
rect 33520 14765 33550 14770
rect 33640 14765 33740 14775
rect 33610 14760 33740 14765
rect 33550 14735 33680 14745
rect 33520 14730 33680 14735
rect 31985 14535 32000 14730
rect 33665 14535 33680 14730
rect 33725 14535 33740 14760
rect 34290 14570 34330 14575
rect 33755 14540 33760 14570
rect 33790 14540 33795 14570
rect 33755 14535 33795 14540
rect 34290 14540 34295 14570
rect 34325 14540 34330 14570
rect 34290 14535 34330 14540
rect 34345 14535 34360 14960
rect 34520 14795 34550 14800
rect 34420 14765 34520 14775
rect 36105 14795 36135 14800
rect 34420 14760 34550 14765
rect 34610 14765 34640 14770
rect 34375 14570 34405 14575
rect 34375 14535 34405 14540
rect 34420 14535 34435 14760
rect 34480 14735 34610 14745
rect 36135 14765 36235 14775
rect 36105 14760 36235 14765
rect 34480 14730 34640 14735
rect 34480 14535 34495 14730
rect 36220 14535 36235 14760
rect 36785 14570 36825 14575
rect 36250 14540 36255 14570
rect 36285 14540 36290 14570
rect 36250 14535 36290 14540
rect 36785 14540 36790 14570
rect 36820 14540 36825 14570
rect 36785 14535 36825 14540
rect 36840 14535 36855 14960
rect 37015 14795 37045 14800
rect 36915 14765 37015 14775
rect 36915 14760 37045 14765
rect 38600 14795 38630 14800
rect 38630 14765 38730 14775
rect 38600 14760 38730 14765
rect 36870 14570 36900 14575
rect 36870 14535 36900 14540
rect 36915 14535 36930 14760
rect 38715 14535 38730 14760
rect 39280 14570 39320 14575
rect 38745 14540 38750 14570
rect 38780 14540 38785 14570
rect 38745 14535 38785 14540
rect 39280 14540 39285 14570
rect 39315 14540 39320 14570
rect 39280 14535 39320 14540
rect 39335 14535 39350 14960
rect 39510 14795 39540 14800
rect 39410 14765 39510 14775
rect 39410 14760 39540 14765
rect 39365 14570 39395 14575
rect 39365 14535 39395 14540
rect 39410 14535 39425 14760
rect 41640 14570 41680 14575
rect 41105 14540 41110 14570
rect 41140 14540 41145 14570
rect 41105 14535 41145 14540
rect 41640 14540 41645 14570
rect 41675 14540 41680 14570
rect 41640 14535 41680 14540
rect 41695 14535 41710 14960
rect 41725 14570 41755 14575
rect 41725 14535 41755 14540
rect -2795 14495 -2655 14525
rect -635 14495 -630 14535
rect -590 14495 -585 14535
rect -635 14490 -585 14495
rect 22185 13665 22200 13680
<< via1 >>
rect 2080 16295 2110 16325
rect 4575 16295 4605 16325
rect 7070 16295 7100 16325
rect 9565 16295 9595 16325
rect 12060 16295 12090 16325
rect 14555 16295 14585 16325
rect 17050 16295 17080 16325
rect 19545 16295 19575 16325
rect 22040 16295 22070 16325
rect 24535 16295 24565 16325
rect 27030 16295 27060 16325
rect 29525 16295 29555 16325
rect 32020 16295 32050 16325
rect 34515 16295 34545 16325
rect 37010 16295 37040 16325
rect 39505 16295 39535 16325
rect 2050 16225 2080 16255
rect 4545 16225 4575 16255
rect 7040 16225 7070 16255
rect 9535 16225 9565 16255
rect 12030 16225 12060 16255
rect 14525 16225 14555 16255
rect 17020 16225 17050 16255
rect 19515 16225 19545 16255
rect 22010 16225 22040 16255
rect 24505 16225 24535 16255
rect 27000 16225 27030 16255
rect 29495 16225 29525 16255
rect 31990 16225 32020 16255
rect 34485 16225 34515 16255
rect 36980 16225 37010 16255
rect 39475 16225 39505 16255
rect 7160 16155 7190 16185
rect 9655 16155 9685 16185
rect 12150 16155 12180 16185
rect 14645 16155 14675 16185
rect 17140 16155 17170 16185
rect 19635 16155 19665 16185
rect 22130 16155 22160 16185
rect 24625 16155 24655 16185
rect 27120 16155 27150 16185
rect 29615 16155 29645 16185
rect 32110 16155 32140 16185
rect 34605 16155 34635 16185
rect 7130 16085 7160 16115
rect 9625 16085 9655 16115
rect 12120 16085 12150 16115
rect 14615 16085 14645 16115
rect 17110 16085 17140 16115
rect 19605 16085 19635 16115
rect 22100 16085 22130 16115
rect 24595 16085 24625 16115
rect 27090 16085 27120 16115
rect 29585 16085 29615 16115
rect 32080 16085 32110 16115
rect 34575 16085 34605 16115
rect 12330 16015 12360 16045
rect 14825 16015 14855 16045
rect 17230 16015 17260 16045
rect 19725 16015 19755 16045
rect 22220 16015 22250 16045
rect 24715 16015 24745 16045
rect 27300 16015 27330 16045
rect 29795 16015 29825 16045
rect 12300 15945 12330 15975
rect 14795 15945 14825 15975
rect 17200 15945 17230 15975
rect 19695 15945 19725 15975
rect 22190 15945 22220 15975
rect 24685 15945 24715 15975
rect 27270 15945 27300 15975
rect 29765 15945 29795 15975
rect 12240 15875 12270 15905
rect 14735 15875 14765 15905
rect 17320 15875 17350 15905
rect 19815 15875 19845 15905
rect 22310 15875 22340 15905
rect 24805 15875 24835 15905
rect 27210 15875 27240 15905
rect 29705 15875 29735 15905
rect 12210 15805 12240 15835
rect 14705 15805 14735 15835
rect 17290 15805 17320 15835
rect 19785 15805 19815 15835
rect 22280 15805 22310 15835
rect 24775 15805 24805 15835
rect 27180 15805 27210 15835
rect 29675 15805 29705 15835
rect 17500 15735 17530 15765
rect 19905 15735 19935 15765
rect 22400 15735 22430 15765
rect 24985 15735 25015 15765
rect 17470 15665 17500 15695
rect 19875 15665 19905 15695
rect 22370 15665 22400 15695
rect 24955 15665 24985 15695
rect 17410 15595 17440 15625
rect 24895 15595 24925 15625
rect 17380 15525 17410 15555
rect 24865 15525 24895 15555
rect 19995 15455 20025 15485
rect 22580 15455 22610 15485
rect 19965 15385 19995 15415
rect 22550 15385 22580 15415
rect 22505 15315 22535 15345
rect 22460 15245 22490 15275
rect 20085 15175 20115 15205
rect 20050 15105 20080 15135
rect -2550 15060 -2520 15090
rect -2755 15030 -2725 15060
rect -425 15030 -395 15060
rect 1935 15030 1965 15060
rect 4430 15030 4460 15060
rect 6925 15030 6955 15060
rect 9420 15030 9450 15060
rect 11915 15030 11945 15060
rect 14410 15030 14440 15060
rect 16905 15030 16935 15060
rect 19400 15030 19430 15060
rect 21895 15030 21925 15060
rect 24390 15030 24420 15060
rect 26885 15030 26915 15060
rect 29380 15030 29410 15060
rect 31875 15030 31905 15060
rect 34370 15030 34400 15060
rect 36865 15030 36895 15060
rect 39360 15030 39390 15060
rect 41720 15030 41750 15060
rect -2620 14965 -2590 14995
rect -2680 14895 -2650 14925
rect 1175 14765 1205 14795
rect -1035 14540 -1005 14570
rect -500 14540 -470 14570
rect -420 14540 -390 14570
rect 1325 14540 1355 14570
rect 1860 14540 1890 14570
rect 2085 14765 2115 14795
rect 3670 14765 3700 14795
rect 1940 14540 1970 14570
rect 3820 14540 3850 14570
rect 4355 14540 4385 14570
rect 4580 14765 4610 14795
rect 4435 14540 4465 14570
rect 6075 14735 6105 14765
rect 6165 14765 6195 14795
rect 6315 14540 6345 14570
rect 6850 14540 6880 14570
rect 7075 14765 7105 14795
rect 6930 14540 6960 14570
rect 7165 14735 7195 14765
rect 8570 14735 8600 14765
rect 8660 14765 8690 14795
rect 8810 14540 8840 14570
rect 9345 14540 9375 14570
rect 9570 14765 9600 14795
rect 9425 14540 9455 14570
rect 9660 14735 9690 14765
rect 10885 14675 10915 14705
rect 10975 14705 11005 14735
rect 11065 14735 11095 14765
rect 11155 14765 11185 14795
rect 11305 14540 11335 14570
rect 11840 14540 11870 14570
rect 12065 14765 12095 14795
rect 11920 14540 11950 14570
rect 12155 14735 12185 14765
rect 12245 14705 12275 14735
rect 12335 14675 12365 14705
rect 13380 14675 13410 14705
rect 13470 14705 13500 14735
rect 13560 14735 13590 14765
rect 13650 14765 13680 14795
rect 13800 14540 13830 14570
rect 14335 14540 14365 14570
rect 14560 14765 14590 14795
rect 14415 14540 14445 14570
rect 14650 14735 14680 14765
rect 14740 14705 14770 14735
rect 14830 14675 14860 14705
rect 15695 14615 15725 14645
rect 15785 14645 15815 14675
rect 15875 14675 15905 14705
rect 15965 14705 15995 14735
rect 16055 14735 16085 14765
rect 16145 14765 16175 14795
rect 16295 14540 16325 14570
rect 16830 14540 16860 14570
rect 17055 14765 17085 14795
rect 16910 14540 16940 14570
rect 17145 14735 17175 14765
rect 17235 14705 17265 14735
rect 17325 14675 17355 14705
rect 17415 14645 17445 14675
rect 17505 14615 17535 14645
rect 18100 14585 18130 14615
rect 18190 14615 18220 14645
rect 18280 14645 18310 14675
rect 18370 14675 18400 14705
rect 18460 14705 18490 14735
rect 18550 14735 18580 14765
rect 18640 14765 18670 14795
rect 18790 14540 18820 14570
rect 19325 14540 19355 14570
rect 19550 14765 19580 14795
rect 19405 14540 19435 14570
rect 19640 14735 19670 14765
rect 19730 14705 19760 14735
rect 19820 14675 19850 14705
rect 19910 14645 19940 14675
rect 20000 14615 20030 14645
rect 20090 14585 20120 14615
rect 20595 14585 20625 14615
rect 20685 14615 20715 14645
rect 20775 14645 20805 14675
rect 20865 14675 20895 14705
rect 20955 14705 20985 14735
rect 21045 14735 21075 14765
rect 21135 14765 21165 14795
rect 21285 14540 21315 14570
rect 21820 14540 21850 14570
rect 22045 14765 22075 14795
rect 21900 14540 21930 14570
rect 22135 14735 22165 14765
rect 22225 14705 22255 14735
rect 22315 14675 22345 14705
rect 22405 14645 22435 14675
rect 22495 14615 22525 14645
rect 22585 14585 22615 14615
rect 23180 14615 23210 14645
rect 23270 14645 23300 14675
rect 23360 14675 23390 14705
rect 23450 14705 23480 14735
rect 23540 14735 23570 14765
rect 23630 14765 23660 14795
rect 23780 14540 23810 14570
rect 24315 14540 24345 14570
rect 24540 14765 24570 14795
rect 24395 14540 24425 14570
rect 24630 14735 24660 14765
rect 24720 14705 24750 14735
rect 24810 14675 24840 14705
rect 24900 14645 24930 14675
rect 25855 14675 25885 14705
rect 25945 14705 25975 14735
rect 26035 14735 26065 14765
rect 26125 14765 26155 14795
rect 24990 14615 25020 14645
rect 26275 14540 26305 14570
rect 26810 14540 26840 14570
rect 27035 14765 27065 14795
rect 26890 14540 26920 14570
rect 27125 14735 27155 14765
rect 27215 14705 27245 14735
rect 27305 14675 27335 14705
rect 28350 14675 28380 14705
rect 28440 14705 28470 14735
rect 28530 14735 28560 14765
rect 28620 14765 28650 14795
rect 28770 14540 28800 14570
rect 29305 14540 29335 14570
rect 29530 14765 29560 14795
rect 29385 14540 29415 14570
rect 29620 14735 29650 14765
rect 29710 14705 29740 14735
rect 31025 14735 31055 14765
rect 31115 14765 31145 14795
rect 29800 14675 29830 14705
rect 31265 14540 31295 14570
rect 31800 14540 31830 14570
rect 32025 14765 32055 14795
rect 31880 14540 31910 14570
rect 32115 14735 32145 14765
rect 33520 14735 33550 14765
rect 33610 14765 33640 14795
rect 33760 14540 33790 14570
rect 34295 14540 34325 14570
rect 34520 14765 34550 14795
rect 34375 14540 34405 14570
rect 34610 14735 34640 14765
rect 36105 14765 36135 14795
rect 36255 14540 36285 14570
rect 36790 14540 36820 14570
rect 37015 14765 37045 14795
rect 38600 14765 38630 14795
rect 36870 14540 36900 14570
rect 38750 14540 38780 14570
rect 39285 14540 39315 14570
rect 39510 14765 39540 14795
rect 39365 14540 39395 14570
rect 41110 14540 41140 14570
rect 41645 14540 41675 14570
rect 41725 14540 41755 14570
rect -630 14495 -590 14535
<< metal2 >>
rect 1175 16330 1215 16335
rect 1175 16300 1180 16330
rect 1210 16300 1215 16330
rect 3670 16330 3710 16335
rect 1175 16295 1215 16300
rect 2075 16295 2080 16325
rect 2110 16295 2115 16325
rect -2765 15060 -2715 15070
rect -2765 15030 -2755 15060
rect -2725 15030 -2715 15060
rect -2765 15020 -2715 15030
rect -2555 15060 -2550 15090
rect -2520 15060 -2515 15090
rect -505 15065 -465 15070
rect -2555 15000 -2540 15060
rect -505 15035 -500 15065
rect -470 15035 -465 15065
rect -505 15030 -465 15035
rect -430 15030 -425 15060
rect -395 15030 -390 15060
rect -2625 14995 -2585 15000
rect -2625 14965 -2620 14995
rect -2590 14965 -2585 14995
rect -2625 14960 -2585 14965
rect -2555 14995 -2515 15000
rect -2555 14965 -2550 14995
rect -2520 14965 -2515 14995
rect -2555 14960 -2515 14965
rect -1040 14995 -1000 15000
rect -1040 14965 -1035 14995
rect -1005 14965 -1000 14995
rect -1040 14960 -1000 14965
rect -2685 14925 -2645 14930
rect -2685 14895 -2680 14925
rect -2650 14895 -2645 14925
rect -2685 14890 -2645 14895
rect -1040 14570 -1005 14960
rect -500 14575 -465 15030
rect -405 14575 -390 15030
rect 1175 14800 1190 16295
rect 1205 16260 1245 16265
rect 1205 16230 1210 16260
rect 1240 16230 1245 16260
rect 1205 16225 1245 16230
rect 2045 16225 2050 16255
rect 2080 16225 2085 16255
rect 1175 14795 1205 14800
rect 1175 14760 1205 14765
rect 1220 14775 1235 16225
rect 1855 15065 1895 15070
rect 1855 15035 1860 15065
rect 1890 15035 1895 15065
rect 1855 15030 1895 15035
rect 1930 15030 1935 15060
rect 1965 15030 1970 15060
rect 1320 14995 1360 15000
rect 1320 14965 1325 14995
rect 1355 14965 1360 14995
rect 1320 14960 1360 14965
rect 1220 14760 1305 14775
rect -505 14570 -465 14575
rect -1040 14540 -1035 14570
rect -1005 14540 -1000 14570
rect -505 14540 -500 14570
rect -470 14540 -465 14570
rect -1040 14535 -1000 14540
rect -635 14535 -585 14540
rect -505 14535 -465 14540
rect -420 14570 -390 14575
rect -420 14535 -390 14540
rect 1290 14535 1305 14760
rect 1320 14570 1355 14960
rect 1860 14575 1895 15030
rect 1955 14575 1970 15030
rect 2055 14775 2070 16225
rect 2100 14800 2115 16295
rect 1855 14570 1895 14575
rect 1320 14540 1325 14570
rect 1355 14540 1360 14570
rect 1320 14535 1360 14540
rect 1855 14540 1860 14570
rect 1890 14540 1895 14570
rect 1855 14535 1895 14540
rect 1940 14570 1970 14575
rect 1940 14535 1970 14540
rect 1985 14760 2070 14775
rect 2085 14795 2115 14800
rect 2085 14760 2115 14765
rect 3670 16300 3675 16330
rect 3705 16300 3710 16330
rect 6165 16330 6205 16335
rect 3670 16295 3710 16300
rect 4570 16295 4575 16325
rect 4605 16295 4610 16325
rect 3670 14800 3685 16295
rect 3700 16260 3740 16265
rect 3700 16230 3705 16260
rect 3735 16230 3740 16260
rect 3700 16225 3740 16230
rect 4540 16225 4545 16255
rect 4575 16225 4580 16255
rect 3670 14795 3700 14800
rect 3670 14760 3700 14765
rect 3715 14775 3730 16225
rect 4350 15065 4390 15070
rect 4350 15035 4355 15065
rect 4385 15035 4390 15065
rect 4350 15030 4390 15035
rect 4425 15030 4430 15060
rect 4460 15030 4465 15060
rect 3815 14995 3855 15000
rect 3815 14965 3820 14995
rect 3850 14965 3855 14995
rect 3815 14960 3855 14965
rect 3715 14760 3800 14775
rect 1985 14535 2000 14760
rect 3785 14535 3800 14760
rect 3815 14570 3850 14960
rect 4355 14575 4390 15030
rect 4450 14575 4465 15030
rect 4550 14775 4565 16225
rect 4595 14800 4610 16295
rect 6165 16300 6170 16330
rect 6200 16300 6205 16330
rect 8660 16330 8700 16335
rect 6165 16295 6205 16300
rect 7065 16295 7070 16325
rect 7100 16295 7105 16325
rect 4350 14570 4390 14575
rect 3815 14540 3820 14570
rect 3850 14540 3855 14570
rect 3815 14535 3855 14540
rect 4350 14540 4355 14570
rect 4385 14540 4390 14570
rect 4350 14535 4390 14540
rect 4435 14570 4465 14575
rect 4435 14535 4465 14540
rect 4480 14760 4565 14775
rect 4580 14795 4610 14800
rect 4580 14760 4610 14765
rect 6075 16190 6115 16195
rect 6075 16160 6080 16190
rect 6110 16160 6115 16190
rect 6075 16155 6115 16160
rect 6075 14770 6090 16155
rect 6105 16120 6145 16125
rect 6105 16090 6110 16120
rect 6140 16090 6145 16120
rect 6105 16085 6145 16090
rect 6075 14765 6105 14770
rect 4480 14535 4495 14760
rect 6075 14730 6105 14735
rect 6120 14745 6135 16085
rect 6165 14800 6180 16295
rect 6195 16260 6235 16265
rect 6195 16230 6200 16260
rect 6230 16230 6235 16260
rect 6195 16225 6235 16230
rect 7035 16225 7040 16255
rect 7070 16225 7075 16255
rect 6165 14795 6195 14800
rect 6165 14760 6195 14765
rect 6210 14775 6225 16225
rect 6845 15065 6885 15070
rect 6845 15035 6850 15065
rect 6880 15035 6885 15065
rect 6845 15030 6885 15035
rect 6920 15030 6925 15060
rect 6955 15030 6960 15060
rect 6310 14995 6350 15000
rect 6310 14965 6315 14995
rect 6345 14965 6350 14995
rect 6310 14960 6350 14965
rect 6210 14760 6295 14775
rect 6120 14730 6235 14745
rect 6220 14535 6235 14730
rect 6280 14535 6295 14760
rect 6310 14570 6345 14960
rect 6850 14575 6885 15030
rect 6945 14575 6960 15030
rect 7045 14775 7060 16225
rect 7090 14800 7105 16295
rect 8660 16300 8665 16330
rect 8695 16300 8700 16330
rect 11155 16330 11195 16335
rect 8660 16295 8700 16300
rect 9560 16295 9565 16325
rect 9595 16295 9600 16325
rect 8570 16190 8610 16195
rect 7155 16155 7160 16185
rect 7190 16155 7195 16185
rect 7125 16085 7130 16115
rect 7160 16085 7165 16115
rect 6845 14570 6885 14575
rect 6310 14540 6315 14570
rect 6345 14540 6350 14570
rect 6310 14535 6350 14540
rect 6845 14540 6850 14570
rect 6880 14540 6885 14570
rect 6845 14535 6885 14540
rect 6930 14570 6960 14575
rect 6930 14535 6960 14540
rect 6975 14760 7060 14775
rect 7075 14795 7105 14800
rect 7075 14760 7105 14765
rect 6975 14535 6990 14760
rect 7135 14745 7150 16085
rect 7180 14770 7195 16155
rect 7035 14730 7150 14745
rect 7165 14765 7195 14770
rect 7165 14730 7195 14735
rect 8570 16160 8575 16190
rect 8605 16160 8610 16190
rect 8570 16155 8610 16160
rect 8570 14770 8585 16155
rect 8600 16120 8640 16125
rect 8600 16090 8605 16120
rect 8635 16090 8640 16120
rect 8600 16085 8640 16090
rect 8570 14765 8600 14770
rect 8570 14730 8600 14735
rect 8615 14745 8630 16085
rect 8660 14800 8675 16295
rect 8690 16260 8730 16265
rect 8690 16230 8695 16260
rect 8725 16230 8730 16260
rect 8690 16225 8730 16230
rect 9530 16225 9535 16255
rect 9565 16225 9570 16255
rect 8660 14795 8690 14800
rect 8660 14760 8690 14765
rect 8705 14775 8720 16225
rect 9340 15065 9380 15070
rect 9340 15035 9345 15065
rect 9375 15035 9380 15065
rect 9340 15030 9380 15035
rect 9415 15030 9420 15060
rect 9450 15030 9455 15060
rect 8805 14995 8845 15000
rect 8805 14965 8810 14995
rect 8840 14965 8845 14995
rect 8805 14960 8845 14965
rect 8705 14760 8790 14775
rect 8615 14730 8730 14745
rect 7035 14535 7050 14730
rect 8715 14535 8730 14730
rect 8775 14535 8790 14760
rect 8805 14570 8840 14960
rect 9345 14575 9380 15030
rect 9440 14575 9455 15030
rect 9540 14775 9555 16225
rect 9585 14800 9600 16295
rect 11155 16300 11160 16330
rect 11190 16300 11195 16330
rect 13650 16330 13690 16335
rect 11155 16295 11195 16300
rect 12055 16295 12060 16325
rect 12090 16295 12095 16325
rect 11065 16190 11105 16195
rect 9650 16155 9655 16185
rect 9685 16155 9690 16185
rect 9620 16085 9625 16115
rect 9655 16085 9660 16115
rect 9340 14570 9380 14575
rect 8805 14540 8810 14570
rect 8840 14540 8845 14570
rect 8805 14535 8845 14540
rect 9340 14540 9345 14570
rect 9375 14540 9380 14570
rect 9340 14535 9380 14540
rect 9425 14570 9455 14575
rect 9425 14535 9455 14540
rect 9470 14760 9555 14775
rect 9570 14795 9600 14800
rect 9570 14760 9600 14765
rect 9470 14535 9485 14760
rect 9630 14745 9645 16085
rect 9675 14770 9690 16155
rect 11065 16160 11070 16190
rect 11100 16160 11105 16190
rect 11065 16155 11105 16160
rect 9530 14730 9645 14745
rect 9660 14765 9690 14770
rect 9660 14730 9690 14735
rect 10885 16050 10925 16055
rect 10885 16020 10890 16050
rect 10920 16020 10925 16050
rect 10885 16015 10925 16020
rect 9530 14535 9545 14730
rect 10885 14710 10900 16015
rect 10915 15980 10955 15985
rect 10915 15950 10920 15980
rect 10950 15950 10955 15980
rect 10915 15945 10955 15950
rect 10885 14705 10915 14710
rect 10885 14670 10915 14675
rect 10930 14685 10945 15945
rect 10975 15910 11015 15915
rect 10975 15880 10980 15910
rect 11010 15880 11015 15910
rect 10975 15875 11015 15880
rect 10975 14740 10990 15875
rect 11005 15840 11045 15845
rect 11005 15810 11010 15840
rect 11040 15810 11045 15840
rect 11005 15805 11045 15810
rect 10975 14735 11005 14740
rect 10975 14700 11005 14705
rect 11020 14715 11035 15805
rect 11065 14770 11080 16155
rect 11095 16120 11135 16125
rect 11095 16090 11100 16120
rect 11130 16090 11135 16120
rect 11095 16085 11135 16090
rect 11065 14765 11095 14770
rect 11065 14730 11095 14735
rect 11110 14745 11125 16085
rect 11155 14800 11170 16295
rect 11185 16260 11225 16265
rect 11185 16230 11190 16260
rect 11220 16230 11225 16260
rect 11185 16225 11225 16230
rect 12025 16225 12030 16255
rect 12060 16225 12065 16255
rect 11155 14795 11185 14800
rect 11155 14760 11185 14765
rect 11200 14775 11215 16225
rect 11835 15065 11875 15070
rect 11835 15035 11840 15065
rect 11870 15035 11875 15065
rect 11835 15030 11875 15035
rect 11910 15030 11915 15060
rect 11945 15030 11950 15060
rect 11300 14995 11340 15000
rect 11300 14965 11305 14995
rect 11335 14965 11340 14995
rect 11300 14960 11340 14965
rect 11200 14760 11285 14775
rect 11110 14730 11225 14745
rect 11020 14700 11165 14715
rect 10930 14670 11105 14685
rect 11090 14535 11105 14670
rect 11150 14535 11165 14700
rect 11210 14535 11225 14730
rect 11270 14535 11285 14760
rect 11300 14570 11335 14960
rect 11840 14575 11875 15030
rect 11935 14575 11950 15030
rect 12035 14775 12050 16225
rect 12080 14800 12095 16295
rect 13650 16300 13655 16330
rect 13685 16300 13690 16330
rect 16145 16330 16185 16335
rect 13650 16295 13690 16300
rect 14550 16295 14555 16325
rect 14585 16295 14590 16325
rect 13560 16190 13600 16195
rect 12145 16155 12150 16185
rect 12180 16155 12185 16185
rect 12115 16085 12120 16115
rect 12150 16085 12155 16115
rect 11835 14570 11875 14575
rect 11300 14540 11305 14570
rect 11335 14540 11340 14570
rect 11300 14535 11340 14540
rect 11835 14540 11840 14570
rect 11870 14540 11875 14570
rect 11835 14535 11875 14540
rect 11920 14570 11950 14575
rect 11920 14535 11950 14540
rect 11965 14760 12050 14775
rect 12065 14795 12095 14800
rect 12065 14760 12095 14765
rect 11965 14535 11980 14760
rect 12125 14745 12140 16085
rect 12170 14770 12185 16155
rect 13560 16160 13565 16190
rect 13595 16160 13600 16190
rect 13560 16155 13600 16160
rect 13380 16050 13420 16055
rect 12325 16015 12330 16045
rect 12360 16015 12365 16045
rect 12295 15945 12300 15975
rect 12330 15945 12335 15975
rect 12235 15875 12240 15905
rect 12270 15875 12275 15905
rect 12205 15805 12210 15835
rect 12240 15805 12245 15835
rect 12025 14730 12140 14745
rect 12155 14765 12185 14770
rect 12155 14730 12185 14735
rect 12025 14535 12040 14730
rect 12215 14715 12230 15805
rect 12260 14740 12275 15875
rect 12085 14700 12230 14715
rect 12245 14735 12275 14740
rect 12245 14700 12275 14705
rect 12085 14535 12100 14700
rect 12305 14685 12320 15945
rect 12350 14710 12365 16015
rect 12145 14670 12320 14685
rect 12335 14705 12365 14710
rect 12335 14670 12365 14675
rect 13380 16020 13385 16050
rect 13415 16020 13420 16050
rect 13380 16015 13420 16020
rect 13380 14710 13395 16015
rect 13410 15980 13450 15985
rect 13410 15950 13415 15980
rect 13445 15950 13450 15980
rect 13410 15945 13450 15950
rect 13380 14705 13410 14710
rect 13380 14670 13410 14675
rect 13425 14685 13440 15945
rect 13470 15910 13510 15915
rect 13470 15880 13475 15910
rect 13505 15880 13510 15910
rect 13470 15875 13510 15880
rect 13470 14740 13485 15875
rect 13500 15840 13540 15845
rect 13500 15810 13505 15840
rect 13535 15810 13540 15840
rect 13500 15805 13540 15810
rect 13470 14735 13500 14740
rect 13470 14700 13500 14705
rect 13515 14715 13530 15805
rect 13560 14770 13575 16155
rect 13590 16120 13630 16125
rect 13590 16090 13595 16120
rect 13625 16090 13630 16120
rect 13590 16085 13630 16090
rect 13560 14765 13590 14770
rect 13560 14730 13590 14735
rect 13605 14745 13620 16085
rect 13650 14800 13665 16295
rect 13680 16260 13720 16265
rect 13680 16230 13685 16260
rect 13715 16230 13720 16260
rect 13680 16225 13720 16230
rect 14520 16225 14525 16255
rect 14555 16225 14560 16255
rect 13650 14795 13680 14800
rect 13650 14760 13680 14765
rect 13695 14775 13710 16225
rect 14330 15065 14370 15070
rect 14330 15035 14335 15065
rect 14365 15035 14370 15065
rect 14330 15030 14370 15035
rect 14405 15030 14410 15060
rect 14440 15030 14445 15060
rect 13795 14995 13835 15000
rect 13795 14965 13800 14995
rect 13830 14965 13835 14995
rect 13795 14960 13835 14965
rect 13695 14760 13780 14775
rect 13605 14730 13720 14745
rect 13515 14700 13660 14715
rect 13425 14670 13600 14685
rect 12145 14535 12160 14670
rect 13585 14535 13600 14670
rect 13645 14535 13660 14700
rect 13705 14535 13720 14730
rect 13765 14535 13780 14760
rect 13795 14570 13830 14960
rect 14335 14575 14370 15030
rect 14430 14575 14445 15030
rect 14530 14775 14545 16225
rect 14575 14800 14590 16295
rect 16145 16300 16150 16330
rect 16180 16300 16185 16330
rect 18640 16330 18680 16335
rect 16145 16295 16185 16300
rect 17045 16295 17050 16325
rect 17080 16295 17085 16325
rect 16055 16190 16095 16195
rect 14640 16155 14645 16185
rect 14675 16155 14680 16185
rect 14610 16085 14615 16115
rect 14645 16085 14650 16115
rect 14330 14570 14370 14575
rect 13795 14540 13800 14570
rect 13830 14540 13835 14570
rect 13795 14535 13835 14540
rect 14330 14540 14335 14570
rect 14365 14540 14370 14570
rect 14330 14535 14370 14540
rect 14415 14570 14445 14575
rect 14415 14535 14445 14540
rect 14460 14760 14545 14775
rect 14560 14795 14590 14800
rect 14560 14760 14590 14765
rect 14460 14535 14475 14760
rect 14620 14745 14635 16085
rect 14665 14770 14680 16155
rect 16055 16160 16060 16190
rect 16090 16160 16095 16190
rect 16055 16155 16095 16160
rect 15965 16050 16005 16055
rect 14820 16015 14825 16045
rect 14855 16015 14860 16045
rect 14790 15945 14795 15975
rect 14825 15945 14830 15975
rect 14730 15875 14735 15905
rect 14765 15875 14770 15905
rect 14700 15805 14705 15835
rect 14735 15805 14740 15835
rect 14520 14730 14635 14745
rect 14650 14765 14680 14770
rect 14650 14730 14680 14735
rect 14520 14535 14535 14730
rect 14710 14715 14725 15805
rect 14755 14740 14770 15875
rect 14580 14700 14725 14715
rect 14740 14735 14770 14740
rect 14740 14700 14770 14705
rect 14580 14535 14595 14700
rect 14800 14685 14815 15945
rect 14845 14710 14860 16015
rect 15965 16020 15970 16050
rect 16000 16020 16005 16050
rect 15965 16015 16005 16020
rect 15875 15910 15915 15915
rect 15875 15880 15880 15910
rect 15910 15880 15915 15910
rect 15875 15875 15915 15880
rect 14640 14670 14815 14685
rect 14830 14705 14860 14710
rect 14830 14670 14860 14675
rect 15695 15770 15735 15775
rect 15695 15740 15700 15770
rect 15730 15740 15735 15770
rect 15695 15735 15735 15740
rect 14640 14535 14655 14670
rect 15695 14650 15710 15735
rect 15725 15700 15765 15705
rect 15725 15670 15730 15700
rect 15760 15670 15765 15700
rect 15725 15665 15765 15670
rect 15695 14645 15725 14650
rect 15695 14610 15725 14615
rect 15740 14625 15755 15665
rect 15785 15630 15825 15635
rect 15785 15600 15790 15630
rect 15820 15600 15825 15630
rect 15785 15595 15825 15600
rect 15785 14680 15800 15595
rect 15815 15560 15855 15565
rect 15815 15530 15820 15560
rect 15850 15530 15855 15560
rect 15815 15525 15855 15530
rect 15785 14675 15815 14680
rect 15785 14640 15815 14645
rect 15830 14655 15845 15525
rect 15875 14710 15890 15875
rect 15905 15840 15945 15845
rect 15905 15810 15910 15840
rect 15940 15810 15945 15840
rect 15905 15805 15945 15810
rect 15875 14705 15905 14710
rect 15875 14670 15905 14675
rect 15920 14685 15935 15805
rect 15965 14740 15980 16015
rect 15995 15980 16035 15985
rect 15995 15950 16000 15980
rect 16030 15950 16035 15980
rect 15995 15945 16035 15950
rect 15965 14735 15995 14740
rect 15965 14700 15995 14705
rect 16010 14715 16025 15945
rect 16055 14770 16070 16155
rect 16085 16120 16125 16125
rect 16085 16090 16090 16120
rect 16120 16090 16125 16120
rect 16085 16085 16125 16090
rect 16055 14765 16085 14770
rect 16055 14730 16085 14735
rect 16100 14745 16115 16085
rect 16145 14800 16160 16295
rect 16175 16260 16215 16265
rect 16175 16230 16180 16260
rect 16210 16230 16215 16260
rect 16175 16225 16215 16230
rect 17015 16225 17020 16255
rect 17050 16225 17055 16255
rect 16145 14795 16175 14800
rect 16145 14760 16175 14765
rect 16190 14775 16205 16225
rect 16825 15065 16865 15070
rect 16825 15035 16830 15065
rect 16860 15035 16865 15065
rect 16825 15030 16865 15035
rect 16900 15030 16905 15060
rect 16935 15030 16940 15060
rect 16290 14995 16330 15000
rect 16290 14965 16295 14995
rect 16325 14965 16330 14995
rect 16290 14960 16330 14965
rect 16190 14760 16275 14775
rect 16100 14730 16215 14745
rect 16010 14700 16155 14715
rect 15920 14670 16095 14685
rect 15830 14640 16035 14655
rect 15740 14610 15975 14625
rect 15960 14535 15975 14610
rect 16020 14535 16035 14640
rect 16080 14535 16095 14670
rect 16140 14535 16155 14700
rect 16200 14535 16215 14730
rect 16260 14535 16275 14760
rect 16290 14570 16325 14960
rect 16830 14575 16865 15030
rect 16925 14575 16940 15030
rect 17025 14775 17040 16225
rect 17070 14800 17085 16295
rect 18640 16300 18645 16330
rect 18675 16300 18680 16330
rect 21135 16330 21175 16335
rect 18640 16295 18680 16300
rect 19540 16295 19545 16325
rect 19575 16295 19580 16325
rect 18550 16190 18590 16195
rect 17135 16155 17140 16185
rect 17170 16155 17175 16185
rect 17105 16085 17110 16115
rect 17140 16085 17145 16115
rect 16825 14570 16865 14575
rect 16290 14540 16295 14570
rect 16325 14540 16330 14570
rect 16290 14535 16330 14540
rect 16825 14540 16830 14570
rect 16860 14540 16865 14570
rect 16825 14535 16865 14540
rect 16910 14570 16940 14575
rect 16910 14535 16940 14540
rect 16955 14760 17040 14775
rect 17055 14795 17085 14800
rect 17055 14760 17085 14765
rect 16955 14535 16970 14760
rect 17115 14745 17130 16085
rect 17160 14770 17175 16155
rect 18550 16160 18555 16190
rect 18585 16160 18590 16190
rect 18550 16155 18590 16160
rect 18460 16050 18500 16055
rect 17225 16015 17230 16045
rect 17260 16015 17265 16045
rect 17195 15945 17200 15975
rect 17230 15945 17235 15975
rect 17015 14730 17130 14745
rect 17145 14765 17175 14770
rect 17145 14730 17175 14735
rect 17015 14535 17030 14730
rect 17205 14715 17220 15945
rect 17250 14740 17265 16015
rect 18460 16020 18465 16050
rect 18495 16020 18500 16050
rect 18460 16015 18500 16020
rect 18370 15910 18410 15915
rect 17315 15875 17320 15905
rect 17350 15875 17355 15905
rect 17285 15805 17290 15835
rect 17320 15805 17325 15835
rect 17075 14700 17220 14715
rect 17235 14735 17265 14740
rect 17235 14700 17265 14705
rect 17075 14535 17090 14700
rect 17295 14685 17310 15805
rect 17340 14710 17355 15875
rect 18370 15880 18375 15910
rect 18405 15880 18410 15910
rect 18370 15875 18410 15880
rect 18280 15770 18320 15775
rect 17495 15735 17500 15765
rect 17530 15735 17535 15765
rect 17465 15665 17470 15695
rect 17500 15665 17505 15695
rect 17405 15595 17410 15625
rect 17440 15595 17445 15625
rect 17375 15525 17380 15555
rect 17410 15525 17415 15555
rect 17135 14670 17310 14685
rect 17325 14705 17355 14710
rect 17325 14670 17355 14675
rect 17135 14535 17150 14670
rect 17385 14655 17400 15525
rect 17430 14680 17445 15595
rect 17195 14640 17400 14655
rect 17415 14675 17445 14680
rect 17415 14640 17445 14645
rect 17195 14535 17210 14640
rect 17475 14625 17490 15665
rect 17520 14650 17535 15735
rect 18280 15740 18285 15770
rect 18315 15740 18320 15770
rect 18280 15735 18320 15740
rect 18190 15490 18230 15495
rect 18190 15460 18195 15490
rect 18225 15460 18230 15490
rect 18190 15455 18230 15460
rect 17255 14610 17490 14625
rect 17505 14645 17535 14650
rect 17505 14610 17535 14615
rect 18100 15210 18140 15215
rect 18100 15180 18105 15210
rect 18135 15180 18140 15210
rect 18100 15175 18140 15180
rect 18100 14620 18115 15175
rect 18130 15140 18170 15145
rect 18130 15110 18135 15140
rect 18165 15110 18170 15140
rect 18130 15105 18170 15110
rect 18100 14615 18130 14620
rect 17255 14535 17270 14610
rect 18100 14580 18130 14585
rect 18145 14595 18160 15105
rect 18190 14650 18205 15455
rect 18220 15420 18260 15425
rect 18220 15390 18225 15420
rect 18255 15390 18260 15420
rect 18220 15385 18260 15390
rect 18190 14645 18220 14650
rect 18190 14610 18220 14615
rect 18235 14625 18250 15385
rect 18280 14680 18295 15735
rect 18310 15700 18350 15705
rect 18310 15670 18315 15700
rect 18345 15670 18350 15700
rect 18310 15665 18350 15670
rect 18280 14675 18310 14680
rect 18280 14640 18310 14645
rect 18325 14655 18340 15665
rect 18370 14710 18385 15875
rect 18400 15840 18440 15845
rect 18400 15810 18405 15840
rect 18435 15810 18440 15840
rect 18400 15805 18440 15810
rect 18370 14705 18400 14710
rect 18370 14670 18400 14675
rect 18415 14685 18430 15805
rect 18460 14740 18475 16015
rect 18490 15980 18530 15985
rect 18490 15950 18495 15980
rect 18525 15950 18530 15980
rect 18490 15945 18530 15950
rect 18460 14735 18490 14740
rect 18460 14700 18490 14705
rect 18505 14715 18520 15945
rect 18550 14770 18565 16155
rect 18580 16120 18620 16125
rect 18580 16090 18585 16120
rect 18615 16090 18620 16120
rect 18580 16085 18620 16090
rect 18550 14765 18580 14770
rect 18550 14730 18580 14735
rect 18595 14745 18610 16085
rect 18640 14800 18655 16295
rect 18670 16260 18710 16265
rect 18670 16230 18675 16260
rect 18705 16230 18710 16260
rect 18670 16225 18710 16230
rect 19510 16225 19515 16255
rect 19545 16225 19550 16255
rect 18640 14795 18670 14800
rect 18640 14760 18670 14765
rect 18685 14775 18700 16225
rect 19320 15065 19360 15070
rect 19320 15035 19325 15065
rect 19355 15035 19360 15065
rect 19320 15030 19360 15035
rect 19395 15030 19400 15060
rect 19430 15030 19435 15060
rect 18785 14995 18825 15000
rect 18785 14965 18790 14995
rect 18820 14965 18825 14995
rect 18785 14960 18825 14965
rect 18685 14760 18770 14775
rect 18595 14730 18710 14745
rect 18505 14700 18650 14715
rect 18415 14670 18590 14685
rect 18325 14640 18530 14655
rect 18235 14610 18470 14625
rect 18145 14580 18410 14595
rect 18395 14535 18410 14580
rect 18455 14535 18470 14610
rect 18515 14535 18530 14640
rect 18575 14535 18590 14670
rect 18635 14535 18650 14700
rect 18695 14535 18710 14730
rect 18755 14535 18770 14760
rect 18785 14570 18820 14960
rect 19325 14575 19360 15030
rect 19420 14575 19435 15030
rect 19520 14775 19535 16225
rect 19565 14800 19580 16295
rect 21135 16300 21140 16330
rect 21170 16300 21175 16330
rect 23630 16330 23670 16335
rect 21135 16295 21175 16300
rect 22035 16295 22040 16325
rect 22070 16295 22075 16325
rect 21045 16190 21085 16195
rect 19630 16155 19635 16185
rect 19665 16155 19670 16185
rect 19600 16085 19605 16115
rect 19635 16085 19640 16115
rect 19320 14570 19360 14575
rect 18785 14540 18790 14570
rect 18820 14540 18825 14570
rect 18785 14535 18825 14540
rect 19320 14540 19325 14570
rect 19355 14540 19360 14570
rect 19320 14535 19360 14540
rect 19405 14570 19435 14575
rect 19405 14535 19435 14540
rect 19450 14760 19535 14775
rect 19550 14795 19580 14800
rect 19550 14760 19580 14765
rect 19450 14535 19465 14760
rect 19610 14745 19625 16085
rect 19655 14770 19670 16155
rect 21045 16160 21050 16190
rect 21080 16160 21085 16190
rect 21045 16155 21085 16160
rect 20955 16050 20995 16055
rect 19720 16015 19725 16045
rect 19755 16015 19760 16045
rect 19690 15945 19695 15975
rect 19725 15945 19730 15975
rect 19510 14730 19625 14745
rect 19640 14765 19670 14770
rect 19640 14730 19670 14735
rect 19510 14535 19525 14730
rect 19700 14715 19715 15945
rect 19745 14740 19760 16015
rect 20955 16020 20960 16050
rect 20990 16020 20995 16050
rect 20955 16015 20995 16020
rect 20865 15910 20905 15915
rect 19810 15875 19815 15905
rect 19845 15875 19850 15905
rect 19780 15805 19785 15835
rect 19815 15805 19820 15835
rect 19570 14700 19715 14715
rect 19730 14735 19760 14740
rect 19730 14700 19760 14705
rect 19570 14535 19585 14700
rect 19790 14685 19805 15805
rect 19835 14710 19850 15875
rect 20865 15880 20870 15910
rect 20900 15880 20905 15910
rect 20865 15875 20905 15880
rect 20775 15770 20815 15775
rect 19900 15735 19905 15765
rect 19935 15735 19940 15765
rect 19870 15665 19875 15695
rect 19905 15665 19910 15695
rect 19630 14670 19805 14685
rect 19820 14705 19850 14710
rect 19820 14670 19850 14675
rect 19630 14535 19645 14670
rect 19880 14655 19895 15665
rect 19925 14680 19940 15735
rect 20775 15740 20780 15770
rect 20810 15740 20815 15770
rect 20775 15735 20815 15740
rect 20595 15490 20635 15495
rect 19990 15455 19995 15485
rect 20025 15455 20030 15485
rect 19960 15385 19965 15415
rect 19995 15385 20000 15415
rect 19690 14640 19895 14655
rect 19910 14675 19940 14680
rect 19910 14640 19940 14645
rect 19690 14535 19705 14640
rect 19970 14625 19985 15385
rect 20015 14650 20030 15455
rect 20595 15460 20600 15490
rect 20630 15460 20635 15490
rect 20595 15455 20635 15460
rect 20080 15175 20085 15205
rect 20115 15175 20120 15205
rect 20045 15105 20050 15135
rect 20080 15105 20085 15135
rect 19750 14610 19985 14625
rect 20000 14645 20030 14650
rect 20000 14610 20030 14615
rect 19750 14535 19765 14610
rect 20060 14595 20075 15105
rect 20105 14620 20120 15175
rect 19810 14580 20075 14595
rect 20090 14615 20120 14620
rect 20090 14580 20120 14585
rect 20595 14620 20610 15455
rect 20625 15420 20665 15425
rect 20625 15390 20630 15420
rect 20660 15390 20665 15420
rect 20625 15385 20665 15390
rect 20595 14615 20625 14620
rect 20595 14580 20625 14585
rect 20640 14595 20655 15385
rect 20670 15350 20710 15355
rect 20670 15320 20675 15350
rect 20705 15320 20710 15350
rect 20670 15315 20710 15320
rect 20685 14650 20700 15315
rect 20715 15280 20755 15285
rect 20715 15250 20720 15280
rect 20750 15250 20755 15280
rect 20715 15245 20755 15250
rect 20685 14645 20715 14650
rect 20685 14610 20715 14615
rect 20730 14625 20745 15245
rect 20775 14680 20790 15735
rect 20805 15700 20845 15705
rect 20805 15670 20810 15700
rect 20840 15670 20845 15700
rect 20805 15665 20845 15670
rect 20775 14675 20805 14680
rect 20775 14640 20805 14645
rect 20820 14655 20835 15665
rect 20865 14710 20880 15875
rect 20895 15840 20935 15845
rect 20895 15810 20900 15840
rect 20930 15810 20935 15840
rect 20895 15805 20935 15810
rect 20865 14705 20895 14710
rect 20865 14670 20895 14675
rect 20910 14685 20925 15805
rect 20955 14740 20970 16015
rect 20985 15980 21025 15985
rect 20985 15950 20990 15980
rect 21020 15950 21025 15980
rect 20985 15945 21025 15950
rect 20955 14735 20985 14740
rect 20955 14700 20985 14705
rect 21000 14715 21015 15945
rect 21045 14770 21060 16155
rect 21075 16120 21115 16125
rect 21075 16090 21080 16120
rect 21110 16090 21115 16120
rect 21075 16085 21115 16090
rect 21045 14765 21075 14770
rect 21045 14730 21075 14735
rect 21090 14745 21105 16085
rect 21135 14800 21150 16295
rect 21165 16260 21205 16265
rect 21165 16230 21170 16260
rect 21200 16230 21205 16260
rect 21165 16225 21205 16230
rect 22005 16225 22010 16255
rect 22040 16225 22045 16255
rect 21135 14795 21165 14800
rect 21135 14760 21165 14765
rect 21180 14775 21195 16225
rect 21815 15065 21855 15070
rect 21815 15035 21820 15065
rect 21850 15035 21855 15065
rect 21815 15030 21855 15035
rect 21890 15030 21895 15060
rect 21925 15030 21930 15060
rect 21280 14995 21320 15000
rect 21280 14965 21285 14995
rect 21315 14965 21320 14995
rect 21280 14960 21320 14965
rect 21180 14760 21265 14775
rect 21090 14730 21205 14745
rect 21000 14700 21145 14715
rect 20910 14670 21085 14685
rect 20820 14640 21025 14655
rect 20730 14610 20965 14625
rect 20640 14580 20905 14595
rect 19810 14535 19825 14580
rect 20890 14535 20905 14580
rect 20950 14535 20965 14610
rect 21010 14535 21025 14640
rect 21070 14535 21085 14670
rect 21130 14535 21145 14700
rect 21190 14535 21205 14730
rect 21250 14535 21265 14760
rect 21280 14570 21315 14960
rect 21820 14575 21855 15030
rect 21915 14575 21930 15030
rect 22015 14775 22030 16225
rect 22060 14800 22075 16295
rect 23630 16300 23635 16330
rect 23665 16300 23670 16330
rect 26125 16330 26165 16335
rect 23630 16295 23670 16300
rect 24530 16295 24535 16325
rect 24565 16295 24570 16325
rect 23540 16190 23580 16195
rect 22125 16155 22130 16185
rect 22160 16155 22165 16185
rect 22095 16085 22100 16115
rect 22130 16085 22135 16115
rect 21815 14570 21855 14575
rect 21280 14540 21285 14570
rect 21315 14540 21320 14570
rect 21280 14535 21320 14540
rect 21815 14540 21820 14570
rect 21850 14540 21855 14570
rect 21815 14535 21855 14540
rect 21900 14570 21930 14575
rect 21900 14535 21930 14540
rect 21945 14760 22030 14775
rect 22045 14795 22075 14800
rect 22045 14760 22075 14765
rect 21945 14535 21960 14760
rect 22105 14745 22120 16085
rect 22150 14770 22165 16155
rect 23540 16160 23545 16190
rect 23575 16160 23580 16190
rect 23540 16155 23580 16160
rect 23450 16050 23490 16055
rect 22215 16015 22220 16045
rect 22250 16015 22255 16045
rect 22185 15945 22190 15975
rect 22220 15945 22225 15975
rect 22005 14730 22120 14745
rect 22135 14765 22165 14770
rect 22135 14730 22165 14735
rect 22005 14535 22020 14730
rect 22195 14715 22210 15945
rect 22240 14740 22255 16015
rect 23450 16020 23455 16050
rect 23485 16020 23490 16050
rect 23450 16015 23490 16020
rect 23360 15910 23400 15915
rect 22305 15875 22310 15905
rect 22340 15875 22345 15905
rect 22275 15805 22280 15835
rect 22310 15805 22315 15835
rect 22065 14700 22210 14715
rect 22225 14735 22255 14740
rect 22225 14700 22255 14705
rect 22065 14535 22080 14700
rect 22285 14685 22300 15805
rect 22330 14710 22345 15875
rect 23360 15880 23365 15910
rect 23395 15880 23400 15910
rect 23360 15875 23400 15880
rect 23180 15770 23220 15775
rect 22395 15735 22400 15765
rect 22430 15735 22435 15765
rect 22365 15665 22370 15695
rect 22400 15665 22405 15695
rect 22125 14670 22300 14685
rect 22315 14705 22345 14710
rect 22315 14670 22345 14675
rect 22125 14535 22140 14670
rect 22375 14655 22390 15665
rect 22420 14680 22435 15735
rect 23180 15740 23185 15770
rect 23215 15740 23220 15770
rect 23180 15735 23220 15740
rect 22575 15455 22580 15485
rect 22610 15455 22615 15485
rect 22545 15385 22550 15415
rect 22580 15385 22585 15415
rect 22500 15315 22505 15345
rect 22535 15315 22540 15345
rect 22455 15245 22460 15275
rect 22490 15245 22495 15275
rect 22185 14640 22390 14655
rect 22405 14675 22435 14680
rect 22405 14640 22435 14645
rect 22185 14535 22200 14640
rect 22465 14625 22480 15245
rect 22510 14650 22525 15315
rect 22245 14610 22480 14625
rect 22495 14645 22525 14650
rect 22495 14610 22525 14615
rect 22245 14535 22260 14610
rect 22555 14595 22570 15385
rect 22600 14620 22615 15455
rect 22305 14580 22570 14595
rect 22585 14615 22615 14620
rect 23180 14650 23195 15735
rect 23210 15700 23250 15705
rect 23210 15670 23215 15700
rect 23245 15670 23250 15700
rect 23210 15665 23250 15670
rect 23180 14645 23210 14650
rect 23180 14610 23210 14615
rect 23225 14625 23240 15665
rect 23270 15630 23310 15635
rect 23270 15600 23275 15630
rect 23305 15600 23310 15630
rect 23270 15595 23310 15600
rect 23270 14680 23285 15595
rect 23300 15560 23340 15565
rect 23300 15530 23305 15560
rect 23335 15530 23340 15560
rect 23300 15525 23340 15530
rect 23270 14675 23300 14680
rect 23270 14640 23300 14645
rect 23315 14655 23330 15525
rect 23360 14710 23375 15875
rect 23390 15840 23430 15845
rect 23390 15810 23395 15840
rect 23425 15810 23430 15840
rect 23390 15805 23430 15810
rect 23360 14705 23390 14710
rect 23360 14670 23390 14675
rect 23405 14685 23420 15805
rect 23450 14740 23465 16015
rect 23480 15980 23520 15985
rect 23480 15950 23485 15980
rect 23515 15950 23520 15980
rect 23480 15945 23520 15950
rect 23450 14735 23480 14740
rect 23450 14700 23480 14705
rect 23495 14715 23510 15945
rect 23540 14770 23555 16155
rect 23570 16120 23610 16125
rect 23570 16090 23575 16120
rect 23605 16090 23610 16120
rect 23570 16085 23610 16090
rect 23540 14765 23570 14770
rect 23540 14730 23570 14735
rect 23585 14745 23600 16085
rect 23630 14800 23645 16295
rect 23660 16260 23700 16265
rect 23660 16230 23665 16260
rect 23695 16230 23700 16260
rect 23660 16225 23700 16230
rect 24500 16225 24505 16255
rect 24535 16225 24540 16255
rect 23630 14795 23660 14800
rect 23630 14760 23660 14765
rect 23675 14775 23690 16225
rect 24310 15065 24350 15070
rect 24310 15035 24315 15065
rect 24345 15035 24350 15065
rect 24310 15030 24350 15035
rect 24385 15030 24390 15060
rect 24420 15030 24425 15060
rect 23775 14995 23815 15000
rect 23775 14965 23780 14995
rect 23810 14965 23815 14995
rect 23775 14960 23815 14965
rect 23675 14760 23760 14775
rect 23585 14730 23700 14745
rect 23495 14700 23640 14715
rect 23405 14670 23580 14685
rect 23315 14640 23520 14655
rect 23225 14610 23460 14625
rect 22585 14580 22615 14585
rect 22305 14535 22320 14580
rect 23445 14535 23460 14610
rect 23505 14535 23520 14640
rect 23565 14535 23580 14670
rect 23625 14535 23640 14700
rect 23685 14535 23700 14730
rect 23745 14535 23760 14760
rect 23775 14570 23810 14960
rect 24315 14575 24350 15030
rect 24410 14575 24425 15030
rect 24510 14775 24525 16225
rect 24555 14800 24570 16295
rect 26125 16300 26130 16330
rect 26160 16300 26165 16330
rect 28620 16330 28660 16335
rect 26125 16295 26165 16300
rect 27025 16295 27030 16325
rect 27060 16295 27065 16325
rect 26035 16190 26075 16195
rect 24620 16155 24625 16185
rect 24655 16155 24660 16185
rect 24590 16085 24595 16115
rect 24625 16085 24630 16115
rect 24310 14570 24350 14575
rect 23775 14540 23780 14570
rect 23810 14540 23815 14570
rect 23775 14535 23815 14540
rect 24310 14540 24315 14570
rect 24345 14540 24350 14570
rect 24310 14535 24350 14540
rect 24395 14570 24425 14575
rect 24395 14535 24425 14540
rect 24440 14760 24525 14775
rect 24540 14795 24570 14800
rect 24540 14760 24570 14765
rect 24440 14535 24455 14760
rect 24600 14745 24615 16085
rect 24645 14770 24660 16155
rect 26035 16160 26040 16190
rect 26070 16160 26075 16190
rect 26035 16155 26075 16160
rect 25855 16050 25895 16055
rect 24710 16015 24715 16045
rect 24745 16015 24750 16045
rect 24680 15945 24685 15975
rect 24715 15945 24720 15975
rect 24500 14730 24615 14745
rect 24630 14765 24660 14770
rect 24630 14730 24660 14735
rect 24500 14535 24515 14730
rect 24690 14715 24705 15945
rect 24735 14740 24750 16015
rect 25855 16020 25860 16050
rect 25890 16020 25895 16050
rect 25855 16015 25895 16020
rect 24800 15875 24805 15905
rect 24835 15875 24840 15905
rect 24770 15805 24775 15835
rect 24805 15805 24810 15835
rect 24560 14700 24705 14715
rect 24720 14735 24750 14740
rect 24720 14700 24750 14705
rect 24560 14535 24575 14700
rect 24780 14685 24795 15805
rect 24825 14710 24840 15875
rect 24980 15735 24985 15765
rect 25015 15735 25020 15765
rect 24950 15665 24955 15695
rect 24985 15665 24990 15695
rect 24890 15595 24895 15625
rect 24925 15595 24930 15625
rect 24860 15525 24865 15555
rect 24895 15525 24900 15555
rect 24620 14670 24795 14685
rect 24810 14705 24840 14710
rect 24810 14670 24840 14675
rect 24620 14535 24635 14670
rect 24870 14655 24885 15525
rect 24915 14680 24930 15595
rect 24680 14640 24885 14655
rect 24900 14675 24930 14680
rect 24900 14640 24930 14645
rect 24680 14535 24695 14640
rect 24960 14625 24975 15665
rect 25005 14650 25020 15735
rect 25855 14710 25870 16015
rect 25885 15980 25925 15985
rect 25885 15950 25890 15980
rect 25920 15950 25925 15980
rect 25885 15945 25925 15950
rect 25855 14705 25885 14710
rect 25855 14670 25885 14675
rect 25900 14685 25915 15945
rect 25945 15910 25985 15915
rect 25945 15880 25950 15910
rect 25980 15880 25985 15910
rect 25945 15875 25985 15880
rect 25945 14740 25960 15875
rect 25975 15840 26015 15845
rect 25975 15810 25980 15840
rect 26010 15810 26015 15840
rect 25975 15805 26015 15810
rect 25945 14735 25975 14740
rect 25945 14700 25975 14705
rect 25990 14715 26005 15805
rect 26035 14770 26050 16155
rect 26065 16120 26105 16125
rect 26065 16090 26070 16120
rect 26100 16090 26105 16120
rect 26065 16085 26105 16090
rect 26035 14765 26065 14770
rect 26035 14730 26065 14735
rect 26080 14745 26095 16085
rect 26125 14800 26140 16295
rect 26155 16260 26195 16265
rect 26155 16230 26160 16260
rect 26190 16230 26195 16260
rect 26155 16225 26195 16230
rect 26995 16225 27000 16255
rect 27030 16225 27035 16255
rect 26125 14795 26155 14800
rect 26125 14760 26155 14765
rect 26170 14775 26185 16225
rect 26805 15065 26845 15070
rect 26805 15035 26810 15065
rect 26840 15035 26845 15065
rect 26805 15030 26845 15035
rect 26880 15030 26885 15060
rect 26915 15030 26920 15060
rect 26270 14995 26310 15000
rect 26270 14965 26275 14995
rect 26305 14965 26310 14995
rect 26270 14960 26310 14965
rect 26170 14760 26255 14775
rect 26080 14730 26195 14745
rect 25990 14700 26135 14715
rect 25900 14670 26075 14685
rect 24740 14610 24975 14625
rect 24990 14645 25020 14650
rect 24990 14610 25020 14615
rect 24740 14535 24755 14610
rect 26060 14535 26075 14670
rect 26120 14535 26135 14700
rect 26180 14535 26195 14730
rect 26240 14535 26255 14760
rect 26270 14570 26305 14960
rect 26810 14575 26845 15030
rect 26905 14575 26920 15030
rect 27005 14775 27020 16225
rect 27050 14800 27065 16295
rect 28620 16300 28625 16330
rect 28655 16300 28660 16330
rect 31115 16330 31155 16335
rect 28620 16295 28660 16300
rect 29520 16295 29525 16325
rect 29555 16295 29560 16325
rect 28530 16190 28570 16195
rect 27115 16155 27120 16185
rect 27150 16155 27155 16185
rect 27085 16085 27090 16115
rect 27120 16085 27125 16115
rect 26805 14570 26845 14575
rect 26270 14540 26275 14570
rect 26305 14540 26310 14570
rect 26270 14535 26310 14540
rect 26805 14540 26810 14570
rect 26840 14540 26845 14570
rect 26805 14535 26845 14540
rect 26890 14570 26920 14575
rect 26890 14535 26920 14540
rect 26935 14760 27020 14775
rect 27035 14795 27065 14800
rect 27035 14760 27065 14765
rect 26935 14535 26950 14760
rect 27095 14745 27110 16085
rect 27140 14770 27155 16155
rect 28530 16160 28535 16190
rect 28565 16160 28570 16190
rect 28530 16155 28570 16160
rect 28350 16050 28390 16055
rect 27295 16015 27300 16045
rect 27330 16015 27335 16045
rect 27265 15945 27270 15975
rect 27300 15945 27305 15975
rect 27205 15875 27210 15905
rect 27240 15875 27245 15905
rect 27175 15805 27180 15835
rect 27210 15805 27215 15835
rect 26995 14730 27110 14745
rect 27125 14765 27155 14770
rect 27125 14730 27155 14735
rect 26995 14535 27010 14730
rect 27185 14715 27200 15805
rect 27230 14740 27245 15875
rect 27055 14700 27200 14715
rect 27215 14735 27245 14740
rect 27215 14700 27245 14705
rect 27055 14535 27070 14700
rect 27275 14685 27290 15945
rect 27320 14710 27335 16015
rect 27115 14670 27290 14685
rect 27305 14705 27335 14710
rect 27305 14670 27335 14675
rect 28350 16020 28355 16050
rect 28385 16020 28390 16050
rect 28350 16015 28390 16020
rect 28350 14710 28365 16015
rect 28380 15980 28420 15985
rect 28380 15950 28385 15980
rect 28415 15950 28420 15980
rect 28380 15945 28420 15950
rect 28350 14705 28380 14710
rect 28350 14670 28380 14675
rect 28395 14685 28410 15945
rect 28440 15910 28480 15915
rect 28440 15880 28445 15910
rect 28475 15880 28480 15910
rect 28440 15875 28480 15880
rect 28440 14740 28455 15875
rect 28470 15840 28510 15845
rect 28470 15810 28475 15840
rect 28505 15810 28510 15840
rect 28470 15805 28510 15810
rect 28440 14735 28470 14740
rect 28440 14700 28470 14705
rect 28485 14715 28500 15805
rect 28530 14770 28545 16155
rect 28560 16120 28600 16125
rect 28560 16090 28565 16120
rect 28595 16090 28600 16120
rect 28560 16085 28600 16090
rect 28530 14765 28560 14770
rect 28530 14730 28560 14735
rect 28575 14745 28590 16085
rect 28620 14800 28635 16295
rect 28650 16260 28690 16265
rect 28650 16230 28655 16260
rect 28685 16230 28690 16260
rect 28650 16225 28690 16230
rect 29490 16225 29495 16255
rect 29525 16225 29530 16255
rect 28620 14795 28650 14800
rect 28620 14760 28650 14765
rect 28665 14775 28680 16225
rect 29300 15065 29340 15070
rect 29300 15035 29305 15065
rect 29335 15035 29340 15065
rect 29300 15030 29340 15035
rect 29375 15030 29380 15060
rect 29410 15030 29415 15060
rect 28765 14995 28805 15000
rect 28765 14965 28770 14995
rect 28800 14965 28805 14995
rect 28765 14960 28805 14965
rect 28665 14760 28750 14775
rect 28575 14730 28690 14745
rect 28485 14700 28630 14715
rect 28395 14670 28570 14685
rect 27115 14535 27130 14670
rect 28555 14535 28570 14670
rect 28615 14535 28630 14700
rect 28675 14535 28690 14730
rect 28735 14535 28750 14760
rect 28765 14570 28800 14960
rect 29305 14575 29340 15030
rect 29400 14575 29415 15030
rect 29500 14775 29515 16225
rect 29545 14800 29560 16295
rect 31115 16300 31120 16330
rect 31150 16300 31155 16330
rect 33610 16330 33650 16335
rect 31115 16295 31155 16300
rect 32015 16295 32020 16325
rect 32050 16295 32055 16325
rect 31025 16190 31065 16195
rect 29610 16155 29615 16185
rect 29645 16155 29650 16185
rect 29580 16085 29585 16115
rect 29615 16085 29620 16115
rect 29300 14570 29340 14575
rect 28765 14540 28770 14570
rect 28800 14540 28805 14570
rect 28765 14535 28805 14540
rect 29300 14540 29305 14570
rect 29335 14540 29340 14570
rect 29300 14535 29340 14540
rect 29385 14570 29415 14575
rect 29385 14535 29415 14540
rect 29430 14760 29515 14775
rect 29530 14795 29560 14800
rect 29530 14760 29560 14765
rect 29430 14535 29445 14760
rect 29590 14745 29605 16085
rect 29635 14770 29650 16155
rect 31025 16160 31030 16190
rect 31060 16160 31065 16190
rect 31025 16155 31065 16160
rect 29790 16015 29795 16045
rect 29825 16015 29830 16045
rect 29760 15945 29765 15975
rect 29795 15945 29800 15975
rect 29700 15875 29705 15905
rect 29735 15875 29740 15905
rect 29670 15805 29675 15835
rect 29705 15805 29710 15835
rect 29490 14730 29605 14745
rect 29620 14765 29650 14770
rect 29620 14730 29650 14735
rect 29490 14535 29505 14730
rect 29680 14715 29695 15805
rect 29725 14740 29740 15875
rect 29550 14700 29695 14715
rect 29710 14735 29740 14740
rect 29710 14700 29740 14705
rect 29550 14535 29565 14700
rect 29770 14685 29785 15945
rect 29815 14710 29830 16015
rect 31025 14770 31040 16155
rect 31055 16120 31095 16125
rect 31055 16090 31060 16120
rect 31090 16090 31095 16120
rect 31055 16085 31095 16090
rect 31025 14765 31055 14770
rect 31025 14730 31055 14735
rect 31070 14745 31085 16085
rect 31115 14800 31130 16295
rect 31145 16260 31185 16265
rect 31145 16230 31150 16260
rect 31180 16230 31185 16260
rect 31145 16225 31185 16230
rect 31985 16225 31990 16255
rect 32020 16225 32025 16255
rect 31115 14795 31145 14800
rect 31115 14760 31145 14765
rect 31160 14775 31175 16225
rect 31795 15065 31835 15070
rect 31795 15035 31800 15065
rect 31830 15035 31835 15065
rect 31795 15030 31835 15035
rect 31870 15030 31875 15060
rect 31905 15030 31910 15060
rect 31260 14995 31300 15000
rect 31260 14965 31265 14995
rect 31295 14965 31300 14995
rect 31260 14960 31300 14965
rect 31160 14760 31245 14775
rect 31070 14730 31185 14745
rect 29610 14670 29785 14685
rect 29800 14705 29830 14710
rect 29800 14670 29830 14675
rect 29610 14535 29625 14670
rect 31170 14535 31185 14730
rect 31230 14535 31245 14760
rect 31260 14570 31295 14960
rect 31800 14575 31835 15030
rect 31895 14575 31910 15030
rect 31995 14775 32010 16225
rect 32040 14800 32055 16295
rect 33610 16300 33615 16330
rect 33645 16300 33650 16330
rect 36105 16330 36145 16335
rect 33610 16295 33650 16300
rect 34510 16295 34515 16325
rect 34545 16295 34550 16325
rect 33520 16190 33560 16195
rect 32105 16155 32110 16185
rect 32140 16155 32145 16185
rect 32075 16085 32080 16115
rect 32110 16085 32115 16115
rect 31795 14570 31835 14575
rect 31260 14540 31265 14570
rect 31295 14540 31300 14570
rect 31260 14535 31300 14540
rect 31795 14540 31800 14570
rect 31830 14540 31835 14570
rect 31795 14535 31835 14540
rect 31880 14570 31910 14575
rect 31880 14535 31910 14540
rect 31925 14760 32010 14775
rect 32025 14795 32055 14800
rect 32025 14760 32055 14765
rect 31925 14535 31940 14760
rect 32085 14745 32100 16085
rect 32130 14770 32145 16155
rect 31985 14730 32100 14745
rect 32115 14765 32145 14770
rect 32115 14730 32145 14735
rect 33520 16160 33525 16190
rect 33555 16160 33560 16190
rect 33520 16155 33560 16160
rect 33520 14770 33535 16155
rect 33550 16120 33590 16125
rect 33550 16090 33555 16120
rect 33585 16090 33590 16120
rect 33550 16085 33590 16090
rect 33520 14765 33550 14770
rect 33520 14730 33550 14735
rect 33565 14745 33580 16085
rect 33610 14800 33625 16295
rect 33640 16260 33680 16265
rect 33640 16230 33645 16260
rect 33675 16230 33680 16260
rect 33640 16225 33680 16230
rect 34480 16225 34485 16255
rect 34515 16225 34520 16255
rect 33610 14795 33640 14800
rect 33610 14760 33640 14765
rect 33655 14775 33670 16225
rect 34290 15065 34330 15070
rect 34290 15035 34295 15065
rect 34325 15035 34330 15065
rect 34290 15030 34330 15035
rect 34365 15030 34370 15060
rect 34400 15030 34405 15060
rect 33755 14995 33795 15000
rect 33755 14965 33760 14995
rect 33790 14965 33795 14995
rect 33755 14960 33795 14965
rect 33655 14760 33740 14775
rect 33565 14730 33680 14745
rect 31985 14535 32000 14730
rect 33665 14535 33680 14730
rect 33725 14535 33740 14760
rect 33755 14570 33790 14960
rect 34295 14575 34330 15030
rect 34390 14575 34405 15030
rect 34490 14775 34505 16225
rect 34535 14800 34550 16295
rect 36105 16300 36110 16330
rect 36140 16300 36145 16330
rect 38600 16330 38640 16335
rect 36105 16295 36145 16300
rect 37005 16295 37010 16325
rect 37040 16295 37045 16325
rect 34600 16155 34605 16185
rect 34635 16155 34640 16185
rect 34570 16085 34575 16115
rect 34605 16085 34610 16115
rect 34290 14570 34330 14575
rect 33755 14540 33760 14570
rect 33790 14540 33795 14570
rect 33755 14535 33795 14540
rect 34290 14540 34295 14570
rect 34325 14540 34330 14570
rect 34290 14535 34330 14540
rect 34375 14570 34405 14575
rect 34375 14535 34405 14540
rect 34420 14760 34505 14775
rect 34520 14795 34550 14800
rect 34520 14760 34550 14765
rect 34420 14535 34435 14760
rect 34580 14745 34595 16085
rect 34625 14770 34640 16155
rect 34480 14730 34595 14745
rect 34610 14765 34640 14770
rect 36105 14800 36120 16295
rect 36135 16260 36175 16265
rect 36135 16230 36140 16260
rect 36170 16230 36175 16260
rect 36135 16225 36175 16230
rect 36975 16225 36980 16255
rect 37010 16225 37015 16255
rect 36105 14795 36135 14800
rect 36105 14760 36135 14765
rect 36150 14775 36165 16225
rect 36785 15065 36825 15070
rect 36785 15035 36790 15065
rect 36820 15035 36825 15065
rect 36785 15030 36825 15035
rect 36860 15030 36865 15060
rect 36895 15030 36900 15060
rect 36250 14995 36290 15000
rect 36250 14965 36255 14995
rect 36285 14965 36290 14995
rect 36250 14960 36290 14965
rect 36150 14760 36235 14775
rect 34610 14730 34640 14735
rect 34480 14535 34495 14730
rect 36220 14535 36235 14760
rect 36250 14570 36285 14960
rect 36790 14575 36825 15030
rect 36885 14575 36900 15030
rect 36985 14775 37000 16225
rect 37030 14800 37045 16295
rect 36785 14570 36825 14575
rect 36250 14540 36255 14570
rect 36285 14540 36290 14570
rect 36250 14535 36290 14540
rect 36785 14540 36790 14570
rect 36820 14540 36825 14570
rect 36785 14535 36825 14540
rect 36870 14570 36900 14575
rect 36870 14535 36900 14540
rect 36915 14760 37000 14775
rect 37015 14795 37045 14800
rect 37015 14760 37045 14765
rect 38600 16300 38605 16330
rect 38635 16300 38640 16330
rect 38600 16295 38640 16300
rect 39500 16295 39505 16325
rect 39535 16295 39540 16325
rect 38600 14800 38615 16295
rect 38630 16260 38670 16265
rect 38630 16230 38635 16260
rect 38665 16230 38670 16260
rect 38630 16225 38670 16230
rect 39470 16225 39475 16255
rect 39505 16225 39510 16255
rect 38600 14795 38630 14800
rect 38600 14760 38630 14765
rect 38645 14775 38660 16225
rect 39280 15065 39320 15070
rect 39280 15035 39285 15065
rect 39315 15035 39320 15065
rect 39280 15030 39320 15035
rect 39355 15030 39360 15060
rect 39390 15030 39395 15060
rect 38745 14995 38785 15000
rect 38745 14965 38750 14995
rect 38780 14965 38785 14995
rect 38745 14960 38785 14965
rect 38645 14760 38730 14775
rect 36915 14535 36930 14760
rect 38715 14535 38730 14760
rect 38745 14570 38780 14960
rect 39285 14575 39320 15030
rect 39380 14575 39395 15030
rect 39480 14775 39495 16225
rect 39525 14800 39540 16295
rect 41640 15065 41680 15070
rect 41640 15035 41645 15065
rect 41675 15035 41680 15065
rect 41640 15030 41680 15035
rect 41715 15030 41720 15060
rect 41750 15030 41755 15060
rect 39280 14570 39320 14575
rect 38745 14540 38750 14570
rect 38780 14540 38785 14570
rect 38745 14535 38785 14540
rect 39280 14540 39285 14570
rect 39315 14540 39320 14570
rect 39280 14535 39320 14540
rect 39365 14570 39395 14575
rect 39365 14535 39395 14540
rect 39410 14760 39495 14775
rect 39510 14795 39540 14800
rect 39510 14760 39540 14765
rect 41105 14995 41145 15000
rect 41105 14965 41110 14995
rect 41140 14965 41145 14995
rect 41105 14960 41145 14965
rect 39410 14535 39425 14760
rect 41105 14570 41140 14960
rect 41645 14575 41680 15030
rect 41740 14575 41755 15030
rect 41640 14570 41680 14575
rect 41105 14540 41110 14570
rect 41140 14540 41145 14570
rect 41105 14535 41145 14540
rect 41640 14540 41645 14570
rect 41675 14540 41680 14570
rect 41640 14535 41680 14540
rect 41725 14570 41755 14575
rect 41725 14535 41755 14540
rect -635 14495 -630 14535
rect -590 14495 -585 14535
rect -635 14490 -585 14495
rect 22185 13665 22200 13680
rect -2395 -870 -2375 0
rect -2395 -875 -1170 -870
rect -2395 -885 -1205 -875
rect -1210 -905 -1205 -885
rect -1175 -905 -1170 -875
rect -1210 -910 -1170 -905
<< via2 >>
rect 1180 16300 1210 16330
rect -2755 15030 -2725 15060
rect -500 15035 -470 15065
rect -2620 14965 -2590 14995
rect -2550 14965 -2520 14995
rect -1035 14965 -1005 14995
rect -2680 14895 -2650 14925
rect 1210 16230 1240 16260
rect 1860 15035 1890 15065
rect 1325 14965 1355 14995
rect 3675 16300 3705 16330
rect 3705 16230 3735 16260
rect 4355 15035 4385 15065
rect 3820 14965 3850 14995
rect 6170 16300 6200 16330
rect 6080 16160 6110 16190
rect 6110 16090 6140 16120
rect 6200 16230 6230 16260
rect 6850 15035 6880 15065
rect 6315 14965 6345 14995
rect 8665 16300 8695 16330
rect 8575 16160 8605 16190
rect 8605 16090 8635 16120
rect 8695 16230 8725 16260
rect 9345 15035 9375 15065
rect 8810 14965 8840 14995
rect 11160 16300 11190 16330
rect 11070 16160 11100 16190
rect 10890 16020 10920 16050
rect 10920 15950 10950 15980
rect 10980 15880 11010 15910
rect 11010 15810 11040 15840
rect 11100 16090 11130 16120
rect 11190 16230 11220 16260
rect 11840 15035 11870 15065
rect 11305 14965 11335 14995
rect 13655 16300 13685 16330
rect 13565 16160 13595 16190
rect 13385 16020 13415 16050
rect 13415 15950 13445 15980
rect 13475 15880 13505 15910
rect 13505 15810 13535 15840
rect 13595 16090 13625 16120
rect 13685 16230 13715 16260
rect 14335 15035 14365 15065
rect 13800 14965 13830 14995
rect 16150 16300 16180 16330
rect 16060 16160 16090 16190
rect 15970 16020 16000 16050
rect 15880 15880 15910 15910
rect 15700 15740 15730 15770
rect 15730 15670 15760 15700
rect 15790 15600 15820 15630
rect 15820 15530 15850 15560
rect 15910 15810 15940 15840
rect 16000 15950 16030 15980
rect 16090 16090 16120 16120
rect 16180 16230 16210 16260
rect 16830 15035 16860 15065
rect 16295 14965 16325 14995
rect 18645 16300 18675 16330
rect 18555 16160 18585 16190
rect 18465 16020 18495 16050
rect 18375 15880 18405 15910
rect 18285 15740 18315 15770
rect 18195 15460 18225 15490
rect 18105 15180 18135 15210
rect 18135 15110 18165 15140
rect 18225 15390 18255 15420
rect 18315 15670 18345 15700
rect 18405 15810 18435 15840
rect 18495 15950 18525 15980
rect 18585 16090 18615 16120
rect 18675 16230 18705 16260
rect 19325 15035 19355 15065
rect 18790 14965 18820 14995
rect 21140 16300 21170 16330
rect 21050 16160 21080 16190
rect 20960 16020 20990 16050
rect 20870 15880 20900 15910
rect 20780 15740 20810 15770
rect 20600 15460 20630 15490
rect 20630 15390 20660 15420
rect 20675 15320 20705 15350
rect 20720 15250 20750 15280
rect 20810 15670 20840 15700
rect 20900 15810 20930 15840
rect 20990 15950 21020 15980
rect 21080 16090 21110 16120
rect 21170 16230 21200 16260
rect 21820 15035 21850 15065
rect 21285 14965 21315 14995
rect 23635 16300 23665 16330
rect 23545 16160 23575 16190
rect 23455 16020 23485 16050
rect 23365 15880 23395 15910
rect 23185 15740 23215 15770
rect 23215 15670 23245 15700
rect 23275 15600 23305 15630
rect 23305 15530 23335 15560
rect 23395 15810 23425 15840
rect 23485 15950 23515 15980
rect 23575 16090 23605 16120
rect 23665 16230 23695 16260
rect 24315 15035 24345 15065
rect 23780 14965 23810 14995
rect 26130 16300 26160 16330
rect 26040 16160 26070 16190
rect 25860 16020 25890 16050
rect 25890 15950 25920 15980
rect 25950 15880 25980 15910
rect 25980 15810 26010 15840
rect 26070 16090 26100 16120
rect 26160 16230 26190 16260
rect 26810 15035 26840 15065
rect 26275 14965 26305 14995
rect 28625 16300 28655 16330
rect 28535 16160 28565 16190
rect 28355 16020 28385 16050
rect 28385 15950 28415 15980
rect 28445 15880 28475 15910
rect 28475 15810 28505 15840
rect 28565 16090 28595 16120
rect 28655 16230 28685 16260
rect 29305 15035 29335 15065
rect 28770 14965 28800 14995
rect 31120 16300 31150 16330
rect 31030 16160 31060 16190
rect 31060 16090 31090 16120
rect 31150 16230 31180 16260
rect 31800 15035 31830 15065
rect 31265 14965 31295 14995
rect 33615 16300 33645 16330
rect 33525 16160 33555 16190
rect 33555 16090 33585 16120
rect 33645 16230 33675 16260
rect 34295 15035 34325 15065
rect 33760 14965 33790 14995
rect 36110 16300 36140 16330
rect 36140 16230 36170 16260
rect 36790 15035 36820 15065
rect 36255 14965 36285 14995
rect 38605 16300 38635 16330
rect 38635 16230 38665 16260
rect 39285 15035 39315 15065
rect 38750 14965 38780 14995
rect 41645 15035 41675 15065
rect 41110 14965 41140 14995
rect -630 14495 -590 14535
rect -1205 -905 -1175 -875
<< metal3 >>
rect 1175 16330 1215 16335
rect 1175 16325 1180 16330
rect -2570 16300 1180 16325
rect 1210 16325 1215 16330
rect 3670 16330 3710 16335
rect 3670 16325 3675 16330
rect 1210 16300 3675 16325
rect 3705 16325 3710 16330
rect 6165 16330 6205 16335
rect 6165 16325 6170 16330
rect 3705 16300 6170 16325
rect 6200 16325 6205 16330
rect 8660 16330 8700 16335
rect 8660 16325 8665 16330
rect 6200 16300 8665 16325
rect 8695 16325 8700 16330
rect 11155 16330 11195 16335
rect 11155 16325 11160 16330
rect 8695 16300 11160 16325
rect 11190 16325 11195 16330
rect 13650 16330 13690 16335
rect 13650 16325 13655 16330
rect 11190 16300 13655 16325
rect 13685 16325 13690 16330
rect 16145 16330 16185 16335
rect 16145 16325 16150 16330
rect 13685 16300 16150 16325
rect 16180 16325 16185 16330
rect 18640 16330 18680 16335
rect 18640 16325 18645 16330
rect 16180 16300 18645 16325
rect 18675 16325 18680 16330
rect 21135 16330 21175 16335
rect 21135 16325 21140 16330
rect 18675 16300 21140 16325
rect 21170 16325 21175 16330
rect 23630 16330 23670 16335
rect 23630 16325 23635 16330
rect 21170 16300 23635 16325
rect 23665 16325 23670 16330
rect 26125 16330 26165 16335
rect 26125 16325 26130 16330
rect 23665 16300 26130 16325
rect 26160 16325 26165 16330
rect 28620 16330 28660 16335
rect 28620 16325 28625 16330
rect 26160 16300 28625 16325
rect 28655 16325 28660 16330
rect 31115 16330 31155 16335
rect 31115 16325 31120 16330
rect 28655 16300 31120 16325
rect 31150 16325 31155 16330
rect 33610 16330 33650 16335
rect 33610 16325 33615 16330
rect 31150 16300 33615 16325
rect 33645 16325 33650 16330
rect 36105 16330 36145 16335
rect 36105 16325 36110 16330
rect 33645 16300 36110 16325
rect 36140 16325 36145 16330
rect 38600 16330 38640 16335
rect 38600 16325 38605 16330
rect 36140 16300 38605 16325
rect 38635 16325 38640 16330
rect 38635 16300 42325 16325
rect -2570 16295 42325 16300
rect 1205 16260 1245 16265
rect 1205 16255 1210 16260
rect -2570 16230 1210 16255
rect 1240 16255 1245 16260
rect 3700 16260 3740 16265
rect 3700 16255 3705 16260
rect 1240 16230 3705 16255
rect 3735 16255 3740 16260
rect 6195 16260 6235 16265
rect 6195 16255 6200 16260
rect 3735 16230 6200 16255
rect 6230 16255 6235 16260
rect 8690 16260 8730 16265
rect 8690 16255 8695 16260
rect 6230 16230 8695 16255
rect 8725 16255 8730 16260
rect 11185 16260 11225 16265
rect 11185 16255 11190 16260
rect 8725 16230 11190 16255
rect 11220 16255 11225 16260
rect 13680 16260 13720 16265
rect 13680 16255 13685 16260
rect 11220 16230 13685 16255
rect 13715 16255 13720 16260
rect 16175 16260 16215 16265
rect 16175 16255 16180 16260
rect 13715 16230 16180 16255
rect 16210 16255 16215 16260
rect 18670 16260 18710 16265
rect 18670 16255 18675 16260
rect 16210 16230 18675 16255
rect 18705 16255 18710 16260
rect 21165 16260 21205 16265
rect 21165 16255 21170 16260
rect 18705 16230 21170 16255
rect 21200 16255 21205 16260
rect 23660 16260 23700 16265
rect 23660 16255 23665 16260
rect 21200 16230 23665 16255
rect 23695 16255 23700 16260
rect 26155 16260 26195 16265
rect 26155 16255 26160 16260
rect 23695 16230 26160 16255
rect 26190 16255 26195 16260
rect 28650 16260 28690 16265
rect 28650 16255 28655 16260
rect 26190 16230 28655 16255
rect 28685 16255 28690 16260
rect 31145 16260 31185 16265
rect 31145 16255 31150 16260
rect 28685 16230 31150 16255
rect 31180 16255 31185 16260
rect 33640 16260 33680 16265
rect 33640 16255 33645 16260
rect 31180 16230 33645 16255
rect 33675 16255 33680 16260
rect 36135 16260 36175 16265
rect 36135 16255 36140 16260
rect 33675 16230 36140 16255
rect 36170 16255 36175 16260
rect 38630 16260 38670 16265
rect 38630 16255 38635 16260
rect 36170 16230 38635 16255
rect 38665 16255 38670 16260
rect 38665 16230 42325 16255
rect -2570 16225 42325 16230
rect 6075 16190 6115 16195
rect 6075 16185 6080 16190
rect -2570 16160 6080 16185
rect 6110 16185 6115 16190
rect 8570 16190 8610 16195
rect 8570 16185 8575 16190
rect 6110 16160 8575 16185
rect 8605 16185 8610 16190
rect 11065 16190 11105 16195
rect 11065 16185 11070 16190
rect 8605 16160 11070 16185
rect 11100 16185 11105 16190
rect 13560 16190 13600 16195
rect 13560 16185 13565 16190
rect 11100 16160 13565 16185
rect 13595 16185 13600 16190
rect 16055 16190 16095 16195
rect 16055 16185 16060 16190
rect 13595 16160 16060 16185
rect 16090 16185 16095 16190
rect 18550 16190 18590 16195
rect 18550 16185 18555 16190
rect 16090 16160 18555 16185
rect 18585 16185 18590 16190
rect 21045 16190 21085 16195
rect 21045 16185 21050 16190
rect 18585 16160 21050 16185
rect 21080 16185 21085 16190
rect 23540 16190 23580 16195
rect 23540 16185 23545 16190
rect 21080 16160 23545 16185
rect 23575 16185 23580 16190
rect 26035 16190 26075 16195
rect 26035 16185 26040 16190
rect 23575 16160 26040 16185
rect 26070 16185 26075 16190
rect 28530 16190 28570 16195
rect 28530 16185 28535 16190
rect 26070 16160 28535 16185
rect 28565 16185 28570 16190
rect 31025 16190 31065 16195
rect 31025 16185 31030 16190
rect 28565 16160 31030 16185
rect 31060 16185 31065 16190
rect 33520 16190 33560 16195
rect 33520 16185 33525 16190
rect 31060 16160 33525 16185
rect 33555 16185 33560 16190
rect 33555 16160 42325 16185
rect -2570 16155 42325 16160
rect 6105 16120 6145 16125
rect 6105 16115 6110 16120
rect -2570 16090 6110 16115
rect 6140 16115 6145 16120
rect 8600 16120 8640 16125
rect 8600 16115 8605 16120
rect 6140 16090 8605 16115
rect 8635 16115 8640 16120
rect 11095 16120 11135 16125
rect 11095 16115 11100 16120
rect 8635 16090 11100 16115
rect 11130 16115 11135 16120
rect 13590 16120 13630 16125
rect 13590 16115 13595 16120
rect 11130 16090 13595 16115
rect 13625 16115 13630 16120
rect 16085 16120 16125 16125
rect 16085 16115 16090 16120
rect 13625 16090 16090 16115
rect 16120 16115 16125 16120
rect 18580 16120 18620 16125
rect 18580 16115 18585 16120
rect 16120 16090 18585 16115
rect 18615 16115 18620 16120
rect 21075 16120 21115 16125
rect 21075 16115 21080 16120
rect 18615 16090 21080 16115
rect 21110 16115 21115 16120
rect 23570 16120 23610 16125
rect 23570 16115 23575 16120
rect 21110 16090 23575 16115
rect 23605 16115 23610 16120
rect 26065 16120 26105 16125
rect 26065 16115 26070 16120
rect 23605 16090 26070 16115
rect 26100 16115 26105 16120
rect 28560 16120 28600 16125
rect 28560 16115 28565 16120
rect 26100 16090 28565 16115
rect 28595 16115 28600 16120
rect 31055 16120 31095 16125
rect 31055 16115 31060 16120
rect 28595 16090 31060 16115
rect 31090 16115 31095 16120
rect 33550 16120 33590 16125
rect 33550 16115 33555 16120
rect 31090 16090 33555 16115
rect 33585 16115 33590 16120
rect 33585 16090 42325 16115
rect -2570 16085 42325 16090
rect 10885 16050 10925 16055
rect 10885 16045 10890 16050
rect -2570 16020 10890 16045
rect 10920 16045 10925 16050
rect 13380 16050 13420 16055
rect 13380 16045 13385 16050
rect 10920 16020 13385 16045
rect 13415 16045 13420 16050
rect 15965 16050 16005 16055
rect 15965 16045 15970 16050
rect 13415 16020 15970 16045
rect 16000 16045 16005 16050
rect 18460 16050 18500 16055
rect 18460 16045 18465 16050
rect 16000 16020 18465 16045
rect 18495 16045 18500 16050
rect 20955 16050 20995 16055
rect 20955 16045 20960 16050
rect 18495 16020 20960 16045
rect 20990 16045 20995 16050
rect 23450 16050 23490 16055
rect 23450 16045 23455 16050
rect 20990 16020 23455 16045
rect 23485 16045 23490 16050
rect 25855 16050 25895 16055
rect 25855 16045 25860 16050
rect 23485 16020 25860 16045
rect 25890 16045 25895 16050
rect 28350 16050 28390 16055
rect 28350 16045 28355 16050
rect 25890 16020 28355 16045
rect 28385 16045 28390 16050
rect 28385 16020 42325 16045
rect -2570 16015 42325 16020
rect 10915 15980 10955 15985
rect 10915 15975 10920 15980
rect -2570 15950 10920 15975
rect 10950 15975 10955 15980
rect 13410 15980 13450 15985
rect 13410 15975 13415 15980
rect 10950 15950 13415 15975
rect 13445 15975 13450 15980
rect 15995 15980 16035 15985
rect 15995 15975 16000 15980
rect 13445 15950 16000 15975
rect 16030 15975 16035 15980
rect 18490 15980 18530 15985
rect 18490 15975 18495 15980
rect 16030 15950 18495 15975
rect 18525 15975 18530 15980
rect 20985 15980 21025 15985
rect 20985 15975 20990 15980
rect 18525 15950 20990 15975
rect 21020 15975 21025 15980
rect 23480 15980 23520 15985
rect 23480 15975 23485 15980
rect 21020 15950 23485 15975
rect 23515 15975 23520 15980
rect 25885 15980 25925 15985
rect 25885 15975 25890 15980
rect 23515 15950 25890 15975
rect 25920 15975 25925 15980
rect 28380 15980 28420 15985
rect 28380 15975 28385 15980
rect 25920 15950 28385 15975
rect 28415 15975 28420 15980
rect 28415 15950 42325 15975
rect -2570 15945 42325 15950
rect 10975 15910 11015 15915
rect 10975 15905 10980 15910
rect -2570 15880 10980 15905
rect 11010 15905 11015 15910
rect 13470 15910 13510 15915
rect 13470 15905 13475 15910
rect 11010 15880 13475 15905
rect 13505 15905 13510 15910
rect 15875 15910 15915 15915
rect 15875 15905 15880 15910
rect 13505 15880 15880 15905
rect 15910 15905 15915 15910
rect 18370 15910 18410 15915
rect 18370 15905 18375 15910
rect 15910 15880 18375 15905
rect 18405 15905 18410 15910
rect 20865 15910 20905 15915
rect 20865 15905 20870 15910
rect 18405 15880 20870 15905
rect 20900 15905 20905 15910
rect 23360 15910 23400 15915
rect 23360 15905 23365 15910
rect 20900 15880 23365 15905
rect 23395 15905 23400 15910
rect 25945 15910 25985 15915
rect 25945 15905 25950 15910
rect 23395 15880 25950 15905
rect 25980 15905 25985 15910
rect 28440 15910 28480 15915
rect 28440 15905 28445 15910
rect 25980 15880 28445 15905
rect 28475 15905 28480 15910
rect 28475 15880 42325 15905
rect -2570 15875 42325 15880
rect 11005 15840 11045 15845
rect 11005 15835 11010 15840
rect -2570 15810 11010 15835
rect 11040 15835 11045 15840
rect 13500 15840 13540 15845
rect 13500 15835 13505 15840
rect 11040 15810 13505 15835
rect 13535 15835 13540 15840
rect 15905 15840 15945 15845
rect 15905 15835 15910 15840
rect 13535 15810 15910 15835
rect 15940 15835 15945 15840
rect 18400 15840 18440 15845
rect 18400 15835 18405 15840
rect 15940 15810 18405 15835
rect 18435 15835 18440 15840
rect 20895 15840 20935 15845
rect 20895 15835 20900 15840
rect 18435 15810 20900 15835
rect 20930 15835 20935 15840
rect 23390 15840 23430 15845
rect 23390 15835 23395 15840
rect 20930 15810 23395 15835
rect 23425 15835 23430 15840
rect 25975 15840 26015 15845
rect 25975 15835 25980 15840
rect 23425 15810 25980 15835
rect 26010 15835 26015 15840
rect 28470 15840 28510 15845
rect 28470 15835 28475 15840
rect 26010 15810 28475 15835
rect 28505 15835 28510 15840
rect 28505 15810 42325 15835
rect -2570 15805 42325 15810
rect 15695 15770 15735 15775
rect 15695 15765 15700 15770
rect -2570 15740 15700 15765
rect 15730 15765 15735 15770
rect 18280 15770 18320 15775
rect 18280 15765 18285 15770
rect 15730 15740 18285 15765
rect 18315 15765 18320 15770
rect 20775 15770 20815 15775
rect 20775 15765 20780 15770
rect 18315 15740 20780 15765
rect 20810 15765 20815 15770
rect 23180 15770 23220 15775
rect 23180 15765 23185 15770
rect 20810 15740 23185 15765
rect 23215 15765 23220 15770
rect 23215 15740 42325 15765
rect -2570 15735 42325 15740
rect 15725 15700 15765 15705
rect 15725 15695 15730 15700
rect -2570 15670 15730 15695
rect 15760 15695 15765 15700
rect 18310 15700 18350 15705
rect 18310 15695 18315 15700
rect 15760 15670 18315 15695
rect 18345 15695 18350 15700
rect 20805 15700 20845 15705
rect 20805 15695 20810 15700
rect 18345 15670 20810 15695
rect 20840 15695 20845 15700
rect 23210 15700 23250 15705
rect 23210 15695 23215 15700
rect 20840 15670 23215 15695
rect 23245 15695 23250 15700
rect 23245 15670 42325 15695
rect -2570 15665 42325 15670
rect 15785 15630 15825 15635
rect 15785 15625 15790 15630
rect -2570 15600 15790 15625
rect 15820 15625 15825 15630
rect 23270 15630 23310 15635
rect 23270 15625 23275 15630
rect 15820 15600 23275 15625
rect 23305 15625 23310 15630
rect 23305 15600 42325 15625
rect -2570 15595 42325 15600
rect 15815 15560 15855 15565
rect 15815 15555 15820 15560
rect -2570 15530 15820 15555
rect 15850 15555 15855 15560
rect 23300 15560 23340 15565
rect 23300 15555 23305 15560
rect 15850 15530 23305 15555
rect 23335 15555 23340 15560
rect 23335 15530 42325 15555
rect -2570 15525 42325 15530
rect 18190 15490 18230 15495
rect 18190 15485 18195 15490
rect -2570 15460 18195 15485
rect 18225 15485 18230 15490
rect 20595 15490 20635 15495
rect 20595 15485 20600 15490
rect 18225 15460 20600 15485
rect 20630 15485 20635 15490
rect 20630 15460 42325 15485
rect -2570 15455 42325 15460
rect 18220 15420 18260 15425
rect 18220 15415 18225 15420
rect -2570 15390 18225 15415
rect 18255 15415 18260 15420
rect 20625 15420 20665 15425
rect 20625 15415 20630 15420
rect 18255 15390 20630 15415
rect 20660 15415 20665 15420
rect 20660 15390 42325 15415
rect -2570 15385 42325 15390
rect 20670 15350 20710 15355
rect 20670 15345 20675 15350
rect -2570 15320 20675 15345
rect 20705 15345 20710 15350
rect 20705 15320 42325 15345
rect -2570 15315 42325 15320
rect 20715 15280 20755 15285
rect 20715 15275 20720 15280
rect -2570 15250 20720 15275
rect 20750 15275 20755 15280
rect 20750 15250 42325 15275
rect -2570 15245 42325 15250
rect 18100 15210 18140 15215
rect 18100 15205 18105 15210
rect -2590 15200 18105 15205
rect -2790 15180 18105 15200
rect 18135 15205 18140 15210
rect 18135 15180 42325 15205
rect -2790 15175 42325 15180
rect -2790 15170 -2570 15175
rect 18130 15140 18170 15145
rect 18130 15135 18135 15140
rect -2590 15130 18135 15135
rect -2790 15110 18135 15130
rect 18165 15135 18170 15140
rect 18165 15110 42325 15135
rect -2790 15105 42325 15110
rect -2790 15100 -2570 15105
rect -2765 15065 -2715 15070
rect -2765 15025 -2760 15065
rect -2720 15025 -2715 15065
rect -505 15065 -465 15070
rect -505 15060 -500 15065
rect -2765 15020 -2715 15025
rect -2685 15035 -500 15060
rect -470 15060 -465 15065
rect 1855 15065 1895 15070
rect 1855 15060 1860 15065
rect -470 15035 1860 15060
rect 1890 15060 1895 15065
rect 4350 15065 4390 15070
rect 4350 15060 4355 15065
rect 1890 15035 4355 15060
rect 4385 15060 4390 15065
rect 6845 15065 6885 15070
rect 6845 15060 6850 15065
rect 4385 15035 6850 15060
rect 6880 15060 6885 15065
rect 9340 15065 9380 15070
rect 9340 15060 9345 15065
rect 6880 15035 9345 15060
rect 9375 15060 9380 15065
rect 11835 15065 11875 15070
rect 11835 15060 11840 15065
rect 9375 15035 11840 15060
rect 11870 15060 11875 15065
rect 14330 15065 14370 15070
rect 14330 15060 14335 15065
rect 11870 15035 14335 15060
rect 14365 15060 14370 15065
rect 16825 15065 16865 15070
rect 16825 15060 16830 15065
rect 14365 15035 16830 15060
rect 16860 15060 16865 15065
rect 19320 15065 19360 15070
rect 19320 15060 19325 15065
rect 16860 15035 19325 15060
rect 19355 15060 19360 15065
rect 21815 15065 21855 15070
rect 21815 15060 21820 15065
rect 19355 15035 21820 15060
rect 21850 15060 21855 15065
rect 24310 15065 24350 15070
rect 24310 15060 24315 15065
rect 21850 15035 24315 15060
rect 24345 15060 24350 15065
rect 26805 15065 26845 15070
rect 26805 15060 26810 15065
rect 24345 15035 26810 15060
rect 26840 15060 26845 15065
rect 29300 15065 29340 15070
rect 29300 15060 29305 15065
rect 26840 15035 29305 15060
rect 29335 15060 29340 15065
rect 31795 15065 31835 15070
rect 31795 15060 31800 15065
rect 29335 15035 31800 15060
rect 31830 15060 31835 15065
rect 34290 15065 34330 15070
rect 34290 15060 34295 15065
rect 31830 15035 34295 15060
rect 34325 15060 34330 15065
rect 36785 15065 36825 15070
rect 36785 15060 36790 15065
rect 34325 15035 36790 15060
rect 36820 15060 36825 15065
rect 39280 15065 39320 15070
rect 39280 15060 39285 15065
rect 36820 15035 39285 15060
rect 39315 15060 39320 15065
rect 41640 15065 41680 15070
rect 41640 15060 41645 15065
rect 39315 15035 41645 15060
rect 41675 15060 41680 15065
rect 41675 15035 42325 15060
rect -2685 15030 42325 15035
rect -3185 14950 -3150 14995
rect -2685 14930 -2655 15030
rect -2625 14995 -2585 15000
rect -2625 14965 -2620 14995
rect -2590 14990 -2585 14995
rect -2555 14995 -2515 15000
rect -2555 14990 -2550 14995
rect -2590 14965 -2550 14990
rect -2520 14990 -2515 14995
rect -1040 14995 -1000 15000
rect -1040 14990 -1035 14995
rect -2520 14965 -1035 14990
rect -1005 14990 -1000 14995
rect 1320 14995 1360 15000
rect 1320 14990 1325 14995
rect -1005 14965 1325 14990
rect 1355 14990 1360 14995
rect 3815 14995 3855 15000
rect 3815 14990 3820 14995
rect 1355 14965 3820 14990
rect 3850 14990 3855 14995
rect 6310 14995 6350 15000
rect 6310 14990 6315 14995
rect 3850 14965 6315 14990
rect 6345 14990 6350 14995
rect 8805 14995 8845 15000
rect 8805 14990 8810 14995
rect 6345 14965 8810 14990
rect 8840 14990 8845 14995
rect 11300 14995 11340 15000
rect 11300 14990 11305 14995
rect 8840 14965 11305 14990
rect 11335 14990 11340 14995
rect 13795 14995 13835 15000
rect 13795 14990 13800 14995
rect 11335 14965 13800 14990
rect 13830 14990 13835 14995
rect 16290 14995 16330 15000
rect 16290 14990 16295 14995
rect 13830 14965 16295 14990
rect 16325 14990 16330 14995
rect 18785 14995 18825 15000
rect 18785 14990 18790 14995
rect 16325 14965 18790 14990
rect 18820 14990 18825 14995
rect 21280 14995 21320 15000
rect 21280 14990 21285 14995
rect 18820 14965 21285 14990
rect 21315 14990 21320 14995
rect 23775 14995 23815 15000
rect 23775 14990 23780 14995
rect 21315 14965 23780 14990
rect 23810 14990 23815 14995
rect 26270 14995 26310 15000
rect 26270 14990 26275 14995
rect 23810 14965 26275 14990
rect 26305 14990 26310 14995
rect 28765 14995 28805 15000
rect 28765 14990 28770 14995
rect 26305 14965 28770 14990
rect 28800 14990 28805 14995
rect 31260 14995 31300 15000
rect 31260 14990 31265 14995
rect 28800 14965 31265 14990
rect 31295 14990 31300 14995
rect 33755 14995 33795 15000
rect 33755 14990 33760 14995
rect 31295 14965 33760 14990
rect 33790 14990 33795 14995
rect 36250 14995 36290 15000
rect 36250 14990 36255 14995
rect 33790 14965 36255 14990
rect 36285 14990 36290 14995
rect 38745 14995 38785 15000
rect 38745 14990 38750 14995
rect 36285 14965 38750 14990
rect 38780 14990 38785 14995
rect 41105 14995 41145 15000
rect 41105 14990 41110 14995
rect 38780 14965 41110 14990
rect 41140 14990 41145 14995
rect 41140 14965 42325 14990
rect -2625 14960 42325 14965
rect -2685 14925 -2645 14930
rect -2685 14895 -2680 14925
rect -2650 14895 -2645 14925
rect -2685 14890 -2645 14895
rect -635 14535 -585 14540
rect -635 14495 -630 14535
rect -590 14495 -585 14535
rect -635 14490 -585 14495
rect -1215 40 -1165 45
rect -1215 0 -1210 40
rect -1170 0 -1165 40
rect -1215 -5 -1165 0
rect 38490 35 38540 40
rect 38490 -5 38495 35
rect 38535 -5 38540 35
rect -1205 -870 -1175 -5
rect 38490 -10 38540 -5
rect -1210 -875 -1170 -870
rect -1210 -905 -1205 -875
rect -1175 -905 -1170 -875
rect -1210 -910 -1170 -905
rect 38500 -935 38530 -10
<< via3 >>
rect -2760 15060 -2720 15065
rect -2760 15030 -2755 15060
rect -2755 15030 -2725 15060
rect -2725 15030 -2720 15060
rect -2760 15025 -2720 15030
rect -630 14495 -590 14535
rect -1210 0 -1170 40
rect 38495 -5 38535 35
<< metal4 >>
rect -2765 15065 -2715 15070
rect -2765 15025 -2760 15065
rect -2720 15025 -2715 15065
rect -3185 14995 -2715 15025
rect -3185 14950 -3150 14995
rect -2845 14775 -2795 14805
rect -2320 14535 39855 14540
rect -2320 14510 -630 14535
rect -2320 -825 -2290 14510
rect -635 14495 -630 14510
rect -590 14510 39855 14535
rect -590 14495 -585 14510
rect -635 14490 -585 14495
rect 40 14440 70 14510
rect 2535 14440 2565 14510
rect 5030 14440 5060 14510
rect 7525 14440 7555 14510
rect 10020 14440 10050 14510
rect 12515 14440 12545 14510
rect 15010 14440 15040 14510
rect 17505 14440 17535 14510
rect 20000 14440 20030 14510
rect 22495 14440 22525 14510
rect 24990 14440 25020 14510
rect 27485 14440 27515 14510
rect 29980 14440 30010 14510
rect 32475 14440 32505 14510
rect 34970 14440 35000 14510
rect 37465 14440 37495 14510
rect -1215 40 -1165 45
rect -1215 0 -1210 40
rect -1170 30 -1165 40
rect 38490 35 38540 40
rect 38490 30 38495 35
rect -1170 0 38495 30
rect -1215 -5 -1165 0
rect 38490 -5 38495 0
rect 38535 -5 38540 35
rect 38490 -10 38540 -5
rect 40 -825 70 -755
rect 2535 -825 2565 -755
rect 5030 -825 5060 -755
rect 7525 -825 7555 -755
rect 10020 -825 10050 -755
rect 12515 -825 12545 -755
rect 15010 -825 15040 -755
rect 17505 -825 17535 -755
rect 20000 -825 20030 -755
rect 22495 -825 22525 -755
rect 24990 -825 25020 -755
rect 27485 -825 27515 -755
rect 29980 -825 30010 -755
rect 32475 -825 32505 -755
rect 34970 -825 35000 -755
rect 37465 -825 37495 -755
rect 39825 -825 39855 14510
rect -2320 -855 39855 -825
use dum_vert  cap_dum_0
timestamp 1730644682
transform 0 1 9280 -1 0 14670
box 135 -1795 990 565
use dum_vert  cap_dum_1
timestamp 1730644682
transform 0 1 21755 -1 0 14670
box 135 -1795 990 565
use dum_vert  cap_dum_2
timestamp 1730644682
transform 0 1 24250 -1 0 14670
box 135 -1795 990 565
use dum_vert  cap_dum_3
timestamp 1730644682
transform 0 1 26745 -1 0 14670
box 135 -1795 990 565
use dum_vert  cap_dum_4
timestamp 1730644682
transform 0 1 29240 -1 0 14670
box 135 -1795 990 565
use dum_vert  cap_dum_5
timestamp 1730644682
transform 0 1 31735 -1 0 14670
box 135 -1795 990 565
use dum_vert  cap_dum_6
timestamp 1730644682
transform 0 1 34230 -1 0 14670
box 135 -1795 990 565
use dum_vert  cap_dum_7
timestamp 1730644682
transform 0 1 36725 -1 0 14670
box 135 -1795 990 565
use dum_vert  cap_dum_8
timestamp 1730644682
transform 0 1 39220 -1 0 14670
box 135 -1795 990 565
use dum_vert  cap_dum_10
timestamp 1730644682
transform 0 1 4290 -1 0 14670
box 135 -1795 990 565
use dum_vert  cap_dum_11
timestamp 1730644682
transform 0 1 6785 -1 0 14670
box 135 -1795 990 565
use dum_vert  cap_dum_12
timestamp 1730644682
transform 0 1 19260 -1 0 14670
box 135 -1795 990 565
use dum_vert  cap_dum_13
timestamp 1730644682
transform 0 1 11775 -1 0 14670
box 135 -1795 990 565
use dum_vert  cap_dum_14
timestamp 1730644682
transform 0 1 14270 -1 0 14670
box 135 -1795 990 565
use dum_vert  cap_dum_15
timestamp 1730644682
transform 0 1 16765 -1 0 14670
box 135 -1795 990 565
use dum_vert  dum_vert_0
timestamp 1730644682
transform 0 1 -565 -1 0 990
box 135 -1795 990 565
use dum_vert  dum_vert_1
timestamp 1730644682
transform 0 1 1795 -1 0 14670
box 135 -1795 990 565
use dum_vert  dum_vert_2
timestamp 1730644682
transform 0 1 -565 -1 0 14670
box 135 -1795 990 565
use dum_vert  dum_vert_3
timestamp 1730644682
transform 0 1 -565 -1 0 13815
box 135 -1795 990 565
use dum_vert  dum_vert_4
timestamp 1730644682
transform 0 1 -565 -1 0 12960
box 135 -1795 990 565
use dum_vert  dum_vert_5
timestamp 1730644682
transform 0 1 -565 -1 0 12105
box 135 -1795 990 565
use dum_vert  dum_vert_6
timestamp 1730644682
transform 0 1 -565 -1 0 11250
box 135 -1795 990 565
use dum_vert  dum_vert_7
timestamp 1730644682
transform 0 1 -565 -1 0 10395
box 135 -1795 990 565
use dum_vert  dum_vert_8
timestamp 1730644682
transform 0 1 -565 -1 0 9540
box 135 -1795 990 565
use dum_vert  dum_vert_9
timestamp 1730644682
transform 0 1 -565 -1 0 8685
box 135 -1795 990 565
use dum_vert  dum_vert_10
timestamp 1730644682
transform 0 1 -565 -1 0 7830
box 135 -1795 990 565
use dum_vert  dum_vert_11
timestamp 1730644682
transform 0 1 -565 -1 0 6975
box 135 -1795 990 565
use dum_vert  dum_vert_12
timestamp 1730644682
transform 0 1 -565 -1 0 6120
box 135 -1795 990 565
use dum_vert  dum_vert_13
timestamp 1730644682
transform 0 1 -565 -1 0 5265
box 135 -1795 990 565
use dum_vert  dum_vert_14
timestamp 1730644682
transform 0 1 -565 -1 0 4410
box 135 -1795 990 565
use dum_vert  dum_vert_15
timestamp 1730644682
transform 0 1 -565 -1 0 3555
box 135 -1795 990 565
use dum_vert  dum_vert_16
timestamp 1730644682
transform 0 1 -565 -1 0 2700
box 135 -1795 990 565
use dum_vert  dum_vert_17
timestamp 1730644682
transform 0 1 -565 -1 0 1845
box 135 -1795 990 565
use dum_vert  dum_vert_18
timestamp 1730644682
transform 0 1 1795 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_19
timestamp 1730644682
transform 0 1 -565 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_20
timestamp 1730644682
transform 0 1 24250 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_21
timestamp 1730644682
transform 0 1 4290 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_22
timestamp 1730644682
transform 0 1 6785 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_23
timestamp 1730644682
transform 0 1 9280 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_24
timestamp 1730644682
transform 0 1 11775 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_25
timestamp 1730644682
transform 0 1 14270 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_26
timestamp 1730644682
transform 0 1 16765 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_27
timestamp 1730644682
transform 0 1 19260 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_28
timestamp 1730644682
transform 0 1 21755 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_29
timestamp 1730644682
transform 0 1 29240 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_30
timestamp 1730644682
transform 0 1 26745 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_31
timestamp 1730644682
transform 0 1 34230 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_32
timestamp 1730644682
transform 0 1 31735 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_33
timestamp 1730644682
transform 0 1 39220 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_34
timestamp 1730644682
transform 0 1 36725 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_35
timestamp 1730644682
transform 0 1 41580 -1 0 6975
box 135 -1795 990 565
use dum_vert  dum_vert_36
timestamp 1730644682
transform 0 1 41580 -1 0 135
box 135 -1795 990 565
use dum_vert  dum_vert_37
timestamp 1730644682
transform 0 1 41580 -1 0 990
box 135 -1795 990 565
use dum_vert  dum_vert_38
timestamp 1730644682
transform 0 1 41580 -1 0 1845
box 135 -1795 990 565
use dum_vert  dum_vert_39
timestamp 1730644682
transform 0 1 41580 -1 0 2700
box 135 -1795 990 565
use dum_vert  dum_vert_40
timestamp 1730644682
transform 0 1 41580 -1 0 3555
box 135 -1795 990 565
use dum_vert  dum_vert_41
timestamp 1730644682
transform 0 1 41580 -1 0 4410
box 135 -1795 990 565
use dum_vert  dum_vert_42
timestamp 1730644682
transform 0 1 41580 -1 0 5265
box 135 -1795 990 565
use dum_vert  dum_vert_43
timestamp 1730644682
transform 0 1 41580 -1 0 6120
box 135 -1795 990 565
use dum_vert  dum_vert_44
timestamp 1730644682
transform 0 1 41580 -1 0 14670
box 135 -1795 990 565
use dum_vert  dum_vert_45
timestamp 1730644682
transform 0 1 41580 -1 0 7830
box 135 -1795 990 565
use dum_vert  dum_vert_46
timestamp 1730644682
transform 0 1 41580 -1 0 8685
box 135 -1795 990 565
use dum_vert  dum_vert_47
timestamp 1730644682
transform 0 1 41580 -1 0 9540
box 135 -1795 990 565
use dum_vert  dum_vert_48
timestamp 1730644682
transform 0 1 41580 -1 0 10395
box 135 -1795 990 565
use dum_vert  dum_vert_49
timestamp 1730644682
transform 0 1 41580 -1 0 11250
box 135 -1795 990 565
use dum_vert  dum_vert_50
timestamp 1730644682
transform 0 1 41580 -1 0 12105
box 135 -1795 990 565
use dum_vert  dum_vert_51
timestamp 1730644682
transform 0 1 41580 -1 0 12960
box 135 -1795 990 565
use dum_vert  dum_vert_52
timestamp 1730644682
transform 0 1 41580 -1 0 13815
box 135 -1795 990 565
use end  end_0
timestamp 1729689530
transform 0 1 0 -1 0 13680
box 0 0 13680 2360
use end  end_1
timestamp 1729689530
transform 0 1 2495 -1 0 13680
box 0 0 13680 2360
use end  end_2
timestamp 1729689530
transform 0 1 34930 -1 0 13680
box 0 0 13680 2360
use end  end_3
timestamp 1729689530
transform 0 1 37425 -1 0 13680
box 0 0 13680 2360
use mid_2  mid_2_0
timestamp 1729709358
transform 1 0 17465 0 1 6840
box 0 -6840 4900 6840
use mid_2to4_  mid_2to4__0
timestamp 1729683266
transform 0 1 14970 -1 0 13680
box 0 0 13680 2360
use mid_2to4_  mid_2to4__1
timestamp 1729683266
transform 0 1 22455 -1 0 13680
box 0 0 13680 2360
use mid_4to8  mid_4to8_0
timestamp 1729685583
transform 0 1 9980 -1 0 13680
box 0 0 13680 2360
use mid_4to8  mid_4to8_1
timestamp 1729685583
transform 0 1 12475 -1 0 13680
box 0 0 13680 2360
use mid_4to8  mid_4to8_2
timestamp 1729685583
transform 0 1 24950 -1 0 13680
box 0 0 13680 2360
use mid_4to8  mid_4to8_3
timestamp 1729685583
transform 0 1 27445 -1 0 13680
box 0 0 13680 2360
use mid_6to8  mid_6to8_0
timestamp 1729688460
transform 0 1 4990 -1 0 13680
box 0 0 13680 2360
use mid_6to8  mid_6to8_1
timestamp 1729688460
transform 0 1 7485 -1 0 13680
box 0 0 13680 2360
use mid_6to8  mid_6to8_2
timestamp 1729688460
transform 0 1 29940 -1 0 13680
box 0 0 13680 2360
use mid_6to8  mid_6to8_3
timestamp 1729688460
transform 0 1 32435 -1 0 13680
box 0 0 13680 2360
use smpl_switch  smpl_switch_1
timestamp 1730647371
transform 1 0 -2990 0 -1 15105
box -400 -95 615 15115
<< labels >>
flabel metal3 -2486 15033 -2431 15058 0 FreeSans 80 0 0 0 vdd
port 18 nsew
flabel metal1 -2406 15031 -2360 15044 0 FreeSans 80 0 0 0 vin
port 60 nsew
flabel metal1 -2395 16296 -2349 16309 0 FreeSans 80 0 0 0 phi2_n7
port 98 nsew
flabel metal1 -2397 16226 -2351 16239 0 FreeSans 80 0 0 0 phi1_n7
port 96 nsew
flabel metal1 -2399 16155 -2353 16168 0 FreeSans 80 0 0 0 phi2_n6
port 94 nsew
flabel metal1 -2397 16085 -2351 16098 0 FreeSans 80 0 0 0 phi1_n6
port 92 nsew
flabel metal1 -2393 16016 -2347 16029 0 FreeSans 80 0 0 0 phi2_n5
port 90 nsew
flabel metal1 -2394 15946 -2348 15959 0 FreeSans 80 0 0 0 phi1_n5
port 88 nsew
flabel metal1 -2395 15876 -2349 15889 0 FreeSans 80 0 0 0 phi2_n4
port 86 nsew
flabel metal1 -2396 15806 -2350 15819 0 FreeSans 80 0 0 0 phi1_n4
port 84 nsew
flabel metal1 -2396 15736 -2350 15749 0 FreeSans 80 0 0 0 phi2_n3
port 82 nsew
flabel metal1 -2397 15666 -2351 15679 0 FreeSans 80 0 0 0 phi1_n3
port 80 nsew
flabel metal1 -2398 15596 -2352 15609 0 FreeSans 80 0 0 0 phi2_n2
port 78 nsew
flabel metal1 -2399 15525 -2353 15538 0 FreeSans 80 0 0 0 phi1_n2
port 76 nsew
flabel metal1 -2400 15456 -2354 15469 0 FreeSans 80 0 0 0 phi2_n1
port 74 nsew
flabel metal1 -2401 15385 -2355 15398 0 FreeSans 80 0 0 0 phi1_n1
port 72 nsew
flabel metal1 -2401 15316 -2355 15329 0 FreeSans 80 0 0 0 phi2_n0
port 70 nsew
flabel metal1 -2401 15245 -2355 15258 0 FreeSans 80 0 0 0 phi1_n0
port 68 nsew
flabel metal1 -2400 15175 -2354 15188 0 FreeSans 80 0 0 0 sphi2_n
port 66 nsew
flabel metal1 -2399 15107 -2353 15120 0 FreeSans 80 0 0 0 sphi1_n
port 64 nsew
flabel metal1 -2411 14960 -2365 14972 0 FreeSans 80 0 0 0 gnd
port 58 nsew
flabel metal3 -2473 16297 -2419 16322 0 FreeSans 80 0 0 0 phi27
port 56 nsew
flabel metal3 -2475 16227 -2421 16252 0 FreeSans 80 0 0 0 phi17
port 54 nsew
flabel metal3 -2477 16157 -2423 16182 0 FreeSans 80 0 0 0 phi26
port 52 nsew
flabel metal3 -2476 16086 -2422 16111 0 FreeSans 80 0 0 0 phi16
port 50 nsew
flabel metal3 -2475 16016 -2421 16041 0 FreeSans 80 0 0 0 phi25
port 48 nsew
flabel metal3 -2477 15948 -2423 15973 0 FreeSans 80 0 0 0 phi15
port 46 nsew
flabel metal3 -2477 15878 -2423 15903 0 FreeSans 80 0 0 0 phi24
port 44 nsew
flabel metal3 -2479 15809 -2425 15834 0 FreeSans 80 0 0 0 phi14
port 42 nsew
flabel metal3 -2478 15737 -2424 15762 0 FreeSans 80 0 0 0 phi23
port 40 nsew
flabel metal3 -2484 15668 -2430 15693 0 FreeSans 80 0 0 0 phi13
port 38 nsew
flabel metal3 -2490 15597 -2436 15622 0 FreeSans 80 0 0 0 phi22
port 36 nsew
flabel metal3 -2487 15527 -2433 15552 0 FreeSans 80 0 0 0 phi12
port 34 nsew
flabel metal3 -2485 15457 -2431 15482 0 FreeSans 80 0 0 0 phi21
port 32 nsew
flabel metal3 -2486 15388 -2432 15413 0 FreeSans 80 0 0 0 phi11
port 30 nsew
flabel metal3 -2487 15318 -2433 15343 0 FreeSans 80 0 0 0 phi20
port 28 nsew
flabel metal3 -2491 15246 -2437 15271 0 FreeSans 80 0 0 0 phi10
port 26 nsew
flabel metal3 -2488 15177 -2436 15204 0 FreeSans 80 0 0 0 sphi2
port 24 nsew
flabel metal3 -2485 15106 -2433 15133 0 FreeSans 80 0 0 0 sphi1
port 22 nsew
flabel metal3 -2487 14962 -2432 14987 0 FreeSans 80 0 0 0 sub
port 14 nsew
<< end >>
