magic
tech sky130A
magscale 1 2
timestamp 1729535358
<< pwell >>
rect 1140 -930 1160 -890
rect 1520 -950 1860 -880
<< locali >>
rect 710 180 1520 200
rect 710 140 840 180
rect 1080 140 1160 180
rect 1400 140 1520 180
rect 710 110 1520 140
rect 710 -890 1520 -860
rect 710 -930 840 -890
rect 1080 -930 1140 -890
rect 1400 -930 1520 -890
rect 710 -950 1520 -930
<< viali >>
rect 840 140 1080 180
rect 1160 140 1400 180
rect 840 -930 1080 -890
rect 1140 -930 1400 -890
<< metal1 >>
rect 390 890 1860 920
rect 390 830 1860 860
rect 390 720 1860 750
rect 390 660 1860 690
rect 390 550 1860 580
rect 390 490 1860 520
rect 390 380 1860 410
rect 390 320 810 350
rect 800 290 810 320
rect 870 320 1860 350
rect 870 290 880 320
rect 1330 260 1340 290
rect 390 230 1340 260
rect 1400 260 1410 290
rect 1400 230 1860 260
rect 390 180 1860 200
rect 390 140 840 180
rect 1080 140 1160 180
rect 1400 140 1860 180
rect 390 130 1860 140
rect 910 70 1010 80
rect 910 10 930 70
rect 990 10 1010 70
rect 910 0 1010 10
rect 1220 70 1320 80
rect 1220 10 1240 70
rect 1300 10 1320 70
rect 1220 0 1320 10
rect 900 -340 930 -220
rect 850 -350 930 -340
rect 850 -410 860 -350
rect 920 -410 930 -350
rect 850 -420 930 -410
rect 900 -540 930 -420
rect 990 -340 1020 -220
rect 1210 -340 1240 -220
rect 990 -350 1240 -340
rect 990 -410 1030 -350
rect 1090 -410 1140 -350
rect 1200 -410 1240 -350
rect 990 -420 1240 -410
rect 990 -540 1020 -420
rect 1210 -540 1240 -420
rect 1300 -340 1330 -220
rect 1300 -350 1380 -340
rect 1300 -410 1310 -350
rect 1370 -410 1380 -350
rect 1300 -420 1380 -410
rect 1300 -540 1330 -420
rect 910 -770 1010 -760
rect 910 -830 930 -770
rect 990 -830 1010 -770
rect 910 -840 1010 -830
rect 1220 -770 1320 -760
rect 1220 -830 1240 -770
rect 1300 -830 1320 -770
rect 1220 -840 1320 -830
rect 390 -890 1860 -880
rect 390 -930 840 -890
rect 1080 -930 1140 -890
rect 1400 -930 1860 -890
rect 390 -950 1860 -930
rect 390 -1010 1860 -980
rect 390 -1120 1860 -1090
rect 390 -1180 1860 -1150
rect 390 -1290 1860 -1260
rect 390 -1350 1860 -1320
rect 390 -1460 1860 -1430
rect 390 -1520 1860 -1490
<< via1 >>
rect 810 290 870 350
rect 1340 230 1400 290
rect 930 10 990 70
rect 1240 10 1300 70
rect 860 -410 920 -350
rect 1030 -410 1090 -350
rect 1140 -410 1200 -350
rect 1310 -410 1370 -350
rect 930 -830 990 -770
rect 1240 -830 1300 -770
<< metal2 >>
rect 800 290 810 350
rect 870 290 880 350
rect 850 -340 880 290
rect 950 80 980 370
rect 1260 80 1290 370
rect 1330 230 1340 290
rect 1400 230 1410 290
rect 920 70 1000 80
rect 920 10 930 70
rect 990 10 1000 70
rect 920 0 1000 10
rect 1230 70 1310 80
rect 1230 10 1240 70
rect 1300 10 1310 70
rect 1230 0 1310 10
rect 1350 -340 1380 230
rect 850 -350 930 -340
rect 850 -410 860 -350
rect 920 -410 930 -350
rect 850 -420 930 -410
rect 1020 -350 1210 -340
rect 1020 -410 1030 -350
rect 1090 -410 1140 -350
rect 1200 -410 1210 -350
rect 1020 -420 1210 -410
rect 1300 -350 1380 -340
rect 1300 -410 1310 -350
rect 1370 -410 1380 -350
rect 1300 -420 1380 -410
rect 920 -770 1000 -760
rect 920 -830 930 -770
rect 990 -830 1000 -770
rect 920 -840 1000 -830
rect 950 -970 980 -840
rect 1100 -1620 1130 -420
rect 1230 -770 1310 -760
rect 1230 -830 1240 -770
rect 1300 -830 1310 -770
rect 1230 -840 1310 -830
rect 1260 -970 1290 -840
rect 1070 -1630 1160 -1620
rect 1070 -1690 1080 -1630
rect 1150 -1690 1160 -1630
rect 1070 -1700 1160 -1690
<< via2 >>
rect 1080 -1690 1150 -1630
<< metal4 >>
rect 471 -3280 541 -3210
use sky130_fd_pr__cap_mim_m3_1_BZXSER  sky130_fd_pr__cap_mim_m3_1_BZXSER_0 /home/imasha
timestamp 1728835232
transform 0 1 1120 1 0 -2484
box -886 -740 886 740
use sky130_fd_pr__nfet_01v8_5WU4M2  sky130_fd_pr__nfet_01v8_5WU4M2_0 ~/final
timestamp 1728804544
transform -1 0 1271 0 -1 -661
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_QKK3FL  sky130_fd_pr__pfet_01v8_QKK3FL_0 ~/final
timestamp 1728804544
transform -1 0 1271 0 -1 -96
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_NKK3FE  XM1 ~/final
timestamp 1728804544
transform 1 0 961 0 1 -96
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_5WP7M2  XM2 ~/final
timestamp 1728804544
transform 1 0 961 0 1 -661
box -211 -279 211 279
<< labels >>
flabel metal1 770 -940 830 -880 0 FreeSans 256 0 0 0 sub
port 6 nsew
flabel metal1 1080 -940 1140 -880 0 FreeSans 256 0 0 0 sub
port 1 nsew
flabel metal1 770 130 830 190 0 FreeSans 256 0 0 0 Vdd
port 3 nsew
flabel metal1 1100 130 1150 190 0 FreeSans 256 0 0 0 Vdd
port 7 nsew
flabel metal1 862 -408 922 -348 0 FreeSans 256 0 0 0 Vin
port 5 nsew
flabel metal1 1312 -408 1372 -348 0 FreeSans 256 0 0 0 GND
port 9 nsew
flabel metal1 928 8 988 68 0 FreeSans 256 0 0 0 phi1_n
port 4 nsew
flabel metal1 1234 12 1294 72 0 FreeSans 256 0 0 0 phi2_n
port 10 nsew
flabel via1 930 -830 990 -770 0 FreeSans 256 0 0 0 phi1
port 2 nsew
flabel via1 1240 -830 1300 -770 0 FreeSans 256 0 0 0 phi2
port 8 nsew
flabel metal4 481 -3270 541 -3210 0 FreeSans 256 0 0 0 com_x
port 0 nsew
<< end >>
