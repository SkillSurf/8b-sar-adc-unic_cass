* SPICE3 file created from dac_top_final.ext - technology: sky130A

X0 dum_vert_52/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1 dum_vert_52/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2 dum_vert_52/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3 dum_vert_52/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4 gnd dum_vert_52/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X5 dum_vert_41/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=113.68 ps=1.01136k w=1 l=0.15
X6 dum_vert_41/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=113.68 ps=1.01136k w=1 l=0.15
X7 dum_vert_41/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8 dum_vert_41/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9 gnd dum_vert_41/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X10 dum_vert_30/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X11 dum_vert_30/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X12 dum_vert_30/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X13 dum_vert_30/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X14 gnd dum_vert_30/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X15 dum_vert_42/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X16 dum_vert_42/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X17 dum_vert_42/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X18 dum_vert_42/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X19 gnd dum_vert_42/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X20 dum_vert_31/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X21 dum_vert_31/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X22 dum_vert_31/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X23 dum_vert_31/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X24 gnd dum_vert_31/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X25 dum_vert_20/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X26 dum_vert_20/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X27 dum_vert_20/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X28 dum_vert_20/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X29 gnd dum_vert_20/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X30 dum_vert_43/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X31 dum_vert_43/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X32 dum_vert_43/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X33 dum_vert_43/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X34 gnd dum_vert_43/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X35 dum_vert_32/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X36 dum_vert_32/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X37 dum_vert_32/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X38 dum_vert_32/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X39 gnd dum_vert_32/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X40 dum_vert_21/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X41 dum_vert_21/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X42 dum_vert_21/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X43 dum_vert_21/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X44 gnd dum_vert_21/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X45 dum_vert_10/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X46 dum_vert_10/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X47 dum_vert_10/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X48 dum_vert_10/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X49 gnd dum_vert_10/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X50 dum_vert_0/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X51 dum_vert_0/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X52 dum_vert_0/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X53 dum_vert_0/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X54 gnd dum_vert_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X55 dum_vert_44/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X56 dum_vert_44/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X57 dum_vert_44/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X58 dum_vert_44/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X59 gnd dum_vert_44/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X60 dum_vert_33/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X61 dum_vert_33/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X62 dum_vert_33/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X63 dum_vert_33/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X64 gnd dum_vert_33/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X65 cap_dum_0/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X66 cap_dum_0/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X67 cap_dum_0/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X68 cap_dum_0/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X69 gnd cap_dum_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X70 dum_vert_22/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X71 dum_vert_22/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X72 dum_vert_22/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X73 dum_vert_22/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X74 gnd dum_vert_22/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X75 dum_vert_1/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X76 dum_vert_1/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X77 dum_vert_1/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X78 dum_vert_1/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X79 gnd dum_vert_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X80 dum_vert_11/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X81 dum_vert_11/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X82 dum_vert_11/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X83 dum_vert_11/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X84 gnd dum_vert_11/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X85 dum_vert_45/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X86 dum_vert_45/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X87 dum_vert_45/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X88 dum_vert_45/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X89 gnd dum_vert_45/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X90 dum_vert_34/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X91 dum_vert_34/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X92 dum_vert_34/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X93 dum_vert_34/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X94 gnd dum_vert_34/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X95 cap_dum_1/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X96 cap_dum_1/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X97 cap_dum_1/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X98 cap_dum_1/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X99 gnd cap_dum_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X100 dum_vert_23/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X101 dum_vert_23/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X102 dum_vert_23/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X103 dum_vert_23/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X104 gnd dum_vert_23/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X105 dum_vert_2/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X106 dum_vert_2/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X107 dum_vert_2/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X108 dum_vert_2/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X109 gnd dum_vert_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X110 dum_vert_12/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X111 dum_vert_12/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X112 dum_vert_12/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X113 dum_vert_12/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X114 gnd dum_vert_12/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X115 dum_vert_47/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X116 dum_vert_47/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X117 dum_vert_47/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X118 dum_vert_47/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X119 gnd dum_vert_47/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X120 dum_vert_46/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X121 dum_vert_46/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X122 dum_vert_46/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X123 dum_vert_46/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X124 gnd dum_vert_46/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X125 dum_vert_35/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X126 dum_vert_35/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X127 dum_vert_35/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X128 dum_vert_35/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X129 gnd dum_vert_35/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X130 dum_vert_36/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X131 dum_vert_36/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X132 dum_vert_36/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X133 dum_vert_36/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X134 gnd dum_vert_36/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X135 cap_dum_3/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X136 cap_dum_3/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X137 cap_dum_3/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X138 cap_dum_3/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X139 gnd cap_dum_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X140 cap_dum_2/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X141 cap_dum_2/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X142 cap_dum_2/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X143 cap_dum_2/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X144 gnd cap_dum_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X145 dum_vert_25/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X146 dum_vert_25/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X147 dum_vert_25/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X148 dum_vert_25/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X149 gnd dum_vert_25/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X150 dum_vert_24/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X151 dum_vert_24/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X152 dum_vert_24/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X153 dum_vert_24/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X154 gnd dum_vert_24/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X155 dum_vert_3/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X156 dum_vert_3/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X157 dum_vert_3/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X158 dum_vert_3/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X159 gnd dum_vert_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X160 dum_vert_14/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X161 dum_vert_14/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X162 dum_vert_14/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X163 dum_vert_14/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X164 gnd dum_vert_14/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X165 dum_vert_13/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X166 dum_vert_13/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X167 dum_vert_13/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X168 dum_vert_13/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X169 gnd dum_vert_13/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X170 dum_vert_48/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X171 dum_vert_48/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X172 dum_vert_48/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X173 dum_vert_48/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X174 gnd dum_vert_48/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X175 dum_vert_37/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X176 dum_vert_37/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X177 dum_vert_37/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X178 dum_vert_37/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X179 gnd dum_vert_37/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X180 cap_dum_4/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X181 cap_dum_4/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X182 cap_dum_4/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X183 cap_dum_4/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X184 gnd cap_dum_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X185 dum_vert_26/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X186 dum_vert_26/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X187 dum_vert_26/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X188 dum_vert_26/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X189 gnd dum_vert_26/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X190 dum_vert_4/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X191 dum_vert_4/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X192 dum_vert_4/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X193 dum_vert_4/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X194 gnd dum_vert_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X195 dum_vert_15/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X196 dum_vert_15/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X197 dum_vert_15/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X198 dum_vert_15/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X199 gnd dum_vert_15/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X200 dum_vert_49/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X201 dum_vert_49/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X202 dum_vert_49/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X203 dum_vert_49/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X204 gnd dum_vert_49/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X205 dum_vert_38/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X206 dum_vert_38/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X207 dum_vert_38/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X208 dum_vert_38/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X209 gnd dum_vert_38/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X210 cap_dum_5/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X211 cap_dum_5/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X212 cap_dum_5/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X213 cap_dum_5/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X214 gnd cap_dum_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X215 dum_vert_27/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X216 dum_vert_27/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X217 dum_vert_27/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X218 dum_vert_27/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X219 gnd dum_vert_27/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X220 dum_vert_5/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X221 dum_vert_5/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X222 dum_vert_5/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X223 dum_vert_5/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X224 gnd dum_vert_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X225 dum_vert_16/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X226 dum_vert_16/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X227 dum_vert_16/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X228 dum_vert_16/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X229 gnd dum_vert_16/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X230 dum_vert_39/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X231 dum_vert_39/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X232 dum_vert_39/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X233 dum_vert_39/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X234 gnd dum_vert_39/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X235 cap_dum_6/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X236 cap_dum_6/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X237 cap_dum_6/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X238 cap_dum_6/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X239 gnd cap_dum_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X240 dum_vert_28/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X241 dum_vert_28/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X242 dum_vert_28/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X243 dum_vert_28/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X244 gnd dum_vert_28/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X245 mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X246 mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X247 mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=80.04 ps=712.08 w=1 l=0.15
X248 mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=80.04 ps=712.08 w=1 l=0.15
X249 smpl_switch_1/smpl_switch_1/Vout mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X250 mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X251 mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X252 mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X253 mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X254 smpl_switch_1/smpl_switch_1/Vout mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X255 mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X256 mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X257 mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X258 mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X259 smpl_switch_1/smpl_switch_1/Vout mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X260 mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X261 mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X262 mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X263 mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X264 smpl_switch_1/smpl_switch_1/Vout mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X265 mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X266 mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X267 mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X268 mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X269 smpl_switch_1/smpl_switch_1/Vout mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X270 mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X271 mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n4 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X272 mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n4 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X273 mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi14 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X274 smpl_switch_1/smpl_switch_1/Vout mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X275 mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X276 mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X277 mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X278 mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X279 smpl_switch_1/smpl_switch_1/Vout mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X280 mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X281 mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X282 mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X283 mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X284 smpl_switch_1/smpl_switch_1/Vout mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X285 mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X286 mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X287 mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X288 mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X289 smpl_switch_1/smpl_switch_1/Vout mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X290 mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X291 mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X292 mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X293 mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X294 smpl_switch_1/smpl_switch_1/Vout mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X295 mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X296 mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X297 mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X298 mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X299 smpl_switch_1/smpl_switch_1/Vout mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X300 mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X301 mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X302 mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X303 mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X304 smpl_switch_1/smpl_switch_1/Vout mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X305 mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X306 mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n4 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X307 mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n4 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X308 mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi14 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X309 smpl_switch_1/smpl_switch_1/Vout mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X310 mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X311 mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X312 mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X313 mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X314 smpl_switch_1/smpl_switch_1/Vout mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X315 mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X316 mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X317 mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X318 mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X319 smpl_switch_1/smpl_switch_1/Vout mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X320 mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X321 mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X322 mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X323 mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X324 smpl_switch_1/smpl_switch_1/Vout mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X325 dum_vert_6/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X326 dum_vert_6/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X327 dum_vert_6/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X328 dum_vert_6/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X329 gnd dum_vert_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X330 dum_vert_17/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X331 dum_vert_17/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X332 dum_vert_17/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X333 dum_vert_17/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X334 gnd dum_vert_17/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X335 cap_dum_7/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X336 cap_dum_7/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X337 cap_dum_7/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X338 cap_dum_7/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X339 gnd cap_dum_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X340 dum_vert_29/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X341 dum_vert_29/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X342 dum_vert_29/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X343 dum_vert_29/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X344 gnd dum_vert_29/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X345 mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X346 mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X347 mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X348 mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X349 smpl_switch_1/smpl_switch_1/Vout mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X350 mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X351 mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X352 mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X353 mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X354 smpl_switch_1/smpl_switch_1/Vout mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X355 mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X356 mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X357 mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X358 mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X359 smpl_switch_1/smpl_switch_1/Vout mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X360 mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X361 mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X362 mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X363 mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X364 smpl_switch_1/smpl_switch_1/Vout mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X365 mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X366 mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X367 mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X368 mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X369 smpl_switch_1/smpl_switch_1/Vout mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X370 mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X371 mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n4 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X372 mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n4 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X373 mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi14 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X374 smpl_switch_1/smpl_switch_1/Vout mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X375 mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X376 mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X377 mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X378 mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X379 smpl_switch_1/smpl_switch_1/Vout mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X380 mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X381 mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X382 mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X383 mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X384 smpl_switch_1/smpl_switch_1/Vout mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X385 mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X386 mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X387 mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X388 mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X389 smpl_switch_1/smpl_switch_1/Vout mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X390 mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X391 mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X392 mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X393 mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X394 smpl_switch_1/smpl_switch_1/Vout mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X395 mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X396 mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X397 mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X398 mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X399 smpl_switch_1/smpl_switch_1/Vout mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X400 mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X401 mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X402 mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X403 mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X404 smpl_switch_1/smpl_switch_1/Vout mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X405 mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X406 mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n4 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X407 mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n4 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X408 mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi14 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X409 smpl_switch_1/smpl_switch_1/Vout mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X410 mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X411 mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X412 mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X413 mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X414 smpl_switch_1/smpl_switch_1/Vout mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X415 mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X416 mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X417 mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X418 mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X419 smpl_switch_1/smpl_switch_1/Vout mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X420 mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X421 mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X422 mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X423 mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X424 smpl_switch_1/smpl_switch_1/Vout mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X425 dum_vert_18/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X426 dum_vert_18/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X427 dum_vert_18/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X428 dum_vert_18/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X429 gnd dum_vert_18/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X430 dum_vert_7/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X431 dum_vert_7/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X432 dum_vert_7/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X433 dum_vert_7/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X434 gnd dum_vert_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X435 cap_dum_8/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X436 cap_dum_8/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X437 cap_dum_8/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X438 cap_dum_8/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X439 gnd cap_dum_8/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X440 mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X441 mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X442 mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X443 mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X444 smpl_switch_1/smpl_switch_1/Vout mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X445 mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X446 mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X447 mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X448 mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X449 smpl_switch_1/smpl_switch_1/Vout mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X450 mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X451 mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X452 mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X453 mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X454 smpl_switch_1/smpl_switch_1/Vout mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X455 mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X456 mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X457 mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X458 mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X459 smpl_switch_1/smpl_switch_1/Vout mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X460 mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X461 mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X462 mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X463 mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X464 smpl_switch_1/smpl_switch_1/Vout mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X465 mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X466 mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n4 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X467 mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n4 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X468 mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi14 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X469 smpl_switch_1/smpl_switch_1/Vout mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X470 mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X471 mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X472 mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X473 mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X474 smpl_switch_1/smpl_switch_1/Vout mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X475 mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X476 mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X477 mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X478 mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X479 smpl_switch_1/smpl_switch_1/Vout mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X480 mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X481 mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X482 mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X483 mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X484 smpl_switch_1/smpl_switch_1/Vout mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X485 mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X486 mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X487 mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X488 mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X489 smpl_switch_1/smpl_switch_1/Vout mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X490 mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X491 mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X492 mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X493 mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X494 smpl_switch_1/smpl_switch_1/Vout mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X495 mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X496 mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X497 mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X498 mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X499 smpl_switch_1/smpl_switch_1/Vout mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X500 mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X501 mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n4 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X502 mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n4 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X503 mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi14 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X504 smpl_switch_1/smpl_switch_1/Vout mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X505 mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X506 mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X507 mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X508 mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X509 smpl_switch_1/smpl_switch_1/Vout mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X510 mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X511 mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X512 mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X513 mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X514 smpl_switch_1/smpl_switch_1/Vout mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X515 mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X516 mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X517 mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X518 mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X519 smpl_switch_1/smpl_switch_1/Vout mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X520 mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X521 mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X522 mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X523 mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X524 smpl_switch_1/smpl_switch_1/Vout mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X525 mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X526 mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X527 mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X528 mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X529 smpl_switch_1/smpl_switch_1/Vout mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X530 mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X531 mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X532 mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X533 mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X534 smpl_switch_1/smpl_switch_1/Vout mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X535 mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X536 mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X537 mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X538 mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X539 smpl_switch_1/smpl_switch_1/Vout mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X540 mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X541 mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X542 mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X543 mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X544 smpl_switch_1/smpl_switch_1/Vout mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X545 mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X546 mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n4 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X547 mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n4 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X548 mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi14 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X549 smpl_switch_1/smpl_switch_1/Vout mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X550 mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X551 mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X552 mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X553 mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X554 smpl_switch_1/smpl_switch_1/Vout mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X555 mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X556 mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X557 mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X558 mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X559 smpl_switch_1/smpl_switch_1/Vout mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X560 mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X561 mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X562 mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X563 mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X564 smpl_switch_1/smpl_switch_1/Vout mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X565 mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X566 mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X567 mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X568 mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X569 smpl_switch_1/smpl_switch_1/Vout mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X570 mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X571 mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X572 mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X573 mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X574 smpl_switch_1/smpl_switch_1/Vout mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X575 mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X576 mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X577 mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X578 mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X579 smpl_switch_1/smpl_switch_1/Vout mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X580 mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X581 mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n4 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X582 mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n4 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X583 mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi14 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X584 smpl_switch_1/smpl_switch_1/Vout mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X585 mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X586 mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X587 mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X588 mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X589 smpl_switch_1/smpl_switch_1/Vout mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X590 mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X591 mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X592 mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X593 mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X594 smpl_switch_1/smpl_switch_1/Vout mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X595 mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X596 mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X597 mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X598 mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X599 smpl_switch_1/smpl_switch_1/Vout mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X600 dum_vert_9/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X601 dum_vert_9/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X602 dum_vert_9/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X603 dum_vert_9/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X604 gnd dum_vert_9/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X605 dum_vert_8/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X606 dum_vert_8/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X607 dum_vert_8/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X608 dum_vert_8/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X609 gnd dum_vert_8/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X610 dum_vert_19/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X611 dum_vert_19/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X612 dum_vert_19/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X613 dum_vert_19/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X614 gnd dum_vert_19/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X615 mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X616 mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X617 mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X618 mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X619 smpl_switch_1/smpl_switch_1/Vout mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X620 mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi23 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X621 mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n3 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X622 mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n3 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X623 mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi13 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X624 smpl_switch_1/smpl_switch_1/Vout mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X625 mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X626 mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X627 mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X628 mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X629 smpl_switch_1/smpl_switch_1/Vout mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X630 mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X631 mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X632 mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X633 mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X634 smpl_switch_1/smpl_switch_1/Vout mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X635 mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X636 mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X637 mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X638 mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X639 smpl_switch_1/smpl_switch_1/Vout mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X640 mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X641 mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X642 mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X643 mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X644 smpl_switch_1/smpl_switch_1/Vout mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X645 mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X646 mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n4 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X647 mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n4 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X648 mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi14 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X649 smpl_switch_1/smpl_switch_1/Vout mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X650 mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi22 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X651 mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n2 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X652 mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n2 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X653 mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi12 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X654 smpl_switch_1/smpl_switch_1/Vout mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X655 mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi23 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X656 mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n3 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X657 mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n3 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X658 mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi13 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X659 smpl_switch_1/smpl_switch_1/Vout mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X660 mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X661 mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X662 mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X663 mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X664 smpl_switch_1/smpl_switch_1/Vout mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X665 mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi22 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X666 mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n2 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X667 mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n2 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X668 mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi12 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X669 smpl_switch_1/smpl_switch_1/Vout mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X670 mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X671 mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n4 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X672 mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n4 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X673 mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi14 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X674 smpl_switch_1/smpl_switch_1/Vout mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X675 mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X676 mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X677 mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X678 mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X679 smpl_switch_1/smpl_switch_1/Vout mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X680 mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X681 mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X682 mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X683 mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X684 smpl_switch_1/smpl_switch_1/Vout mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X685 mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X686 mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X687 mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X688 mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X689 smpl_switch_1/smpl_switch_1/Vout mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X690 mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X691 mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X692 mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X693 mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X694 smpl_switch_1/smpl_switch_1/Vout mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X695 mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X696 mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X697 mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X698 mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X699 smpl_switch_1/smpl_switch_1/Vout mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X700 mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi23 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X701 mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n3 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X702 mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n3 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X703 mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi13 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X704 smpl_switch_1/smpl_switch_1/Vout mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X705 mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X706 mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X707 mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X708 mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X709 smpl_switch_1/smpl_switch_1/Vout mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X710 mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X711 mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X712 mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X713 mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X714 smpl_switch_1/smpl_switch_1/Vout mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X715 mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X716 mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X717 mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X718 mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X719 smpl_switch_1/smpl_switch_1/Vout mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X720 mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X721 mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X722 mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X723 mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X724 smpl_switch_1/smpl_switch_1/Vout mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X725 mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X726 mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n4 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X727 mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n4 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X728 mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi14 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X729 smpl_switch_1/smpl_switch_1/Vout mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X730 mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi22 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X731 mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n2 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X732 mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n2 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X733 mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi12 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X734 smpl_switch_1/smpl_switch_1/Vout mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X735 mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi23 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X736 mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n3 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X737 mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n3 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X738 mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi13 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X739 smpl_switch_1/smpl_switch_1/Vout mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X740 mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X741 mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X742 mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X743 mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X744 smpl_switch_1/smpl_switch_1/Vout mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X745 mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi22 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X746 mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n2 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X747 mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n2 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X748 mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi12 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X749 smpl_switch_1/smpl_switch_1/Vout mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X750 mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X751 mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n4 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X752 mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n4 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X753 mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi14 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X754 smpl_switch_1/smpl_switch_1/Vout mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X755 mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X756 mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X757 mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X758 mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X759 smpl_switch_1/smpl_switch_1/Vout mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X760 mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X761 mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X762 mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X763 mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X764 smpl_switch_1/smpl_switch_1/Vout mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X765 mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X766 mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X767 mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X768 mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X769 smpl_switch_1/smpl_switch_1/Vout mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X770 mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X771 mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X772 mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X773 mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X774 smpl_switch_1/smpl_switch_1/Vout mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X775 mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X776 mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X777 mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X778 mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X779 smpl_switch_1/smpl_switch_1/Vout mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X780 mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X781 mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X782 mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X783 mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X784 smpl_switch_1/smpl_switch_1/Vout mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X785 mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X786 mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X787 mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X788 mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X789 smpl_switch_1/smpl_switch_1/Vout mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X790 mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X791 mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X792 mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X793 mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X794 smpl_switch_1/smpl_switch_1/Vout mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X795 mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X796 mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X797 mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X798 mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X799 smpl_switch_1/smpl_switch_1/Vout mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X800 mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X801 mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X802 mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X803 mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X804 smpl_switch_1/smpl_switch_1/Vout mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X805 mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X806 mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X807 mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X808 mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X809 smpl_switch_1/smpl_switch_1/Vout mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X810 mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X811 mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X812 mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X813 mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X814 smpl_switch_1/smpl_switch_1/Vout mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X815 mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X816 mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X817 mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X818 mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X819 smpl_switch_1/smpl_switch_1/Vout mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X820 mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X821 mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X822 mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X823 mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X824 smpl_switch_1/smpl_switch_1/Vout mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X825 mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X826 mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X827 mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X828 mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X829 smpl_switch_1/smpl_switch_1/Vout mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X830 mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X831 mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X832 mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X833 mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X834 smpl_switch_1/smpl_switch_1/Vout mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X835 mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X836 mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X837 mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X838 mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X839 smpl_switch_1/smpl_switch_1/Vout mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X840 mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X841 mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X842 mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X843 mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X844 smpl_switch_1/smpl_switch_1/Vout mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X845 mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X846 mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X847 mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X848 mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X849 smpl_switch_1/smpl_switch_1/Vout mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X850 mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X851 mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X852 mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X853 mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X854 smpl_switch_1/smpl_switch_1/Vout mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X855 end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X856 end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X857 end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X858 end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X859 smpl_switch_1/smpl_switch_1/Vout end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X860 end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X861 end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X862 end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X863 end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X864 smpl_switch_1/smpl_switch_1/Vout end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X865 end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X866 end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X867 end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X868 end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X869 smpl_switch_1/smpl_switch_1/Vout end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X870 end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X871 end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X872 end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X873 end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X874 smpl_switch_1/smpl_switch_1/Vout end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X875 end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X876 end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X877 end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X878 end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X879 smpl_switch_1/smpl_switch_1/Vout end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X880 end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X881 end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X882 end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X883 end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X884 smpl_switch_1/smpl_switch_1/Vout end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X885 end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X886 end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X887 end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X888 end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X889 smpl_switch_1/smpl_switch_1/Vout end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X890 end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X891 end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X892 end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X893 end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X894 smpl_switch_1/smpl_switch_1/Vout end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X895 end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X896 end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X897 end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X898 end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X899 smpl_switch_1/smpl_switch_1/Vout end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X900 end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X901 end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X902 end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X903 end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X904 smpl_switch_1/smpl_switch_1/Vout end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X905 end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X906 end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X907 end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X908 end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X909 smpl_switch_1/smpl_switch_1/Vout end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X910 end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X911 end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X912 end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X913 end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X914 smpl_switch_1/smpl_switch_1/Vout end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X915 end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X916 end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X917 end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X918 end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X919 smpl_switch_1/smpl_switch_1/Vout end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X920 end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X921 end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X922 end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X923 end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X924 smpl_switch_1/smpl_switch_1/Vout end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X925 end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X926 end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X927 end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X928 end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X929 smpl_switch_1/smpl_switch_1/Vout end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X930 end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X931 end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X932 end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X933 end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X934 smpl_switch_1/smpl_switch_1/Vout end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X935 mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X936 mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X937 mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X938 mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X939 smpl_switch_1/smpl_switch_1/Vout mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X940 mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X941 mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X942 mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X943 mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X944 smpl_switch_1/smpl_switch_1/Vout mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X945 mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X946 mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X947 mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X948 mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X949 smpl_switch_1/smpl_switch_1/Vout mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X950 mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X951 mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X952 mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X953 mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X954 smpl_switch_1/smpl_switch_1/Vout mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X955 mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X956 mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X957 mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X958 mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X959 smpl_switch_1/smpl_switch_1/Vout mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X960 mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X961 mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X962 mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X963 mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X964 smpl_switch_1/smpl_switch_1/Vout mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X965 mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X966 mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X967 mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X968 mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X969 smpl_switch_1/smpl_switch_1/Vout mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X970 mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X971 mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X972 mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X973 mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X974 smpl_switch_1/smpl_switch_1/Vout mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X975 mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X976 mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X977 mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X978 mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X979 smpl_switch_1/smpl_switch_1/Vout mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X980 mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X981 mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X982 mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X983 mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X984 smpl_switch_1/smpl_switch_1/Vout mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X985 mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X986 mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X987 mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X988 mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X989 smpl_switch_1/smpl_switch_1/Vout mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X990 mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X991 mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X992 mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X993 mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X994 smpl_switch_1/smpl_switch_1/Vout mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X995 mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X996 mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X997 mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X998 mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X999 smpl_switch_1/smpl_switch_1/Vout mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1000 mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1001 mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1002 mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1003 mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1004 smpl_switch_1/smpl_switch_1/Vout mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1005 mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1006 mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1007 mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1008 mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1009 smpl_switch_1/smpl_switch_1/Vout mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1010 mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1011 mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1012 mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1013 mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1014 smpl_switch_1/smpl_switch_1/Vout mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1015 end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1016 end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1017 end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1018 end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1019 smpl_switch_1/smpl_switch_1/Vout end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1020 end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1021 end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1022 end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1023 end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1024 smpl_switch_1/smpl_switch_1/Vout end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1025 end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1026 end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1027 end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1028 end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1029 smpl_switch_1/smpl_switch_1/Vout end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1030 end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1031 end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1032 end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1033 end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1034 smpl_switch_1/smpl_switch_1/Vout end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1035 end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1036 end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1037 end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1038 end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1039 smpl_switch_1/smpl_switch_1/Vout end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1040 end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1041 end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1042 end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1043 end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1044 smpl_switch_1/smpl_switch_1/Vout end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1045 end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1046 end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1047 end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1048 end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1049 smpl_switch_1/smpl_switch_1/Vout end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1050 end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1051 end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1052 end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1053 end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1054 smpl_switch_1/smpl_switch_1/Vout end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1055 end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1056 end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1057 end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1058 end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1059 smpl_switch_1/smpl_switch_1/Vout end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1060 end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1061 end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1062 end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1063 end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1064 smpl_switch_1/smpl_switch_1/Vout end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1065 end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1066 end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1067 end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1068 end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1069 smpl_switch_1/smpl_switch_1/Vout end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1070 end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1071 end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1072 end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1073 end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1074 smpl_switch_1/smpl_switch_1/Vout end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1075 end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1076 end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1077 end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1078 end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1079 smpl_switch_1/smpl_switch_1/Vout end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1080 end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1081 end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1082 end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1083 end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1084 smpl_switch_1/smpl_switch_1/Vout end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1085 end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1086 end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1087 end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1088 end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1089 smpl_switch_1/smpl_switch_1/Vout end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1090 end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1091 end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1092 end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1093 end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1094 smpl_switch_1/smpl_switch_1/Vout end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1095 end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1096 end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1097 end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1098 end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1099 smpl_switch_1/smpl_switch_1/Vout end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1100 end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1101 end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1102 end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1103 end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1104 smpl_switch_1/smpl_switch_1/Vout end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1105 end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1106 end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1107 end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1108 end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1109 smpl_switch_1/smpl_switch_1/Vout end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1110 end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1111 end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1112 end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1113 end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1114 smpl_switch_1/smpl_switch_1/Vout end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1115 end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1116 end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1117 end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1118 end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1119 smpl_switch_1/smpl_switch_1/Vout end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1120 end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1121 end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1122 end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1123 end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1124 smpl_switch_1/smpl_switch_1/Vout end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1125 end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1126 end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1127 end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1128 end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1129 smpl_switch_1/smpl_switch_1/Vout end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1130 end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1131 end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1132 end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1133 end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1134 smpl_switch_1/smpl_switch_1/Vout end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1135 end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1136 end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1137 end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1138 end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1139 smpl_switch_1/smpl_switch_1/Vout end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1140 end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1141 end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1142 end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1143 end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1144 smpl_switch_1/smpl_switch_1/Vout end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1145 end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1146 end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1147 end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1148 end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1149 smpl_switch_1/smpl_switch_1/Vout end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1150 end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1151 end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1152 end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1153 end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1154 smpl_switch_1/smpl_switch_1/Vout end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1155 end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1156 end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1157 end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1158 end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1159 smpl_switch_1/smpl_switch_1/Vout end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1160 end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1161 end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1162 end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1163 end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1164 smpl_switch_1/smpl_switch_1/Vout end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1165 end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1166 end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1167 end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1168 end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1169 smpl_switch_1/smpl_switch_1/Vout end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1170 end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1171 end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1172 end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1173 end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1174 smpl_switch_1/smpl_switch_1/Vout end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1175 mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1176 mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1177 mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1178 mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1179 smpl_switch_1/smpl_switch_1/Vout mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1180 mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1181 mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1182 mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1183 mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1184 smpl_switch_1/smpl_switch_1/Vout mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1185 mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1186 mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1187 mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1188 mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1189 smpl_switch_1/smpl_switch_1/Vout mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1190 mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1191 mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1192 mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1193 mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1194 smpl_switch_1/smpl_switch_1/Vout mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1195 mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1196 mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1197 mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1198 mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1199 smpl_switch_1/smpl_switch_1/Vout mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1200 mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1201 mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1202 mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1203 mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1204 smpl_switch_1/smpl_switch_1/Vout mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1205 mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1206 mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1207 mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1208 mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1209 smpl_switch_1/smpl_switch_1/Vout mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1210 mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1211 mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1212 mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1213 mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1214 smpl_switch_1/smpl_switch_1/Vout mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1215 mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1216 mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1217 mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1218 mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1219 smpl_switch_1/smpl_switch_1/Vout mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1220 mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1221 mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1222 mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1223 mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1224 smpl_switch_1/smpl_switch_1/Vout mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1225 mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1226 mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1227 mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1228 mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1229 smpl_switch_1/smpl_switch_1/Vout mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1230 mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1231 mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1232 mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1233 mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1234 smpl_switch_1/smpl_switch_1/Vout mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1235 mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1236 mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1237 mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1238 mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1239 smpl_switch_1/smpl_switch_1/Vout mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1240 mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1241 mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1242 mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1243 mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1244 smpl_switch_1/smpl_switch_1/Vout mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1245 mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1246 mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1247 mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1248 mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1249 smpl_switch_1/smpl_switch_1/Vout mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1250 mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1251 mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1252 mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1253 mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1254 smpl_switch_1/smpl_switch_1/Vout mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1255 cap_dum_10/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1256 cap_dum_10/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1257 cap_dum_10/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1258 cap_dum_10/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1259 gnd cap_dum_10/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1260 smpl_switch_1/smpl_switch_2/Vout sphi2_n smpl_switch_1/smpl_switch_0/Vin vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1261 smpl_switch_1/smpl_switch_2/Vout sphi2_n smpl_switch_1/smpl_switch_0/Vin vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1262 smpl_switch_1/smpl_switch_2/Vout sphi2 smpl_switch_1/smpl_switch_0/Vin sub sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1263 smpl_switch_1/smpl_switch_2/Vout sphi2 smpl_switch_1/smpl_switch_0/Vin sub sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1264 smpl_switch_1/smpl_switch_2/Vout sphi2_n smpl_switch_1/smpl_switch_0/Vin vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1265 smpl_switch_1/smpl_switch_2/Vout sphi2_n smpl_switch_1/smpl_switch_0/Vin vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1266 smpl_switch_1/smpl_switch_2/Vout sphi2 smpl_switch_1/smpl_switch_0/Vin sub sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1267 smpl_switch_1/smpl_switch_2/Vout sphi2 smpl_switch_1/smpl_switch_0/Vin sub sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1268 smpl_switch_1/smpl_switch_2/Vout sphi2_n smpl_switch_1/smpl_switch_0/Vin vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1269 smpl_switch_1/smpl_switch_2/Vout sphi2_n smpl_switch_1/smpl_switch_0/Vin vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1270 smpl_switch_1/smpl_switch_2/Vout sphi2 smpl_switch_1/smpl_switch_0/Vin sub sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1271 smpl_switch_1/smpl_switch_2/Vout sphi2_n smpl_switch_1/smpl_switch_0/Vin vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1272 smpl_switch_1/smpl_switch_2/Vout sphi2 smpl_switch_1/smpl_switch_0/Vin sub sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1273 smpl_switch_1/smpl_switch_2/Vout sphi2 smpl_switch_1/smpl_switch_0/Vin sub sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1274 smpl_switch_1/smpl_switch_2/Vout sphi2_n smpl_switch_1/smpl_switch_0/Vin vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1275 smpl_switch_1/smpl_switch_2/Vout sphi2_n smpl_switch_1/smpl_switch_0/Vin vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1276 smpl_switch_1/smpl_switch_2/Vout sphi2 smpl_switch_1/smpl_switch_0/Vin sub sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1277 smpl_switch_1/smpl_switch_2/Vout sphi2 smpl_switch_1/smpl_switch_0/Vin sub sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1278 smpl_switch_1/smpl_switch_2/Vout sphi2_n smpl_switch_1/smpl_switch_0/Vin vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1279 smpl_switch_1/smpl_switch_2/Vout sphi2 smpl_switch_1/smpl_switch_0/Vin sub sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1280 smpl_switch_1/smpl_switch_1/Vout sample_n smpl_switch_1/vcm vdd sky130_fd_pr__pfet_01v8 ad=2.9 pd=25.8 as=2.9 ps=25.8 w=1 l=0.15
X1281 smpl_switch_1/smpl_switch_1/Vout sample_n smpl_switch_1/vcm vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1282 smpl_switch_1/smpl_switch_1/Vout sample smpl_switch_1/vcm sub sky130_fd_pr__nfet_01v8 ad=2.9 pd=25.8 as=2.9 ps=25.8 w=1 l=0.15
X1283 smpl_switch_1/smpl_switch_1/Vout sample smpl_switch_1/vcm sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1284 smpl_switch_1/smpl_switch_1/Vout sample_n smpl_switch_1/vcm vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1285 smpl_switch_1/smpl_switch_1/Vout sample_n smpl_switch_1/vcm vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1286 smpl_switch_1/smpl_switch_1/Vout sample smpl_switch_1/vcm sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1287 smpl_switch_1/smpl_switch_1/Vout sample smpl_switch_1/vcm sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1288 smpl_switch_1/smpl_switch_1/Vout sample_n smpl_switch_1/vcm vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1289 smpl_switch_1/smpl_switch_1/Vout sample_n smpl_switch_1/vcm vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1290 smpl_switch_1/smpl_switch_1/Vout sample smpl_switch_1/vcm sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1291 smpl_switch_1/smpl_switch_1/Vout sample_n smpl_switch_1/vcm vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1292 smpl_switch_1/smpl_switch_1/Vout sample smpl_switch_1/vcm sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1293 smpl_switch_1/smpl_switch_1/Vout sample smpl_switch_1/vcm sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1294 smpl_switch_1/smpl_switch_1/Vout sample_n smpl_switch_1/vcm vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1295 smpl_switch_1/smpl_switch_1/Vout sample_n smpl_switch_1/vcm vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1296 smpl_switch_1/smpl_switch_1/Vout sample smpl_switch_1/vcm sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1297 smpl_switch_1/smpl_switch_1/Vout sample smpl_switch_1/vcm sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1298 smpl_switch_1/smpl_switch_1/Vout sample_n smpl_switch_1/vcm vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1299 smpl_switch_1/smpl_switch_1/Vout sample smpl_switch_1/vcm sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1300 smpl_switch_1/smpl_switch_2/Vout sphi1_n smpl_switch_1/vref vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=2.9 ps=25.8 w=1 l=0.15
X1301 smpl_switch_1/smpl_switch_2/Vout sphi1_n smpl_switch_1/vref vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1302 smpl_switch_1/smpl_switch_2/Vout sphi1 smpl_switch_1/vref sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=2.9 ps=25.8 w=1 l=0.15
X1303 smpl_switch_1/smpl_switch_2/Vout sphi1 smpl_switch_1/vref sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1304 smpl_switch_1/smpl_switch_2/Vout sphi1_n smpl_switch_1/vref vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1305 smpl_switch_1/smpl_switch_2/Vout sphi1_n smpl_switch_1/vref vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1306 smpl_switch_1/smpl_switch_2/Vout sphi1 smpl_switch_1/vref sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1307 smpl_switch_1/smpl_switch_2/Vout sphi1 smpl_switch_1/vref sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1308 smpl_switch_1/smpl_switch_2/Vout sphi1_n smpl_switch_1/vref vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1309 smpl_switch_1/smpl_switch_2/Vout sphi1_n smpl_switch_1/vref vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1310 smpl_switch_1/smpl_switch_2/Vout sphi1 smpl_switch_1/vref sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1311 smpl_switch_1/smpl_switch_2/Vout sphi1_n smpl_switch_1/vref vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1312 smpl_switch_1/smpl_switch_2/Vout sphi1 smpl_switch_1/vref sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1313 smpl_switch_1/smpl_switch_2/Vout sphi1 smpl_switch_1/vref sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1314 smpl_switch_1/smpl_switch_2/Vout sphi1_n smpl_switch_1/vref vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1315 smpl_switch_1/smpl_switch_2/Vout sphi1_n smpl_switch_1/vref vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1316 smpl_switch_1/smpl_switch_2/Vout sphi1 smpl_switch_1/vref sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1317 smpl_switch_1/smpl_switch_2/Vout sphi1 smpl_switch_1/vref sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1318 smpl_switch_1/smpl_switch_2/Vout sphi1_n smpl_switch_1/vref vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1319 smpl_switch_1/smpl_switch_2/Vout sphi1 smpl_switch_1/vref sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1320 end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1321 end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1322 end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1323 end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1324 smpl_switch_1/smpl_switch_1/Vout end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1325 end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1326 end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1327 end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1328 end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1329 smpl_switch_1/smpl_switch_1/Vout end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1330 end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1331 end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1332 end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1333 end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1334 smpl_switch_1/smpl_switch_1/Vout end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1335 end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1336 end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1337 end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1338 end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1339 smpl_switch_1/smpl_switch_1/Vout end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1340 end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1341 end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1342 end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1343 end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1344 smpl_switch_1/smpl_switch_1/Vout end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1345 end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1346 end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1347 end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1348 end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1349 smpl_switch_1/smpl_switch_1/Vout end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1350 end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1351 end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1352 end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1353 end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1354 smpl_switch_1/smpl_switch_1/Vout end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1355 end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1356 end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1357 end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1358 end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1359 smpl_switch_1/smpl_switch_1/Vout end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1360 end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1361 end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1362 end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1363 end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1364 smpl_switch_1/smpl_switch_1/Vout end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1365 end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1366 end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1367 end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1368 end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1369 smpl_switch_1/smpl_switch_1/Vout end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1370 end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1371 end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1372 end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1373 end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1374 smpl_switch_1/smpl_switch_1/Vout end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1375 end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1376 end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1377 end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1378 end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1379 smpl_switch_1/smpl_switch_1/Vout end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1380 end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1381 end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1382 end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1383 end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1384 smpl_switch_1/smpl_switch_1/Vout end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1385 end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1386 end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1387 end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1388 end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1389 smpl_switch_1/smpl_switch_1/Vout end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1390 end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1391 end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1392 end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1393 end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1394 smpl_switch_1/smpl_switch_1/Vout end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1395 end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1396 end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1397 end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1398 end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1399 smpl_switch_1/smpl_switch_1/Vout end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1400 mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1401 mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1402 mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1403 mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1404 smpl_switch_1/smpl_switch_1/Vout mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1405 mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1406 mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1407 mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1408 mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1409 smpl_switch_1/smpl_switch_1/Vout mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1410 mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1411 mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1412 mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1413 mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1414 smpl_switch_1/smpl_switch_1/Vout mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1415 mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1416 mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1417 mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1418 mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1419 smpl_switch_1/smpl_switch_1/Vout mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1420 mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1421 mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1422 mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1423 mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1424 smpl_switch_1/smpl_switch_1/Vout mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1425 mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1426 mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1427 mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1428 mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1429 smpl_switch_1/smpl_switch_1/Vout mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1430 mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1431 mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1432 mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1433 mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1434 smpl_switch_1/smpl_switch_1/Vout mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1435 mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1436 mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1437 mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1438 mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1439 smpl_switch_1/smpl_switch_1/Vout mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1440 mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1441 mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1442 mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1443 mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1444 smpl_switch_1/smpl_switch_1/Vout mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1445 mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1446 mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1447 mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1448 mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1449 smpl_switch_1/smpl_switch_1/Vout mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1450 mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1451 mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1452 mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1453 mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1454 smpl_switch_1/smpl_switch_1/Vout mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1455 mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1456 mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1457 mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1458 mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1459 smpl_switch_1/smpl_switch_1/Vout mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1460 mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1461 mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1462 mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1463 mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1464 smpl_switch_1/smpl_switch_1/Vout mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1465 mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1466 mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1467 mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1468 mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1469 smpl_switch_1/smpl_switch_1/Vout mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1470 mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1471 mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1472 mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1473 mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1474 smpl_switch_1/smpl_switch_1/Vout mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1475 mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1476 mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1477 mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1478 mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1479 smpl_switch_1/smpl_switch_1/Vout mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1480 cap_dum_12/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1481 cap_dum_12/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1482 cap_dum_12/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1483 cap_dum_12/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1484 gnd cap_dum_12/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1485 cap_dum_11/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1486 cap_dum_11/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1487 cap_dum_11/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1488 cap_dum_11/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1489 gnd cap_dum_11/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1490 cap_dum_13/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1491 cap_dum_13/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1492 cap_dum_13/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1493 cap_dum_13/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1494 gnd cap_dum_13/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1495 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1496 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1497 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1498 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1499 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1500 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi21 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1501 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n1 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1502 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n1 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1503 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi11 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1504 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1505 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1506 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1507 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1508 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1509 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1510 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1511 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1512 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1513 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1514 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1515 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1516 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1517 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1518 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1519 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1520 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1521 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1522 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1523 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1524 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1525 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1526 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n4 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1527 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n4 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1528 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi14 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1529 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1530 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi23 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1531 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n3 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1532 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n3 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1533 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi13 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1534 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1535 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1536 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1537 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1538 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1539 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1540 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi20 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1541 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n0 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1542 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n0 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1543 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi10 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1544 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1545 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1546 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1547 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1548 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1549 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1550 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1551 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1552 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1553 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1554 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1555 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1556 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1557 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1558 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1559 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1560 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1561 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1562 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1563 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1564 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1565 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1566 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n4 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1567 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n4 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1568 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi14 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1569 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1570 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi23 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1571 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n3 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1572 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n3 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1573 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi13 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1574 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1575 mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sphi2 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1576 mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sphi2_n gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1577 mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sphi1_n smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1578 mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sphi1 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1579 smpl_switch_1/smpl_switch_1/Vout mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1580 mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1581 mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1582 mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1583 mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1584 smpl_switch_1/smpl_switch_1/Vout mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1585 mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi23 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1586 mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n3 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1587 mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n3 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1588 mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi13 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1589 smpl_switch_1/smpl_switch_1/Vout mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1590 mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1591 mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n4 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1592 mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n4 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1593 mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi14 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1594 smpl_switch_1/smpl_switch_1/Vout mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1595 mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1596 mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1597 mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1598 mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1599 smpl_switch_1/smpl_switch_1/Vout mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1600 mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1601 mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1602 mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1603 mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1604 smpl_switch_1/smpl_switch_1/Vout mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1605 mid_2_0/m4_2410_n9430# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1606 mid_2_0/m4_2410_n9430# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1607 mid_2_0/m4_2410_n9430# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1608 mid_2_0/m4_2410_n9430# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1609 smpl_switch_1/smpl_switch_1/Vout mid_2_0/m4_2410_n9430# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1610 mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1611 mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1612 mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1613 mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1614 smpl_switch_1/smpl_switch_1/Vout mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1615 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi21 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1616 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n1 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1617 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n1 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1618 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi11 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1619 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1620 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1621 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1622 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1623 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1624 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1625 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi23 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1626 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n3 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1627 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n3 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1628 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi13 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1629 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1630 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1631 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n4 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1632 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n4 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1633 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi14 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1634 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1635 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1636 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n5 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1637 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n5 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1638 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi15 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1639 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1640 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1641 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1642 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1643 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1644 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1645 mid_2_0/mid_2_low_0/m4_2410_n9430# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1646 mid_2_0/mid_2_low_0/m4_2410_n9430# phi2_n6 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1647 mid_2_0/mid_2_low_0/m4_2410_n9430# phi1_n6 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1648 mid_2_0/mid_2_low_0/m4_2410_n9430# phi16 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1649 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_low_0/m4_2410_n9430# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1650 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1651 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n7 gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1652 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n7 smpl_switch_1/smpl_switch_2/Vout vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1653 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi17 smpl_switch_1/smpl_switch_2/Vout sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1654 smpl_switch_1/smpl_switch_1/Vout mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1655 cap_dum_14/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1656 cap_dum_14/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1657 cap_dum_14/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1658 cap_dum_14/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1659 gnd cap_dum_14/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1660 cap_dum_15/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1661 cap_dum_15/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1662 cap_dum_15/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1663 cap_dum_15/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1664 gnd cap_dum_15/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1665 dum_vert_50/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1666 dum_vert_50/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1667 dum_vert_50/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1668 dum_vert_50/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1669 gnd dum_vert_50/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1670 dum_vert_51/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1671 dum_vert_51/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1672 dum_vert_51/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1673 dum_vert_51/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1674 gnd dum_vert_51/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1675 dum_vert_40/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1676 dum_vert_40/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1677 dum_vert_40/m1_990_n540# gnd gnd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1678 dum_vert_40/m1_990_n540# vdd gnd sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1679 gnd dum_vert_40/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
