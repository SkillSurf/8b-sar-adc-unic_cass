* SPICE3 file created from mid_6to8.ext - technology: sky130A

X0 8_cap_array_final_0/cap_final_0/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi2 8_cap_array_final_1/cap_final_7/GND SUB sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1 8_cap_array_final_0/cap_final_0/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi2_n 8_cap_array_final_1/cap_final_7/GND 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2 8_cap_array_final_0/cap_final_0/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi1_n 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3 8_cap_array_final_0/cap_final_0/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi1 8_cap_array_final_1/cap_final_7/Vin SUB sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4 8_cap_array_final_1/cap_final_7/com_x 8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X5 8_cap_array_final_0/cap_final_1/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi2 8_cap_array_final_1/cap_final_7/GND SUB sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=4.64 ps=41.28 w=1 l=0.15
X6 8_cap_array_final_0/cap_final_1/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi2_n 8_cap_array_final_1/cap_final_7/GND 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=4.64 ps=41.28 w=1 l=0.15
X7 8_cap_array_final_0/cap_final_1/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi1_n 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=4.64 ps=41.28 w=1 l=0.15
X8 8_cap_array_final_0/cap_final_1/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi1 8_cap_array_final_1/cap_final_7/Vin SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=4.64 ps=41.28 w=1 l=0.15
X9 8_cap_array_final_1/cap_final_7/com_x 8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X10 8_cap_array_final_0/cap_final_2/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi2 8_cap_array_final_1/cap_final_7/GND SUB sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X11 8_cap_array_final_0/cap_final_2/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi2_n 8_cap_array_final_1/cap_final_7/GND 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X12 8_cap_array_final_0/cap_final_2/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi1_n 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X13 8_cap_array_final_0/cap_final_2/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi1 8_cap_array_final_1/cap_final_7/Vin SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X14 8_cap_array_final_1/cap_final_7/com_x 8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X15 8_cap_array_final_0/cap_final_3/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi2 8_cap_array_final_1/cap_final_7/GND SUB sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X16 8_cap_array_final_0/cap_final_3/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi2_n 8_cap_array_final_1/cap_final_7/GND 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X17 8_cap_array_final_0/cap_final_3/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi1_n 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X18 8_cap_array_final_0/cap_final_3/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi1 8_cap_array_final_1/cap_final_7/Vin SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X19 8_cap_array_final_1/cap_final_7/com_x 8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X20 8_cap_array_final_0/cap_final_4/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi2 8_cap_array_final_1/cap_final_7/GND SUB sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X21 8_cap_array_final_0/cap_final_4/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi2_n 8_cap_array_final_1/cap_final_7/GND 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X22 8_cap_array_final_0/cap_final_4/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi1_n 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X23 8_cap_array_final_0/cap_final_4/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi1 8_cap_array_final_1/cap_final_7/Vin SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X24 8_cap_array_final_1/cap_final_7/com_x 8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X25 8_cap_array_final_0/cap_final_5/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi2 8_cap_array_final_1/cap_final_7/GND SUB sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X26 8_cap_array_final_0/cap_final_5/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi2_n 8_cap_array_final_1/cap_final_7/GND 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X27 8_cap_array_final_0/cap_final_5/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi1_n 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X28 8_cap_array_final_0/cap_final_5/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi1 8_cap_array_final_1/cap_final_7/Vin SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X29 8_cap_array_final_1/cap_final_7/com_x 8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X30 8_cap_array_final_0/cap_final_6/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi2 8_cap_array_final_1/cap_final_7/GND SUB sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X31 8_cap_array_final_0/cap_final_6/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi2_n 8_cap_array_final_1/cap_final_7/GND 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X32 8_cap_array_final_0/cap_final_6/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi1_n 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X33 8_cap_array_final_0/cap_final_6/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi1 8_cap_array_final_1/cap_final_7/Vin SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X34 8_cap_array_final_1/cap_final_7/com_x 8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X35 8_cap_array_final_0/cap_final_7/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi2 8_cap_array_final_1/cap_final_7/GND SUB sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X36 8_cap_array_final_0/cap_final_7/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi2_n 8_cap_array_final_1/cap_final_7/GND 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X37 8_cap_array_final_0/cap_final_7/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi1_n 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X38 8_cap_array_final_0/cap_final_7/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi1 8_cap_array_final_1/cap_final_7/Vin SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X39 8_cap_array_final_1/cap_final_7/com_x 8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X40 8_cap_array_final_1/cap_final_0/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi2 8_cap_array_final_1/cap_final_7/GND SUB sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X41 8_cap_array_final_1/cap_final_0/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi2_n 8_cap_array_final_1/cap_final_7/GND 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X42 8_cap_array_final_1/cap_final_0/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi1_n 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X43 8_cap_array_final_1/cap_final_0/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi1 8_cap_array_final_1/cap_final_7/Vin SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X44 8_cap_array_final_1/cap_final_7/com_x 8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X45 8_cap_array_final_1/cap_final_1/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi2 8_cap_array_final_1/cap_final_7/GND SUB sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X46 8_cap_array_final_1/cap_final_1/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi2_n 8_cap_array_final_1/cap_final_7/GND 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X47 8_cap_array_final_1/cap_final_1/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi1_n 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X48 8_cap_array_final_1/cap_final_1/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi1 8_cap_array_final_1/cap_final_7/Vin SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X49 8_cap_array_final_1/cap_final_7/com_x 8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X50 8_cap_array_final_1/cap_final_2/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi2 8_cap_array_final_1/cap_final_7/GND SUB sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X51 8_cap_array_final_1/cap_final_2/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi2_n 8_cap_array_final_1/cap_final_7/GND 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X52 8_cap_array_final_1/cap_final_2/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi1_n 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X53 8_cap_array_final_1/cap_final_2/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi1 8_cap_array_final_1/cap_final_7/Vin SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X54 8_cap_array_final_1/cap_final_7/com_x 8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X55 8_cap_array_final_1/cap_final_3/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi2 8_cap_array_final_1/cap_final_7/GND SUB sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X56 8_cap_array_final_1/cap_final_3/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi2_n 8_cap_array_final_1/cap_final_7/GND 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X57 8_cap_array_final_1/cap_final_3/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi1_n 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X58 8_cap_array_final_1/cap_final_3/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi1 8_cap_array_final_1/cap_final_7/Vin SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X59 8_cap_array_final_1/cap_final_7/com_x 8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X60 8_cap_array_final_1/cap_final_4/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi2 8_cap_array_final_1/cap_final_7/GND SUB sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X61 8_cap_array_final_1/cap_final_4/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi2_n 8_cap_array_final_1/cap_final_7/GND 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X62 8_cap_array_final_1/cap_final_4/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi1_n 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X63 8_cap_array_final_1/cap_final_4/m1_990_n540# 8_cap_array_final_1/cap_final_4/phi1 8_cap_array_final_1/cap_final_7/Vin SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X64 8_cap_array_final_1/cap_final_7/com_x 8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X65 8_cap_array_final_1/cap_final_5/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi2 8_cap_array_final_1/cap_final_7/GND SUB sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X66 8_cap_array_final_1/cap_final_5/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi2_n 8_cap_array_final_1/cap_final_7/GND 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X67 8_cap_array_final_1/cap_final_5/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi1_n 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X68 8_cap_array_final_1/cap_final_5/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi1 8_cap_array_final_1/cap_final_7/Vin SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X69 8_cap_array_final_1/cap_final_7/com_x 8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X70 8_cap_array_final_1/cap_final_6/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi2 8_cap_array_final_1/cap_final_7/GND SUB sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X71 8_cap_array_final_1/cap_final_6/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi2_n 8_cap_array_final_1/cap_final_7/GND 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X72 8_cap_array_final_1/cap_final_6/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi1_n 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X73 8_cap_array_final_1/cap_final_6/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi1 8_cap_array_final_1/cap_final_7/Vin SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X74 8_cap_array_final_1/cap_final_7/com_x 8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X75 8_cap_array_final_1/cap_final_7/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi2 8_cap_array_final_1/cap_final_7/GND SUB sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X76 8_cap_array_final_1/cap_final_7/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi2_n 8_cap_array_final_1/cap_final_7/GND 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X77 8_cap_array_final_1/cap_final_7/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi1_n 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X78 8_cap_array_final_1/cap_final_7/m1_990_n540# 8_cap_array_final_1/cap_final_7/phi1 8_cap_array_final_1/cap_final_7/Vin SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X79 8_cap_array_final_1/cap_final_7/com_x 8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
C0 8_cap_array_final_1/cap_final_1/m1_990_n540# 8_cap_array_final_1/cap_final_7/com_x 4.980186f
C1 8_cap_array_final_1/cap_final_4/phi1_n 8_cap_array_final_1/cap_final_4/phi2_n 3.503955f
C2 8_cap_array_final_1/cap_final_7/Vdd 8_cap_array_final_1/cap_final_7/GND 17.829754f
C3 8_cap_array_final_1/cap_final_7/phi1_n 8_cap_array_final_1/cap_final_7/Vin 2.491869f
C4 8_cap_array_final_1/cap_final_7/Vdd 8_cap_array_final_1/cap_final_4/phi2_n 2.025186f
C5 8_cap_array_final_1/cap_final_7/phi1_n 8_cap_array_final_1/cap_final_7/phi2_n 2.458625f
C6 8_cap_array_final_0/cap_final_6/m1_990_n540# 8_cap_array_final_1/cap_final_7/com_x 5.002494f
C7 8_cap_array_final_1/cap_final_7/Vdd 8_cap_array_final_1/cap_final_4/phi1_n 2.260308f
C8 8_cap_array_final_1/cap_final_2/m1_990_n540# 8_cap_array_final_1/cap_final_7/com_x 5.002493f
C9 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/GND 13.130507f
C10 8_cap_array_final_1/cap_final_4/phi2 8_cap_array_final_1/m1_n130_2110# 8.66167f
C11 8_cap_array_final_1/m1_n130_1870# 8_cap_array_final_1/m1_n130_1990# 8.59886f
C12 8_cap_array_final_1/cap_final_7/phi2_n 8_cap_array_final_1/cap_final_4/phi2_n 8.877353f
C13 8_cap_array_final_1/m1_n130_1750# 8_cap_array_final_1/m1_n130_1870# 8.59886f
C14 8_cap_array_final_0/cap_final_1/m1_990_n540# 8_cap_array_final_1/cap_final_7/com_x 5.002494f
C15 8_cap_array_final_1/cap_final_7/phi2 8_cap_array_final_1/cap_final_4/phi2 8.88377f
C16 8_cap_array_final_0/cap_final_3/m1_990_n540# 8_cap_array_final_1/cap_final_7/com_x 5.002493f
C17 8_cap_array_final_1/cap_final_3/m1_990_n540# 8_cap_array_final_1/cap_final_7/com_x 5.002493f
C18 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_4/phi1_n 2.030011f
C19 8_cap_array_final_1/cap_final_7/Vdd 8_cap_array_final_1/cap_final_7/Vin 2.515294f
C20 8_cap_array_final_1/m1_n130_4220# 8_cap_array_final_1/m1_n130_4340# 8.59886f
C21 8_cap_array_final_0/cap_final_0/m1_990_n540# 8_cap_array_final_1/cap_final_7/com_x 4.979833f
C22 8_cap_array_final_0/cap_final_2/m1_990_n540# 8_cap_array_final_1/cap_final_7/com_x 5.002493f
C23 8_cap_array_final_0/cap_final_7/m1_990_n540# 8_cap_array_final_1/cap_final_7/com_x 5.002493f
C24 8_cap_array_final_1/cap_final_7/Vdd 8_cap_array_final_1/cap_final_7/phi2_n 2.0731f
C25 8_cap_array_final_1/cap_final_0/m1_990_n540# 8_cap_array_final_1/cap_final_7/com_x 5.002494f
C26 8_cap_array_final_0/cap_final_4/m1_990_n540# 8_cap_array_final_1/cap_final_7/com_x 5.002494f
C27 8_cap_array_final_1/cap_final_5/m1_990_n540# 8_cap_array_final_1/cap_final_7/com_x 5.002494f
C28 8_cap_array_final_1/m1_n130_1630# 8_cap_array_final_1/m1_n130_1750# 8.59886f
C29 8_cap_array_final_1/cap_final_4/phi1 8_cap_array_final_1/cap_final_7/phi1 8.870674f
C30 8_cap_array_final_1/m1_n130_4220# 8_cap_array_final_1/m1_n130_4100# 8.59886f
C31 8_cap_array_final_1/cap_final_7/Vin 8_cap_array_final_1/cap_final_7/phi2_n 15.316741f
C32 8_cap_array_final_1/cap_final_6/m1_990_n540# 8_cap_array_final_1/cap_final_7/com_x 5.002494f
C33 8_cap_array_final_1/m1_n130_4460# 8_cap_array_final_1/m1_n130_4340# 8.59886f
C34 8_cap_array_final_1/cap_final_7/m1_990_n540# 8_cap_array_final_1/cap_final_7/com_x 5.002493f
C35 8_cap_array_final_1/m1_n130_2110# 8_cap_array_final_1/m1_n130_1990# 8.59886f
C36 8_cap_array_final_1/cap_final_7/phi1_n 8_cap_array_final_1/cap_final_4/phi1_n 8.855645f
C37 8_cap_array_final_1/cap_final_7/phi1_n 8_cap_array_final_1/cap_final_7/Vdd 3.189947f
C38 8_cap_array_final_1/cap_final_4/phi1 8_cap_array_final_1/cap_final_4/phi2 3.359025f
C39 8_cap_array_final_1/cap_final_4/phi2_n 8_cap_array_final_1/m1_n130_3980# 8.661217f
C40 8_cap_array_final_1/cap_final_4/m1_990_n540# 8_cap_array_final_1/cap_final_7/com_x 5.002494f
C41 8_cap_array_final_1/cap_final_7/phi2 8_cap_array_final_1/cap_final_7/phi1 2.316001f
C42 8_cap_array_final_0/cap_final_5/m1_990_n540# 8_cap_array_final_1/cap_final_7/com_x 5.002494f
C43 8_cap_array_final_1/m1_n130_4100# 8_cap_array_final_1/m1_n130_3980# 8.59886f
C44 8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C45 8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.340515f **FLOATING
C46 8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.340515f **FLOATING
C47 8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.34045f **FLOATING
C48 8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.34045f **FLOATING
C49 8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.34045f **FLOATING
C50 8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.337859f **FLOATING
C51 8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.34045f **FLOATING
C52 8_cap_array_final_1/m1_n130_1630# SUB 6.902993f
C53 8_cap_array_final_1/m1_n130_1750# SUB 2.161048f
C54 8_cap_array_final_1/m1_n130_1870# SUB 2.165453f
C55 8_cap_array_final_1/m1_n130_1990# SUB 2.174098f
C56 8_cap_array_final_1/m1_n130_2110# SUB 2.192258f
C57 8_cap_array_final_1/cap_final_4/phi2_n SUB 4.644181f
C58 8_cap_array_final_1/m1_n130_3980# SUB 2.149859f
C59 8_cap_array_final_1/m1_n130_4100# SUB 2.152169f
C60 8_cap_array_final_1/m1_n130_4220# SUB 2.152169f
C61 8_cap_array_final_1/m1_n130_4340# SUB 2.152169f
C62 8_cap_array_final_1/m1_n130_4460# SUB 6.896649f
C63 8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.34045f **FLOATING
C64 8_cap_array_final_0/cap_final_6/m1_990_n540# SUB 3.34045f **FLOATING
C65 8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.34045f **FLOATING
C66 8_cap_array_final_1/cap_final_4/phi1 SUB 7.006198f
C67 8_cap_array_final_1/cap_final_4/phi1_n SUB 5.552203f
C68 8_cap_array_final_1/cap_final_4/phi2 SUB 6.49607f
C69 8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.340515f **FLOATING
C70 8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.340515f **FLOATING
C71 8_cap_array_final_1/cap_final_7/phi2 SUB 20.081455f
C72 8_cap_array_final_1/cap_final_7/phi2_n SUB 2.4866f
C73 8_cap_array_final_1/cap_final_7/com_x SUB 6.880803f
C74 8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C75 8_cap_array_final_1/cap_final_7/Vin SUB 6.648837f
C76 8_cap_array_final_1/cap_final_7/Vdd SUB 27.949762f
C77 8_cap_array_final_1/cap_final_7/GND SUB 6.423724f
C78 8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.34045f **FLOATING
C79 8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.339785f **FLOATING
C80 8_cap_array_final_1/cap_final_7/phi1 SUB 7.405069f
C81 8_cap_array_final_1/cap_final_7/phi1_n SUB 4.957194f
