* SPICE3 file created from dac_top_name.ext - technology: sky130A

X0 mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1 mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2 mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3 mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X5 mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=74.24 ps=660.48 w=1 l=0.15
X6 mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=74.24 ps=660.48 w=1 l=0.15
X7 mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=74.24 ps=660.48 w=1 l=0.15
X8 mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=74.24 ps=660.48 w=1 l=0.15
X9 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X10 mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X11 mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X12 mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X13 mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X14 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X15 mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X16 mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X17 mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X18 mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X19 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X20 mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X21 mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X22 mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X23 mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X24 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X25 mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X26 mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n4 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X27 mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n4 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X28 mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi14 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X29 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X30 mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X31 mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X32 mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X33 mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X34 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X35 mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X36 mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X37 mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X38 mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X39 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X40 mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X41 mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X42 mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X43 mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X44 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X45 mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X46 mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X47 mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X48 mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X49 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X50 mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X51 mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X52 mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X53 mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X54 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X55 mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X56 mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X57 mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X58 mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X59 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X60 mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X61 mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n4 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X62 mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n4 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X63 mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi14 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X64 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X65 mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X66 mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X67 mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X68 mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X69 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X70 mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X71 mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X72 mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X73 mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X74 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X75 mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X76 mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X77 mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X78 mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X79 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X80 mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X81 mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X82 mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X83 mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X84 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X85 mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X86 mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X87 mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X88 mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X89 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X90 mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X91 mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X92 mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X93 mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X94 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X95 mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X96 mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X97 mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X98 mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X99 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X100 mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X101 mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X102 mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X103 mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X104 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X105 mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X106 mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n4 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X107 mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n4 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X108 mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi14 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X109 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X110 mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X111 mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X112 mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X113 mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X114 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X115 mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X116 mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X117 mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X118 mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X119 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X120 mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X121 mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X122 mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X123 mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X124 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X125 mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X126 mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X127 mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X128 mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X129 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X130 mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X131 mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X132 mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X133 mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X134 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X135 mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X136 mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X137 mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X138 mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X139 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X140 mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X141 mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n4 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X142 mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n4 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X143 mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi14 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X144 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X145 mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X146 mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X147 mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X148 mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X149 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X150 mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X151 mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X152 mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X153 mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X154 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X155 mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X156 mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X157 mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X158 mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X159 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X160 mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X161 mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X162 mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X163 mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X164 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X165 mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X166 mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X167 mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X168 mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X169 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X170 mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X171 mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X172 mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X173 mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X174 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X175 mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X176 mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X177 mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X178 mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X179 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X180 mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X181 mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X182 mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X183 mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X184 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X185 mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X186 mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n4 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X187 mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n4 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X188 mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi14 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X189 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X190 mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X191 mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X192 mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X193 mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X194 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X195 mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X196 mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X197 mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X198 mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X199 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X200 mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X201 mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X202 mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X203 mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X204 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X205 mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X206 mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X207 mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X208 mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X209 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X210 mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X211 mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X212 mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X213 mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X214 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X215 mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X216 mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X217 mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X218 mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X219 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X220 mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X221 mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n4 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X222 mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n4 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X223 mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi14 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X224 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X225 mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X226 mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X227 mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X228 mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X229 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X230 mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X231 mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X232 mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X233 mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X234 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X235 mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X236 mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X237 mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X238 mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X239 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X240 mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X241 mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X242 mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X243 mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X244 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X245 mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X246 mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X247 mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X248 mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X249 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X250 mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X251 mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X252 mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X253 mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X254 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X255 mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X256 mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X257 mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X258 mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X259 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X260 mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X261 mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X262 mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X263 mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X264 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X265 mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X266 mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n4 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X267 mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n4 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X268 mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi14 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X269 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X270 mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X271 mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X272 mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X273 mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X274 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X275 mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X276 mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X277 mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X278 mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X279 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X280 mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X281 mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X282 mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X283 mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X284 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X285 mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X286 mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X287 mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X288 mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X289 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X290 mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X291 mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X292 mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X293 mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X294 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X295 mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X296 mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X297 mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X298 mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X299 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X300 mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X301 mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n4 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X302 mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n4 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X303 mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi14 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X304 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X305 mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X306 mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X307 mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X308 mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X309 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X310 mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X311 mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X312 mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X313 mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X314 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X315 mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X316 mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X317 mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X318 mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X319 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X320 mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X321 mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X322 mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X323 mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X324 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X325 mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi23 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X326 mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n3 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X327 mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n3 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X328 mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi13 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X329 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X330 mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X331 mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X332 mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X333 mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X334 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X335 mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X336 mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X337 mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X338 mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X339 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X340 mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X341 mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X342 mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X343 mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X344 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X345 mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X346 mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X347 mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X348 mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X349 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X350 mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X351 mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n4 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X352 mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n4 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X353 mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi14 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X354 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X355 mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi22 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X356 mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n2 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X357 mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n2 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X358 mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi12 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X359 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X360 mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi23 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X361 mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n3 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X362 mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n3 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X363 mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi13 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X364 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X365 mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X366 mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X367 mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X368 mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X369 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X370 mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi22 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X371 mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n2 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X372 mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n2 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X373 mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi12 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X374 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X375 mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X376 mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n4 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X377 mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n4 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X378 mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi14 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X379 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X380 mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X381 mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X382 mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X383 mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X384 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X385 mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X386 mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X387 mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X388 mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X389 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X390 mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X391 mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X392 mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X393 mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X394 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X395 mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X396 mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X397 mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X398 mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X399 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X400 mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X401 mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X402 mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X403 mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X404 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X405 mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi23 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X406 mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n3 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X407 mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n3 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X408 mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi13 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X409 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X410 mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X411 mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X412 mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X413 mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X414 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X415 mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X416 mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X417 mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X418 mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X419 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X420 mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X421 mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X422 mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X423 mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X424 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X425 mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X426 mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X427 mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X428 mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X429 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X430 mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X431 mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n4 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X432 mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n4 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X433 mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi14 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X434 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X435 mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi22 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X436 mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n2 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X437 mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n2 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X438 mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi12 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X439 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X440 mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi23 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X441 mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n3 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X442 mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n3 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X443 mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi13 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X444 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X445 mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X446 mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X447 mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X448 mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X449 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X450 mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi22 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X451 mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n2 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X452 mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n2 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X453 mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi12 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X454 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X455 mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X456 mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n4 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X457 mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n4 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X458 mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi14 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X459 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X460 mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X461 mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X462 mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X463 mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X464 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X465 mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X466 mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X467 mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X468 mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X469 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X470 mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X471 mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X472 mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X473 mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X474 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X475 mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X476 mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X477 mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X478 mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X479 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X480 mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X481 mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X482 mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X483 mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X484 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X485 mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X486 mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X487 mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X488 mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X489 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X490 mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X491 mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X492 mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X493 mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X494 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X495 mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X496 mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X497 mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X498 mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X499 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X500 mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X501 mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X502 mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X503 mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X504 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X505 mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X506 mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X507 mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X508 mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X509 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X510 mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X511 mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X512 mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X513 mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X514 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X515 mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X516 mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X517 mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X518 mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X519 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X520 mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X521 mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X522 mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X523 mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X524 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X525 mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X526 mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X527 mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X528 mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X529 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X530 mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X531 mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X532 mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X533 mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X534 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X535 mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X536 mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X537 mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X538 mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X539 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X540 mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X541 mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X542 mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X543 mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X544 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X545 mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X546 mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X547 mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X548 mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X549 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X550 mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X551 mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X552 mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X553 mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X554 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X555 mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X556 mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X557 mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X558 mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X559 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X560 end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X561 end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X562 end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X563 end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X564 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X565 end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X566 end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X567 end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X568 end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X569 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X570 end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X571 end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X572 end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X573 end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X574 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X575 end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X576 end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X577 end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X578 end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X579 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X580 end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X581 end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X582 end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X583 end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X584 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X585 end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X586 end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X587 end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X588 end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X589 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X590 end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X591 end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X592 end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X593 end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X594 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X595 end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X596 end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X597 end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X598 end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X599 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X600 end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X601 end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X602 end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X603 end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X604 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X605 end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X606 end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X607 end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X608 end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X609 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X610 end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X611 end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X612 end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X613 end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X614 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X615 end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X616 end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X617 end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X618 end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X619 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X620 end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X621 end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X622 end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X623 end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X624 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X625 end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X626 end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X627 end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X628 end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X629 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X630 end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X631 end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X632 end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X633 end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X634 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X635 end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X636 end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X637 end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X638 end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X639 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X640 mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X641 mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X642 mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X643 mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X644 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X645 mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X646 mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X647 mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X648 mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X649 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X650 mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X651 mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X652 mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X653 mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X654 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X655 mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X656 mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X657 mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X658 mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X659 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X660 mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X661 mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X662 mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X663 mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X664 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X665 mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X666 mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X667 mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X668 mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X669 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X670 mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X671 mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X672 mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X673 mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X674 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X675 mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X676 mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X677 mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X678 mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X679 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X680 mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X681 mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X682 mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X683 mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X684 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X685 mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X686 mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X687 mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X688 mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X689 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X690 mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X691 mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X692 mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X693 mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X694 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X695 mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X696 mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X697 mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X698 mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X699 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X700 mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X701 mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X702 mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X703 mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X704 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X705 mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X706 mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X707 mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X708 mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X709 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X710 mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X711 mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X712 mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X713 mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X714 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X715 mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X716 mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X717 mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X718 mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X719 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X720 end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X721 end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X722 end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X723 end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X724 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X725 end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X726 end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X727 end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X728 end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X729 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X730 end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X731 end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X732 end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X733 end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X734 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X735 end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X736 end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X737 end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X738 end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X739 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X740 end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X741 end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X742 end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X743 end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X744 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X745 end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X746 end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X747 end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X748 end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X749 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X750 end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X751 end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X752 end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X753 end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X754 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X755 end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X756 end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X757 end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X758 end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X759 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X760 end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X761 end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X762 end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X763 end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X764 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X765 end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X766 end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X767 end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X768 end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X769 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X770 end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X771 end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X772 end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X773 end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X774 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X775 end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X776 end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X777 end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X778 end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X779 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X780 end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X781 end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X782 end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X783 end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X784 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X785 end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X786 end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X787 end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X788 end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X789 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X790 end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X791 end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X792 end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X793 end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X794 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X795 end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X796 end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X797 end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X798 end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X799 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X800 end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X801 end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X802 end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X803 end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X804 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X805 end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X806 end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X807 end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X808 end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X809 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X810 end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X811 end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X812 end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X813 end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X814 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X815 end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X816 end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X817 end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X818 end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X819 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X820 end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X821 end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X822 end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X823 end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X824 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X825 end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X826 end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X827 end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X828 end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X829 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X830 end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X831 end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X832 end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X833 end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X834 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X835 end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X836 end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X837 end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X838 end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X839 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X840 end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X841 end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X842 end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X843 end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X844 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X845 end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X846 end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X847 end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X848 end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X849 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X850 end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X851 end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X852 end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X853 end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X854 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X855 end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X856 end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X857 end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X858 end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X859 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X860 end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X861 end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X862 end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X863 end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X864 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X865 end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X866 end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X867 end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X868 end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X869 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X870 end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X871 end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X872 end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X873 end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X874 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X875 end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X876 end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X877 end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X878 end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X879 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X880 mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X881 mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X882 mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X883 mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X884 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X885 mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X886 mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X887 mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X888 mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X889 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X890 mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X891 mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X892 mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X893 mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X894 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X895 mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X896 mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X897 mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X898 mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X899 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X900 mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X901 mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X902 mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X903 mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X904 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X905 mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X906 mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X907 mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X908 mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X909 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X910 mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X911 mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X912 mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X913 mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X914 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X915 mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X916 mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X917 mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X918 mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X919 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X920 mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X921 mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X922 mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X923 mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X924 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X925 mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X926 mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X927 mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X928 mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X929 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X930 mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X931 mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X932 mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X933 mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X934 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X935 mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X936 mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X937 mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X938 mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X939 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X940 mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X941 mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X942 mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X943 mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X944 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X945 mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X946 mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X947 mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X948 mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X949 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X950 mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X951 mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X952 mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X953 mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X954 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X955 mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X956 mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X957 mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X958 mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X959 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X960 end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X961 end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X962 end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X963 end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X964 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X965 end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X966 end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X967 end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X968 end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X969 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X970 end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X971 end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X972 end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X973 end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X974 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X975 end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X976 end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X977 end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X978 end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X979 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X980 end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X981 end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X982 end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X983 end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X984 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X985 end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X986 end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X987 end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X988 end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X989 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X990 end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X991 end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X992 end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X993 end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X994 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X995 end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X996 end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X997 end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X998 end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X999 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1000 end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1001 end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1002 end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1003 end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1004 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1005 end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1006 end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1007 end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1008 end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1009 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1010 end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1011 end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1012 end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1013 end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1014 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1015 end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1016 end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1017 end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1018 end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1019 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1020 end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1021 end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1022 end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1023 end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1024 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1025 end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1026 end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1027 end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1028 end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1029 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1030 end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1031 end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1032 end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1033 end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1034 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1035 end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1036 end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1037 end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1038 end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1039 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1040 mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1041 mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1042 mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1043 mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1044 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1045 mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1046 mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1047 mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1048 mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1049 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1050 mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1051 mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1052 mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1053 mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1054 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1055 mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1056 mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1057 mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1058 mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1059 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1060 mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1061 mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1062 mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1063 mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1064 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1065 mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1066 mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1067 mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1068 mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1069 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1070 mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1071 mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1072 mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1073 mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1074 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1075 mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1076 mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1077 mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1078 mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1079 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1080 mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1081 mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1082 mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1083 mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1084 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1085 mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1086 mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1087 mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1088 mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1089 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1090 mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1091 mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1092 mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1093 mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1094 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1095 mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1096 mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1097 mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1098 mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1099 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1100 mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1101 mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1102 mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1103 mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1104 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1105 mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1106 mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1107 mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1108 mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1109 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1110 mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1111 mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1112 mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1113 mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1114 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1115 mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1116 mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1117 mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1118 mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1119 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1120 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1121 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1122 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1123 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1124 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1125 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi21 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1126 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n1 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1127 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n1 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1128 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# phi11 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1129 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1130 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1131 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1132 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1133 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1134 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1135 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1136 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1137 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1138 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1139 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1140 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1141 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1142 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1143 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1144 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1145 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1146 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1147 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1148 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1149 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1150 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1151 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n4 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1152 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n4 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1153 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# phi14 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1154 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1155 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi23 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1156 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n3 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1157 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n3 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1158 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# phi13 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1159 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1160 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1161 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1162 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1163 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1164 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1165 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi20 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1166 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi2_n0 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1167 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi1_n0 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1168 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# phi10 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1169 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1170 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1171 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1172 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1173 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1174 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1175 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1176 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1177 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1178 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1179 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1180 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1181 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1182 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1183 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1184 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1185 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1186 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1187 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1188 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1189 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1190 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1191 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi2_n4 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1192 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi1_n4 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1193 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# phi14 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1194 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1195 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi23 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1196 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi2_n3 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1197 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi1_n3 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1198 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# phi13 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1199 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1200 mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# smpl_n_d12 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1201 mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# smpl_n_d12_out_n gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1202 mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_0/phi1_n vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1203 mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# smpl vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1204 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1205 mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1206 mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1207 mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1208 mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1209 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1210 mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi23 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1211 mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n3 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1212 mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n3 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1213 mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi13 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1214 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1215 mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1216 mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n4 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1217 mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n4 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1218 mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi14 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1219 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1220 mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1221 mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1222 mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1223 mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1224 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1225 mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1226 mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1227 mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1228 mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1229 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1230 mid_2_0/m4_2410_n9430# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1231 mid_2_0/m4_2410_n9430# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1232 mid_2_0/m4_2410_n9430# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1233 mid_2_0/m4_2410_n9430# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1234 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/m4_2410_n9430# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1235 mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1236 mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1237 mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1238 mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1239 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1240 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi21 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1241 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi2_n1 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1242 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi1_n1 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1243 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# phi11 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1244 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1245 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1246 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1247 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1248 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1249 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1250 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi23 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1251 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi2_n3 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1252 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi1_n3 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1253 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# phi13 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1254 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1255 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi24 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1256 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi2_n4 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1257 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi1_n4 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1258 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# phi14 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1259 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1260 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi25 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1261 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi2_n5 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1262 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi1_n5 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1263 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# phi15 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1264 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1265 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1266 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1267 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1268 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1269 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1270 mid_2_0/mid_2_low_0/m4_2410_n9430# phi26 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1271 mid_2_0/mid_2_low_0/m4_2410_n9430# phi2_n6 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1272 mid_2_0/mid_2_low_0/m4_2410_n9430# phi1_n6 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1273 mid_2_0/mid_2_low_0/m4_2410_n9430# phi16 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1274 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/m4_2410_n9430# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1275 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi27 gnd sub sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1276 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi2_n7 gnd Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1277 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi1_n7 vin Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1278 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# phi17 vin sub sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1279 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
C0 mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C1 mid_6to8_3/8_cap_array_final_1/m1_n130_1870# mid_6to8_3/8_cap_array_final_1/m1_n130_1750# 8.59886f
C2 phi13 phi14 20.084393f
C3 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# 5.002839f
C4 mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C5 phi26 mid_6to8_2/8_cap_array_final_1/m1_n130_2110# 8.66467f
C6 phi1_n4 phi2_n4 50.327557f
C7 phi14 phi24 64.99351f
C8 vin phi1_n5 7.361336f
C9 phi17 gnd 2.178203f
C10 Vdd phi2_n5 8.281558f
C11 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# 5.002839f
C12 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# 5.002838f
C13 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C14 mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C15 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# 5.002838f
C16 end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C17 end_2/8_cap_array_final_1/m1_n130_4460# end_2/8_cap_array_final_1/m1_n130_4340# 8.59886f
C18 mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C19 mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C20 mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C21 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C22 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# 5.002838f
C23 end_1/8_cap_array_final_1/m1_n130_1750# end_1/8_cap_array_final_1/m1_n130_1630# 8.59886f
C24 end_0/8_cap_array_final_1/m1_n130_1870# end_0/8_cap_array_final_1/m1_n130_1750# 8.59886f
C25 mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C26 mid_4to8_2/8_cap_array_final_1/m1_n130_4460# mid_4to8_2/8_cap_array_final_1/m1_n130_4340# 8.59886f
C27 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# 5.002494f
C28 phi2_n0 phi20 2.616692f
C29 end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C30 end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C31 mid_6to8_3/8_cap_array_final_1/m1_n130_1750# mid_6to8_3/8_cap_array_final_1/m1_n130_1630# 8.59886f
C32 end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C33 phi27 end_3/8_cap_array_final_1/m1_n130_2230# 8.728627f
C34 mid_6to8_2/8_cap_array_final_1/m1_n130_2110# mid_6to8_2/8_cap_array_final_1/m1_n130_1990# 8.59886f
C35 mid_4to8_3/8_cap_array_final_1/m1_n130_4340# mid_4to8_3/8_cap_array_final_1/m1_n130_4460# 8.59886f
C36 phi14 phi12 19.728592f
C37 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# 5.002838f
C38 phi1_n3 phi1_n2 18.339928f
C39 mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C40 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C41 gnd phi1_n7 12.560539f
C42 mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C43 phi15 phi25 69.67804f
C44 phi11 phi1_n1 2.693908f
C45 mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C46 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# 5.002839f
C47 mid_2to4__1/8_cap_array_final_1/m1_n130_1630# phi23 8.62096f
C48 phi2_n1 smpl_n_d12_out_n 9.007117f
C49 phi2_n4 Vdd 4.265811f
C50 vin mid_2_0/8_cap_array_final_0/cap_final_0/phi1_n 22.264622f
C51 phi2_n3 phi2_n2 17.995602f
C52 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# 5.002839f
C53 mid_4to8_1/8_cap_array_final_1/m1_n130_1870# phi25 8.649647f
C54 mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C55 phi13 phi24 2.68972f
C56 phi2_n3 phi2_n0 9.046399f
C57 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# 5.002838f
C58 phi1_n4 phi1_n3 20.080708f
C59 phi27 end_1/8_cap_array_final_1/m1_n130_2230# 8.728627f
C60 end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C61 end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C62 phi14 phi23 37.595497f
C63 mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C64 mid_6to8_1/8_cap_array_final_1/m1_n130_4220# mid_6to8_1/8_cap_array_final_1/m1_n130_4100# 8.59886f
C65 smpl_n_d12 smpl_n_d12_out_n 2.639232f
C66 phi23 phi20 9.051891f
C67 mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C68 end_0/8_cap_array_final_1/m1_n130_1750# end_0/8_cap_array_final_1/m1_n130_1630# 8.59886f
C69 phi14 phi25 6.49583f
C70 phi21 phi20 8.979368f
C71 mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C72 phi2_n6 phi1_n7 28.057055f
C73 mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C74 mid_4to8_3/8_cap_array_final_1/m1_n130_1870# mid_4to8_3/8_cap_array_final_1/m1_n130_1750# 8.59886f
C75 mid_6to8_2/8_cap_array_final_1/m1_n130_1990# mid_6to8_2/8_cap_array_final_1/m1_n130_1870# 8.59886f
C76 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# 5.272134f
C77 mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C78 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# 5.272134f
C79 end_3/8_cap_array_final_1/cap_final_7/com_x Vdd 2.644652f
C80 mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C81 phi2_n7 end_1/8_cap_array_final_1/m1_n130_3860# 8.726839f
C82 phi1_n6 phi2_n5 24.056414f
C83 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# 5.002839f
C84 end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272134f
C85 phi13 phi12 18.34155f
C86 phi2_n3 phi23 3.018898f
C87 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C88 phi1_n7 phi2_n7 83.35087f
C89 gnd vin 0.234499p
C90 phi12 phi24 2.222702f
C91 end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C92 mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C93 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# 5.002838f
C94 end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C95 mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C96 phi1_n3 Vdd 2.178562f
C97 mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C98 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# 5.002838f
C99 mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272134f
C100 mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C101 mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272134f
C102 mid_4to8_2/8_cap_array_final_1/m1_n130_4220# mid_4to8_2/8_cap_array_final_1/m1_n130_4340# 8.59886f
C103 mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C104 phi13 phi23 52.877754f
C105 mid_4to8_3/8_cap_array_final_1/m1_n130_1750# mid_4to8_3/8_cap_array_final_1/m1_n130_1630# 8.59886f
C106 mid_6to8_2/8_cap_array_final_1/m1_n130_1870# mid_6to8_2/8_cap_array_final_1/m1_n130_1750# 8.59886f
C107 phi2_n6 mid_6to8_2/8_cap_array_final_1/m1_n130_3980# 8.664217f
C108 phi16 phi27 21.651308f
C109 mid_4to8_1/8_cap_array_final_1/m1_n130_4220# phi2_n5 8.649531f
C110 phi2_n6 phi1_n5 7.061357f
C111 smpl mid_2_0/8_cap_array_final_0/cap_final_0/phi1_n 2.612654f
C112 mid_6to8_3/8_cap_array_final_1/m1_n130_3980# mid_6to8_3/8_cap_array_final_1/m1_n130_4100# 8.59886f
C113 phi23 phi24 18.28477f
C114 mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C115 phi26 phi27 0.108955p
C116 mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C117 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# 5.002838f
C118 end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002494f
C119 phi2_n6 vin 2.262305f
C120 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# 5.002839f
C121 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# 5.002839f
C122 mid_6to8_2/8_cap_array_final_1/m1_n130_4340# mid_6to8_2/8_cap_array_final_1/m1_n130_4220# 8.59886f
C123 end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C124 phi1_n4 phi1_n7 2.231639f
C125 phi1_n0 phi2_n0 25.457558f
C126 phi25 phi24 72.199745f
C127 mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C128 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# 5.002838f
C129 phi2_n3 phi2_n1 9.101527f
C130 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# 5.002839f
C131 end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C132 end_3/8_cap_array_final_1/m1_n130_4340# end_3/8_cap_array_final_1/m1_n130_4220# 8.59886f
C133 end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.27179f
C134 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# 5.002838f
C135 mid_6to8_2/8_cap_array_final_1/m1_n130_3980# mid_6to8_2/8_cap_array_final_1/m1_n130_4100# 8.59886f
C136 mid_6to8_1/8_cap_array_final_1/m1_n130_3980# mid_6to8_1/8_cap_array_final_1/m1_n130_4100# 8.59886f
C137 phi17 Vdd 4.889181f
C138 end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C139 mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C140 mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C141 phi16 phi1_n6 4.236728f
C142 vin phi2_n7 0.246419p
C143 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# 5.002494f
C144 mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C145 end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C146 phi1_n4 phi14 3.267454f
C147 end_1/8_cap_array_final_1/m1_n130_4460# end_1/8_cap_array_final_1/m1_n130_4340# 8.59886f
C148 mid_6to8_2/8_cap_array_final_1/m1_n130_1750# mid_6to8_2/8_cap_array_final_1/m1_n130_1630# 8.59886f
C149 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# 5.002493f
C150 phi12 phi21 36.954197f
C151 phi1_n1 phi1_n3 9.312764f
C152 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# 5.002838f
C153 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# 5.272134f
C154 phi2_n4 phi2_n5 72.16842f
C155 mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272134f
C156 end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.979833f
C157 phi25 mid_4to8_0/8_cap_array_final_1/m1_n130_1870# 8.649647f
C158 mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C159 mid_6to8_3/8_cap_array_final_1/m1_n130_4220# mid_6to8_3/8_cap_array_final_1/m1_n130_4100# 8.59886f
C160 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C161 phi10 phi20 40.411327f
C162 phi1_n4 phi1_n5 84.23691f
C163 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# 5.272134f
C164 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# 5.002839f
C165 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# 5.002839f
C166 phi1_n7 Vdd 51.499027f
C167 phi23 phi21 9.110596f
C168 mid_4to8_1/8_cap_array_final_1/m1_n130_4340# mid_4to8_1/8_cap_array_final_1/m1_n130_4460# 8.59886f
C169 phi1_n4 phi2_n3 22.606203f
C170 phi1_n4 vin 4.006585f
C171 end_2/8_cap_array_final_1/m1_n130_3980# end_2/8_cap_array_final_1/m1_n130_4100# 8.59886f
C172 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# 5.002839f
C173 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# 5.272134f
C174 end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C175 phi2_n1 phi2_n0 8.973002f
C176 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# 5.002838f
C177 end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C178 phi17 phi27 96.231766f
C179 end_1/8_cap_array_final_1/m1_n130_3980# end_1/8_cap_array_final_1/m1_n130_4100# 8.59886f
C180 phi26 mid_6to8_0/8_cap_array_final_1/m1_n130_2110# 8.66467f
C181 mid_6to8_2/8_cap_array_final_1/m1_n130_4220# mid_6to8_2/8_cap_array_final_1/m1_n130_4100# 8.59886f
C182 mid_6to8_1/8_cap_array_final_1/m1_n130_2110# mid_6to8_1/8_cap_array_final_1/m1_n130_1990# 8.59886f
C183 end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C184 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# 5.002838f
C185 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# 5.002838f
C186 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# 5.002839f
C187 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# 5.002839f
C188 phi2_n2 phi1_n2 29.428595f
C189 mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C190 mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C191 end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C192 mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C193 mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C194 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# 5.002838f
C195 gnd phi2_n6 13.09726f
C196 mid_4to8_1/8_cap_array_final_1/m1_n130_1870# mid_4to8_1/8_cap_array_final_1/m1_n130_1750# 8.59886f
C197 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C198 mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C199 mid_6to8_0/8_cap_array_final_1/m1_n130_1990# mid_6to8_0/8_cap_array_final_1/m1_n130_1870# 8.59886f
C200 end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C201 mid_6to8_3/8_cap_array_final_1/m1_n130_2110# phi26 8.66467f
C202 mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C203 phi13 phi10 9.170131f
C204 Vdd phi1_n5 8.691263f
C205 end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C206 smpl_n_d12 smpl 40.532215f
C207 phi2_n1 phi21 2.753754f
C208 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# 5.002838f
C209 phi12 phi1_n2 2.727744f
C210 phi2_n3 Vdd 2.116855f
C211 mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C212 mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C213 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C214 vin Vdd 48.83908f
C215 gnd phi2_n7 27.94766f
C216 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# 5.002839f
C217 end_2/8_cap_array_final_1/m1_n130_3980# end_2/8_cap_array_final_1/m1_n130_3860# 8.59886f
C218 end_2/8_cap_array_final_1/m1_n130_4220# end_2/8_cap_array_final_1/m1_n130_4100# 8.59886f
C219 mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C220 mid_6to8_1/8_cap_array_final_1/m1_n130_1990# mid_6to8_1/8_cap_array_final_1/m1_n130_1870# 8.59886f
C221 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# 5.002838f
C222 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# 5.002838f
C223 mid_4to8_0/8_cap_array_final_1/m1_n130_4340# mid_4to8_0/8_cap_array_final_1/m1_n130_4220# 8.59886f
C224 smpl_n_d12 phi21 9.010565f
C225 end_1/8_cap_array_final_1/m1_n130_3980# end_1/8_cap_array_final_1/m1_n130_3860# 8.59886f
C226 end_1/8_cap_array_final_1/m1_n130_4220# end_1/8_cap_array_final_1/m1_n130_4100# 8.59886f
C227 end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C228 end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002493f
C229 mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C230 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# 5.002838f
C231 phi16 phi26 83.13197f
C232 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# 5.002838f
C233 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# 5.002838f
C234 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# 5.002839f
C235 mid_6to8_3/8_cap_array_final_1/m1_n130_4220# mid_6to8_3/8_cap_array_final_1/m1_n130_4340# 8.59886f
C236 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C237 mid_4to8_1/8_cap_array_final_1/m1_n130_1750# mid_4to8_1/8_cap_array_final_1/m1_n130_1630# 8.59886f
C238 mid_6to8_0/8_cap_array_final_1/m1_n130_1870# mid_6to8_0/8_cap_array_final_1/m1_n130_1750# 8.59886f
C239 mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C240 phi1_n7 phi1_n6 0.130461p
C241 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C242 end_0/8_cap_array_final_1/m1_n130_3980# end_0/8_cap_array_final_1/m1_n130_4100# 8.59886f
C243 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# 5.002838f
C244 phi1_n3 phi2_n4 2.654304f
C245 phi2_n6 phi2_n7 0.108858p
C246 mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C247 mid_4to8_3/8_cap_array_final_1/m1_n130_1870# phi25 8.649647f
C248 mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C249 mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C250 phi1_n0 phi10 2.606045f
C251 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C252 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# 5.002838f
C253 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# 5.002838f
C254 mid_6to8_1/8_cap_array_final_1/m1_n130_1870# mid_6to8_1/8_cap_array_final_1/m1_n130_1750# 8.59886f
C255 mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C256 end_2/8_cap_array_final_1/m1_n130_2230# end_2/8_cap_array_final_1/m1_n130_2110# 8.59886f
C257 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# 5.002839f
C258 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# 5.002494f
C259 end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C260 mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C261 phi2_n3 mid_2to4__0/8_cap_array_final_1/m1_n130_4460# 8.620945f
C262 end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C263 mid_2_0/mid_2_low_0/m4_2410_n9430# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C264 mid_6to8_0/8_cap_array_final_1/m1_n130_4340# mid_6to8_0/8_cap_array_final_1/m1_n130_4460# 8.59886f
C265 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# 5.002839f
C266 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C267 mid_6to8_0/8_cap_array_final_1/m1_n130_1750# mid_6to8_0/8_cap_array_final_1/m1_n130_1630# 8.59886f
C268 mid_6to8_1/8_cap_array_final_1/m1_n130_4460# mid_6to8_1/8_cap_array_final_1/m1_n130_4340# 8.59886f
C269 mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C270 phi2_n1 phi1_n2 21.987999f
C271 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# 5.002839f
C272 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C273 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C274 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# 5.002838f
C275 mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C276 end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C277 mid_4to8_0/8_cap_array_final_1/m1_n130_4460# mid_4to8_0/8_cap_array_final_1/m1_n130_4340# 8.59886f
C278 phi1_n4 phi2_n6 6.004341f
C279 mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C280 smpl Vdd 37.06365f
C281 mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C282 phi1_n6 phi1_n5 42.957775f
C283 mid_6to8_0/8_cap_array_final_1/m1_n130_1990# mid_6to8_0/8_cap_array_final_1/m1_n130_2110# 8.59886f
C284 mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C285 phi11 phi20 37.760708f
C286 vin phi1_n6 16.566456f
C287 end_0/8_cap_array_final_1/m1_n130_3980# end_0/8_cap_array_final_1/m1_n130_3860# 8.59886f
C288 end_0/8_cap_array_final_1/m1_n130_4220# end_0/8_cap_array_final_1/m1_n130_4100# 8.59886f
C289 mid_4to8_0/8_cap_array_final_1/m1_n130_4220# phi2_n5 8.649531f
C290 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# 5.002839f
C291 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# 5.002838f
C292 gnd Vdd 0.288759p
C293 mid_6to8_1/8_cap_array_final_1/m1_n130_1750# mid_6to8_1/8_cap_array_final_1/m1_n130_1630# 8.59886f
C294 mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C295 mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C296 phi17 phi16 0.130666p
C297 end_2/8_cap_array_final_1/m1_n130_2110# end_2/8_cap_array_final_1/m1_n130_1990# 8.59886f
C298 mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C299 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# 4.980177f
C300 end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002493f
C301 phi17 phi26 43.303696f
C302 phi1_n1 mid_2_0/8_cap_array_final_0/cap_final_0/phi1_n 8.91752f
C303 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# 5.002838f
C304 end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C305 mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C306 phi1_n1 phi2_n0 22.7846f
C307 mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C308 mid_6to8_3/8_cap_array_final_1/m1_n130_4460# mid_6to8_3/8_cap_array_final_1/m1_n130_4340# 8.59886f
C309 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# 5.002839f
C310 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# 5.002838f
C311 phi1_n4 phi1_n2 19.731527f
C312 end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C313 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# 5.002839f
C314 phi2_n5 phi1_n5 55.251938f
C315 end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C316 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# 5.002838f
C317 phi2_n6 Vdd 16.618898f
C318 smpl_n_d12 phi10 36.9208f
C319 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# 5.002839f
C320 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# 5.002838f
C321 phi15 phi16 42.98026f
C322 phi11 phi13 9.289417f
C323 end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C324 mid_4to8_2/8_cap_array_final_1/m1_n130_1870# mid_4to8_2/8_cap_array_final_1/m1_n130_1750# 8.59886f
C325 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# 5.002838f
C326 phi15 phi26 7.159061f
C327 phi1_n0 phi1_n1 8.918006f
C328 mid_6to8_1/8_cap_array_final_1/m1_n130_2110# phi26 8.66467f
C329 end_0/8_cap_array_final_1/m1_n130_2230# phi27 8.728627f
C330 end_2/8_cap_array_final_1/m1_n130_1990# end_2/8_cap_array_final_1/m1_n130_1870# 8.59886f
C331 phi22 phi13 39.22582f
C332 mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C333 end_2/8_cap_array_final_1/m1_n130_3860# phi2_n7 8.726839f
C334 gnd phi27 5.607867f
C335 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# 5.002838f
C336 mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C337 mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C338 mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C339 Vdd phi2_n7 33.527f
C340 phi22 phi24 18.10835f
C341 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# 5.002838f
C342 mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C343 phi16 phi14 42.41868f
C344 end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C345 phi14 phi26 6.085594f
C346 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# 5.002838f
C347 phi2_n4 phi1_n5 28.517515f
C348 mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C349 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# 5.002838f
C350 phi2_n6 mid_6to8_3/8_cap_array_final_1/m1_n130_3980# 8.664217f
C351 phi22 phi2_n2 2.730589f
C352 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# 5.002838f
C353 mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C354 end_3/8_cap_array_final_1/m1_n130_2230# end_3/8_cap_array_final_1/m1_n130_2110# 8.59886f
C355 phi2_n3 phi2_n4 18.272886f
C356 mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272135f
C357 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C358 mid_4to8_2/8_cap_array_final_1/m1_n130_1750# mid_4to8_2/8_cap_array_final_1/m1_n130_1630# 8.59886f
C359 phi23 mid_2to4__0/8_cap_array_final_1/m1_n130_1630# 8.62096f
C360 mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C361 gnd phi1_n6 3.445286f
C362 mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C363 mid_6to8_1/8_cap_array_final_1/m1_n130_4340# mid_6to8_1/8_cap_array_final_1/m1_n130_4220# 8.59886f
C364 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# 5.002838f
C365 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# 5.002494f
C366 mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C367 end_2/8_cap_array_final_1/m1_n130_1870# end_2/8_cap_array_final_1/m1_n130_1750# 8.59886f
C368 phi11 smpl 8.929021f
C369 phi2_n7 end_0/8_cap_array_final_1/m1_n130_3860# 8.726839f
C370 end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C371 mid_6to8_0/8_cap_array_final_1/m1_n130_3980# mid_6to8_0/8_cap_array_final_1/m1_n130_4100# 8.59886f
C372 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272135f
C373 phi1_n4 Vdd 4.686877f
C374 phi22 phi12 44.305923f
C375 mid_4to8_2/8_cap_array_final_1/m1_n130_1870# phi25 8.649647f
C376 mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C377 phi16 vin 3.020648f
C378 mid_2_0/m4_2410_n9430# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C379 mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C380 phi2_n1 phi1_n1 29.470316f
C381 phi2_n4 phi24 3.332905f
C382 mid_4to8_1/8_cap_array_final_1/m1_n130_4340# mid_4to8_1/8_cap_array_final_1/m1_n130_4220# 8.59886f
C383 mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C384 phi27 phi2_n7 5.805571f
C385 phi2_n5 mid_4to8_3/8_cap_array_final_1/m1_n130_4220# 8.649531f
C386 phi11 phi21 44.41444f
C387 mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C388 mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C389 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# 5.002838f
C390 end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C391 phi17 phi15 3.002692f
C392 end_3/8_cap_array_final_1/m1_n130_2110# end_3/8_cap_array_final_1/m1_n130_1990# 8.59886f
C393 phi2_n6 phi1_n6 69.25696f
C394 phi22 phi23 18.010555f
C395 mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272134f
C396 phi17 phi1_n7 24.895061f
C397 end_1/8_cap_array_final_1/m1_n130_2230# end_1/8_cap_array_final_1/m1_n130_2110# 8.59886f
C398 phi2_n2 phi2_n4 18.107841f
C399 gnd phi2_n5 6.603709f
C400 mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C401 end_2/8_cap_array_final_1/m1_n130_4340# end_2/8_cap_array_final_1/m1_n130_4220# 8.59886f
C402 end_2/8_cap_array_final_1/m1_n130_1750# end_2/8_cap_array_final_1/m1_n130_1630# 8.59886f
C403 mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C404 phi26 phi24 36.360214f
C405 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C406 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# 5.002838f
C407 phi25 phi2_n5 3.67012f
C408 end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002493f
C409 mid_4to8_0/8_cap_array_final_1/m1_n130_1870# mid_4to8_0/8_cap_array_final_1/m1_n130_1750# 8.59886f
C410 phi2_n3 phi1_n3 38.04705f
C411 end_1/8_cap_array_final_1/m1_n130_4340# end_1/8_cap_array_final_1/m1_n130_4220# 8.59886f
C412 mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C413 mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C414 phi1_n6 phi2_n7 21.364698f
C415 mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272134f
C416 phi17 phi14 2.300412f
C417 mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C418 end_3/8_cap_array_final_1/m1_n130_3980# end_3/8_cap_array_final_1/m1_n130_4100# 8.59886f
C419 mid_4to8_3/8_cap_array_final_1/m1_n130_4340# mid_4to8_3/8_cap_array_final_1/m1_n130_4220# 8.59886f
C420 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# 5.002838f
C421 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# 5.002838f
C422 mid_6to8_0/8_cap_array_final_1/m1_n130_4220# mid_6to8_0/8_cap_array_final_1/m1_n130_4100# 8.59886f
C423 mid_6to8_0/8_cap_array_final_1/m1_n130_3980# phi2_n6 8.664217f
C424 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# 5.002838f
C425 end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C426 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# 5.002839f
C427 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# 5.002839f
C428 mid_6to8_1/8_cap_array_final_1/m1_n130_3980# phi2_n6 8.664217f
C429 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# 5.002839f
C430 mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C431 mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C432 phi2_n6 phi2_n5 36.905354f
C433 phi13 phi1_n3 2.932781f
C434 mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C435 end_3/8_cap_array_final_1/m1_n130_1990# end_3/8_cap_array_final_1/m1_n130_1870# 8.59886f
C436 end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272133f
C437 mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C438 end_1/8_cap_array_final_1/m1_n130_2110# end_1/8_cap_array_final_1/m1_n130_1990# 8.59886f
C439 end_0/8_cap_array_final_1/m1_n130_2230# end_0/8_cap_array_final_1/m1_n130_2110# 8.59886f
C440 mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C441 gnd phi2_n4 3.442492f
C442 mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C443 mid_6to8_3/8_cap_array_final_1/m1_n130_2110# mid_6to8_3/8_cap_array_final_1/m1_n130_1990# 8.59886f
C444 phi15 phi14 84.24828f
C445 end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002493f
C446 mid_4to8_0/8_cap_array_final_1/m1_n130_1750# mid_4to8_0/8_cap_array_final_1/m1_n130_1630# 8.59886f
C447 mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C448 phi17 vin 6.758001f
C449 phi1_n4 phi1_n6 42.41612f
C450 end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C451 phi2_n2 phi1_n3 24.224823f
C452 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# 5.002839f
C453 end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002494f
C454 end_3/8_cap_array_final_1/m1_n130_4340# end_3/8_cap_array_final_1/m1_n130_4460# 8.59886f
C455 mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C456 end_3/8_cap_array_final_1/m1_n130_3860# phi2_n7 8.726839f
C457 mid_4to8_2/8_cap_array_final_1/m1_n130_4220# phi2_n5 8.649531f
C458 end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002494f
C459 gnd phi26 2.737761f
C460 mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C461 mid_6to8_2/8_cap_array_final_1/m1_n130_4460# mid_6to8_2/8_cap_array_final_1/m1_n130_4340# 8.59886f
C462 phi16 phi25 39.08674f
C463 end_3/8_cap_array_final_1/m1_n130_3980# end_3/8_cap_array_final_1/m1_n130_3860# 8.59886f
C464 end_3/8_cap_array_final_1/m1_n130_4220# end_3/8_cap_array_final_1/m1_n130_4100# 8.59886f
C465 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# 5.002839f
C466 phi2_n6 phi2_n4 36.33864f
C467 end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002494f
C468 end_3/8_cap_array_final_1/m1_n130_1870# end_3/8_cap_array_final_1/m1_n130_1750# 8.59886f
C469 mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C470 phi15 phi1_n5 3.571209f
C471 mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C472 phi26 phi25 36.94984f
C473 mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C474 phi1_n7 phi1_n5 2.907911f
C475 end_1/8_cap_array_final_1/m1_n130_1990# end_1/8_cap_array_final_1/m1_n130_1870# 8.59886f
C476 end_0/8_cap_array_final_1/m1_n130_2110# end_0/8_cap_array_final_1/m1_n130_1990# 8.59886f
C477 phi2_n3 mid_2to4__1/8_cap_array_final_1/m1_n130_4460# 8.620945f
C478 end_0/8_cap_array_final_1/m1_n130_4340# end_0/8_cap_array_final_1/m1_n130_4220# 8.59886f
C479 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# 5.002838f
C480 mid_6to8_0/8_cap_array_final_1/m1_n130_4340# mid_6to8_0/8_cap_array_final_1/m1_n130_4220# 8.59886f
C481 mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272134f
C482 mid_6to8_3/8_cap_array_final_1/m1_n130_1990# mid_6to8_3/8_cap_array_final_1/m1_n130_1870# 8.59886f
C483 phi1_n7 vin 46.440384f
C484 phi1_n0 phi1_n3 9.193998f
C485 end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C486 mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C487 smpl_n_d12_out_n mid_2_0/8_cap_array_final_0/cap_final_0/phi1_n 25.579062f
C488 mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C489 phi1_n4 phi2_n5 6.385192f
C490 phi11 phi10 8.931144f
C491 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# 5.002838f
C492 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# 5.002839f
C493 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# 5.002838f
C494 mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C495 phi2_n6 phi26 4.41222f
C496 mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C497 mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C498 end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C499 phi1_n6 Vdd 18.423512f
C500 end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C501 mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C502 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# 5.002839f
C503 end_0/8_cap_array_final_1/m1_n130_4460# end_0/8_cap_array_final_1/m1_n130_4340# 8.59886f
C504 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# 4.980177f
C505 phi15 phi24 43.602276f
C506 mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C507 phi2_n4 phi1_n2 2.193301f
C508 end_3/8_cap_array_final_1/m1_n130_1750# end_3/8_cap_array_final_1/m1_n130_1630# 8.59886f
C509 end_2/8_cap_array_final_1/m1_n130_2230# phi27 8.728627f
C510 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# 5.002839f
C511 mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C512 mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C513 mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C514 end_1/8_cap_array_final_1/m1_n130_1870# end_1/8_cap_array_final_1/m1_n130_1750# 8.59886f
C515 end_0/8_cap_array_final_1/m1_n130_1990# end_0/8_cap_array_final_1/m1_n130_1870# 8.59886f
C516 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# 5.002493f
C517 phi1_n0 smpl_n_d12_out_n 21.9671f
C518 smpl_n_d12 SUB 2.977575f
C519 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C520 mid_2_0/mid_2_low_0/m4_2410_n9430# SUB 3.134649f **FLOATING
C521 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.34045f **FLOATING
C522 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.34039f **FLOATING
C523 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.340337f **FLOATING
C524 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340289f **FLOATING
C525 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.33782f **FLOATING
C526 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.340238f **FLOATING
C527 phi2_n1 SUB 18.851517f
C528 mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C529 mid_2_0/m4_2410_n9430# SUB 3.134649f **FLOATING
C530 mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.34045f **FLOATING
C531 mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.34039f **FLOATING
C532 mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.340337f **FLOATING
C533 mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340289f **FLOATING
C534 mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.33782f **FLOATING
C535 mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.340237f **FLOATING
C536 smpl SUB 6.026207f
C537 mid_2_0/8_cap_array_final_0/cap_final_0/phi1_n SUB 6.313595f
C538 smpl_n_d12_out_n SUB 10.418909f
C539 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340289f **FLOATING
C540 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.340337f **FLOATING
C541 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.340391f **FLOATING
C542 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.34045f **FLOATING
C543 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.34045f **FLOATING
C544 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C545 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.340247f **FLOATING
C546 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.475443f **FLOATING
C547 phi21 SUB 6.518417f
C548 phi23 SUB 10.791802f
C549 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340289f **FLOATING
C550 phi13 SUB 13.502681f
C551 phi1_n3 SUB 17.066725f
C552 phi2_n3 SUB 17.588808f
C553 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.340337f **FLOATING
C554 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.340391f **FLOATING
C555 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.34045f **FLOATING
C556 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.34045f **FLOATING
C557 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C558 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.340247f **FLOATING
C559 phi11 SUB 10.145213f
C560 phi1_n1 SUB 14.422091f
C561 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.475442f **FLOATING
C562 mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C563 mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.340515f **FLOATING
C564 mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.340515f **FLOATING
C565 mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.34045f **FLOATING
C566 mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.34045f **FLOATING
C567 mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.34045f **FLOATING
C568 mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.337859f **FLOATING
C569 mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.34045f **FLOATING
C570 mid_6to8_3/8_cap_array_final_1/m1_n130_1630# SUB 6.903774f
C571 mid_6to8_3/8_cap_array_final_1/m1_n130_1750# SUB 2.161829f
C572 mid_6to8_3/8_cap_array_final_1/m1_n130_1870# SUB 2.166234f
C573 mid_6to8_3/8_cap_array_final_1/m1_n130_1990# SUB 2.174879f
C574 mid_6to8_3/8_cap_array_final_1/m1_n130_2110# SUB 2.193039f
C575 mid_6to8_3/8_cap_array_final_1/m1_n130_3980# SUB 2.15064f
C576 mid_6to8_3/8_cap_array_final_1/m1_n130_4100# SUB 2.15295f
C577 mid_6to8_3/8_cap_array_final_1/m1_n130_4220# SUB 2.15295f
C578 mid_6to8_3/8_cap_array_final_1/m1_n130_4340# SUB 2.15295f
C579 mid_6to8_3/8_cap_array_final_1/m1_n130_4460# SUB 6.89743f
C580 mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.34045f **FLOATING
C581 mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# SUB 3.34045f **FLOATING
C582 mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.34045f **FLOATING
C583 mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.340515f **FLOATING
C584 mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.340515f **FLOATING
C585 mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C586 mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.34045f **FLOATING
C587 mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.47539f **FLOATING
C588 end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C589 end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.340515f **FLOATING
C590 end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.340515f **FLOATING
C591 end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.340515f **FLOATING
C592 end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.340515f **FLOATING
C593 end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C594 end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.337859f **FLOATING
C595 end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.340514f **FLOATING
C596 end_3/8_cap_array_final_1/m1_n130_1630# SUB 6.903774f
C597 end_3/8_cap_array_final_1/m1_n130_1750# SUB 2.161829f
C598 end_3/8_cap_array_final_1/m1_n130_1870# SUB 2.166234f
C599 end_3/8_cap_array_final_1/m1_n130_1990# SUB 2.174879f
C600 end_3/8_cap_array_final_1/m1_n130_2110# SUB 2.195349f
C601 end_3/8_cap_array_final_1/m1_n130_2230# SUB 3.840402f
C602 end_3/8_cap_array_final_1/m1_n130_3860# SUB 3.732141f
C603 end_3/8_cap_array_final_1/m1_n130_3980# SUB 2.15295f
C604 end_3/8_cap_array_final_1/m1_n130_4100# SUB 2.15295f
C605 end_3/8_cap_array_final_1/m1_n130_4220# SUB 2.15295f
C606 end_3/8_cap_array_final_1/m1_n130_4340# SUB 2.15295f
C607 end_3/8_cap_array_final_1/m1_n130_4460# SUB 6.89743f
C608 end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C609 end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# SUB 3.340515f **FLOATING
C610 end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.340515f **FLOATING
C611 end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.340515f **FLOATING
C612 end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.340515f **FLOATING
C613 end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C614 end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.340514f **FLOATING
C615 end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.47539f **FLOATING
C616 mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C617 mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.340515f **FLOATING
C618 mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.340515f **FLOATING
C619 mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.34045f **FLOATING
C620 mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.34045f **FLOATING
C621 mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.34045f **FLOATING
C622 mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.337859f **FLOATING
C623 mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.34045f **FLOATING
C624 mid_6to8_2/8_cap_array_final_1/m1_n130_1630# SUB 6.903774f
C625 mid_6to8_2/8_cap_array_final_1/m1_n130_1750# SUB 2.161829f
C626 mid_6to8_2/8_cap_array_final_1/m1_n130_1870# SUB 2.166234f
C627 mid_6to8_2/8_cap_array_final_1/m1_n130_1990# SUB 2.174879f
C628 mid_6to8_2/8_cap_array_final_1/m1_n130_2110# SUB 2.193039f
C629 mid_6to8_2/8_cap_array_final_1/m1_n130_3980# SUB 2.15064f
C630 mid_6to8_2/8_cap_array_final_1/m1_n130_4100# SUB 2.15295f
C631 mid_6to8_2/8_cap_array_final_1/m1_n130_4220# SUB 2.15295f
C632 mid_6to8_2/8_cap_array_final_1/m1_n130_4340# SUB 2.15295f
C633 mid_6to8_2/8_cap_array_final_1/m1_n130_4460# SUB 6.89743f
C634 mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.34045f **FLOATING
C635 mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# SUB 3.34045f **FLOATING
C636 mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.34045f **FLOATING
C637 mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.340515f **FLOATING
C638 mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.340515f **FLOATING
C639 mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C640 mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.34045f **FLOATING
C641 mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.47539f **FLOATING
C642 end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C643 end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.340515f **FLOATING
C644 end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.340515f **FLOATING
C645 end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.340515f **FLOATING
C646 end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.340515f **FLOATING
C647 end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C648 end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.337859f **FLOATING
C649 end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.340514f **FLOATING
C650 end_2/8_cap_array_final_1/m1_n130_1630# SUB 6.903774f
C651 end_2/8_cap_array_final_1/m1_n130_1750# SUB 2.161829f
C652 end_2/8_cap_array_final_1/m1_n130_1870# SUB 2.166234f
C653 end_2/8_cap_array_final_1/m1_n130_1990# SUB 2.174879f
C654 end_2/8_cap_array_final_1/m1_n130_2110# SUB 2.195349f
C655 end_2/8_cap_array_final_1/m1_n130_2230# SUB 3.840402f
C656 end_2/8_cap_array_final_1/m1_n130_3860# SUB 3.732141f
C657 end_2/8_cap_array_final_1/m1_n130_3980# SUB 2.15295f
C658 end_2/8_cap_array_final_1/m1_n130_4100# SUB 2.15295f
C659 end_2/8_cap_array_final_1/m1_n130_4220# SUB 2.15295f
C660 end_2/8_cap_array_final_1/m1_n130_4340# SUB 2.15295f
C661 end_2/8_cap_array_final_1/m1_n130_4460# SUB 6.89743f
C662 end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C663 end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# SUB 3.340515f **FLOATING
C664 end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.340515f **FLOATING
C665 end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.340515f **FLOATING
C666 end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.340515f **FLOATING
C667 end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C668 end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.340514f **FLOATING
C669 end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.47539f **FLOATING
C670 end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C671 end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.340515f **FLOATING
C672 end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.340515f **FLOATING
C673 end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.340515f **FLOATING
C674 end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.340515f **FLOATING
C675 end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C676 end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.337859f **FLOATING
C677 end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.340514f **FLOATING
C678 end_1/8_cap_array_final_1/m1_n130_1630# SUB 6.903774f
C679 end_1/8_cap_array_final_1/m1_n130_1750# SUB 2.161829f
C680 end_1/8_cap_array_final_1/m1_n130_1870# SUB 2.166234f
C681 end_1/8_cap_array_final_1/m1_n130_1990# SUB 2.174879f
C682 end_1/8_cap_array_final_1/m1_n130_2110# SUB 2.195349f
C683 end_1/8_cap_array_final_1/m1_n130_2230# SUB 3.840402f
C684 end_1/8_cap_array_final_1/m1_n130_3860# SUB 3.732141f
C685 end_1/8_cap_array_final_1/m1_n130_3980# SUB 2.15295f
C686 end_1/8_cap_array_final_1/m1_n130_4100# SUB 2.15295f
C687 end_1/8_cap_array_final_1/m1_n130_4220# SUB 2.15295f
C688 end_1/8_cap_array_final_1/m1_n130_4340# SUB 2.15295f
C689 end_1/8_cap_array_final_1/m1_n130_4460# SUB 6.89743f
C690 end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C691 end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# SUB 3.340515f **FLOATING
C692 end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.340515f **FLOATING
C693 end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.340515f **FLOATING
C694 end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.340515f **FLOATING
C695 end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C696 end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.340514f **FLOATING
C697 end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.47539f **FLOATING
C698 mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C699 mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.340515f **FLOATING
C700 mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.340515f **FLOATING
C701 mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.34045f **FLOATING
C702 mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.34045f **FLOATING
C703 mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.34045f **FLOATING
C704 mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.337859f **FLOATING
C705 mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.34045f **FLOATING
C706 mid_6to8_1/8_cap_array_final_1/m1_n130_1630# SUB 6.903774f
C707 mid_6to8_1/8_cap_array_final_1/m1_n130_1750# SUB 2.161829f
C708 mid_6to8_1/8_cap_array_final_1/m1_n130_1870# SUB 2.166234f
C709 mid_6to8_1/8_cap_array_final_1/m1_n130_1990# SUB 2.174879f
C710 mid_6to8_1/8_cap_array_final_1/m1_n130_2110# SUB 2.193039f
C711 mid_6to8_1/8_cap_array_final_1/m1_n130_3980# SUB 2.15064f
C712 mid_6to8_1/8_cap_array_final_1/m1_n130_4100# SUB 2.15295f
C713 mid_6to8_1/8_cap_array_final_1/m1_n130_4220# SUB 2.15295f
C714 mid_6to8_1/8_cap_array_final_1/m1_n130_4340# SUB 2.15295f
C715 mid_6to8_1/8_cap_array_final_1/m1_n130_4460# SUB 6.89743f
C716 mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.34045f **FLOATING
C717 mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# SUB 3.34045f **FLOATING
C718 mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.34045f **FLOATING
C719 mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.340515f **FLOATING
C720 mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.340515f **FLOATING
C721 mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C722 mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.34045f **FLOATING
C723 mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.47539f **FLOATING
C724 end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C725 end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.340515f **FLOATING
C726 end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.340515f **FLOATING
C727 end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.340515f **FLOATING
C728 end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.340515f **FLOATING
C729 end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C730 end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.337859f **FLOATING
C731 end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.340514f **FLOATING
C732 end_0/8_cap_array_final_1/m1_n130_1630# SUB 6.903774f
C733 end_0/8_cap_array_final_1/m1_n130_1750# SUB 2.161829f
C734 end_0/8_cap_array_final_1/m1_n130_1870# SUB 2.166234f
C735 end_0/8_cap_array_final_1/m1_n130_1990# SUB 2.174879f
C736 end_0/8_cap_array_final_1/m1_n130_2110# SUB 2.195349f
C737 end_0/8_cap_array_final_1/m1_n130_2230# SUB 3.840402f
C738 end_0/8_cap_array_final_1/m1_n130_3860# SUB 3.732141f
C739 end_0/8_cap_array_final_1/m1_n130_3980# SUB 2.15295f
C740 end_0/8_cap_array_final_1/m1_n130_4100# SUB 2.15295f
C741 end_0/8_cap_array_final_1/m1_n130_4220# SUB 2.15295f
C742 end_0/8_cap_array_final_1/m1_n130_4340# SUB 2.15295f
C743 end_0/8_cap_array_final_1/m1_n130_4460# SUB 6.89743f
C744 end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C745 end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# SUB 3.340515f **FLOATING
C746 end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.340515f **FLOATING
C747 end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.340515f **FLOATING
C748 end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.340515f **FLOATING
C749 phi27 SUB 0.349636p
C750 phi2_n7 SUB 68.62492f
C751 end_3/8_cap_array_final_1/cap_final_7/com_x SUB 0.124406p
C752 end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C753 vin SUB 0.115031p
C754 Vdd SUB 0.491736p
C755 gnd SUB 0.125852p
C756 end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.340514f **FLOATING
C757 end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.475423f **FLOATING
C758 phi17 SUB 0.137742p
C759 phi1_n7 SUB 95.30315f
C760 mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C761 mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.340515f **FLOATING
C762 mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.340515f **FLOATING
C763 mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.34045f **FLOATING
C764 mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.34045f **FLOATING
C765 mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.34045f **FLOATING
C766 mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.337859f **FLOATING
C767 mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.34045f **FLOATING
C768 mid_6to8_0/8_cap_array_final_1/m1_n130_1630# SUB 6.903774f
C769 mid_6to8_0/8_cap_array_final_1/m1_n130_1750# SUB 2.161829f
C770 mid_6to8_0/8_cap_array_final_1/m1_n130_1870# SUB 2.166234f
C771 mid_6to8_0/8_cap_array_final_1/m1_n130_1990# SUB 2.174879f
C772 mid_6to8_0/8_cap_array_final_1/m1_n130_2110# SUB 2.193039f
C773 phi2_n6 SUB 60.42595f
C774 mid_6to8_0/8_cap_array_final_1/m1_n130_3980# SUB 2.15064f
C775 mid_6to8_0/8_cap_array_final_1/m1_n130_4100# SUB 2.15295f
C776 mid_6to8_0/8_cap_array_final_1/m1_n130_4220# SUB 2.15295f
C777 mid_6to8_0/8_cap_array_final_1/m1_n130_4340# SUB 2.15295f
C778 mid_6to8_0/8_cap_array_final_1/m1_n130_4460# SUB 6.89743f
C779 mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.34045f **FLOATING
C780 mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# SUB 3.34045f **FLOATING
C781 mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.34045f **FLOATING
C782 phi16 SUB 60.440945f
C783 phi1_n6 SUB 53.428093f
C784 phi26 SUB 75.38205f
C785 mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.340515f **FLOATING
C786 mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.340515f **FLOATING
C787 mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C788 mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.34045f **FLOATING
C789 mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.47539f **FLOATING
C790 mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C791 mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.34045f **FLOATING
C792 mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.34045f **FLOATING
C793 mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.34039f **FLOATING
C794 mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.340337f **FLOATING
C795 mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.340289f **FLOATING
C796 mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.337859f **FLOATING
C797 mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.340247f **FLOATING
C798 mid_2to4__1/8_cap_array_final_1/m1_n130_1630# SUB 6.902235f
C799 mid_2to4__1/8_cap_array_final_1/m1_n130_4460# SUB 6.89589f
C800 mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.340289f **FLOATING
C801 mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# SUB 3.340337f **FLOATING
C802 mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.34039f **FLOATING
C803 mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.34045f **FLOATING
C804 mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.34045f **FLOATING
C805 mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C806 mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.340247f **FLOATING
C807 mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.47539f **FLOATING
C808 phi22 SUB 6.805904f
C809 mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C810 mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.34045f **FLOATING
C811 mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.34045f **FLOATING
C812 mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.34039f **FLOATING
C813 mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.340337f **FLOATING
C814 mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.340289f **FLOATING
C815 mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.337859f **FLOATING
C816 mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.340247f **FLOATING
C817 mid_2to4__0/8_cap_array_final_1/m1_n130_1630# SUB 6.902235f
C818 mid_2to4__0/8_cap_array_final_1/m1_n130_4460# SUB 6.89589f
C819 mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.340289f **FLOATING
C820 phi12 SUB 6.635001f
C821 phi1_n2 SUB 10.978977f
C822 phi2_n2 SUB 10.279954f
C823 mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# SUB 3.340337f **FLOATING
C824 mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.34039f **FLOATING
C825 mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.34045f **FLOATING
C826 mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.34045f **FLOATING
C827 mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C828 mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.340247f **FLOATING
C829 mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.47539f **FLOATING
C830 mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C831 mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.34045f **FLOATING
C832 mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.34045f **FLOATING
C833 mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.34039f **FLOATING
C834 mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.340337f **FLOATING
C835 mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.340337f **FLOATING
C836 mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.337859f **FLOATING
C837 mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.340337f **FLOATING
C838 mid_4to8_3/8_cap_array_final_1/m1_n130_1630# SUB 6.903774f
C839 mid_4to8_3/8_cap_array_final_1/m1_n130_1750# SUB 2.161829f
C840 mid_4to8_3/8_cap_array_final_1/m1_n130_1870# SUB 2.163925f
C841 mid_4to8_3/8_cap_array_final_1/m1_n130_4220# SUB 2.15064f
C842 mid_4to8_3/8_cap_array_final_1/m1_n130_4340# SUB 2.15295f
C843 mid_4to8_3/8_cap_array_final_1/m1_n130_4460# SUB 6.89743f
C844 mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.340337f **FLOATING
C845 mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# SUB 3.340337f **FLOATING
C846 mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.34039f **FLOATING
C847 mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.34045f **FLOATING
C848 mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.34045f **FLOATING
C849 mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C850 mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.340337f **FLOATING
C851 mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.47539f **FLOATING
C852 mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C853 mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.34045f **FLOATING
C854 mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.34045f **FLOATING
C855 mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.34039f **FLOATING
C856 mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.340337f **FLOATING
C857 mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.340337f **FLOATING
C858 mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.337859f **FLOATING
C859 mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.340337f **FLOATING
C860 mid_4to8_2/8_cap_array_final_1/m1_n130_1630# SUB 6.903774f
C861 mid_4to8_2/8_cap_array_final_1/m1_n130_1750# SUB 2.161829f
C862 mid_4to8_2/8_cap_array_final_1/m1_n130_1870# SUB 2.163925f
C863 mid_4to8_2/8_cap_array_final_1/m1_n130_4220# SUB 2.15064f
C864 mid_4to8_2/8_cap_array_final_1/m1_n130_4340# SUB 2.15295f
C865 mid_4to8_2/8_cap_array_final_1/m1_n130_4460# SUB 6.89743f
C866 mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.340337f **FLOATING
C867 mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# SUB 3.340337f **FLOATING
C868 mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.34039f **FLOATING
C869 mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.34045f **FLOATING
C870 mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.34045f **FLOATING
C871 mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C872 mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.340337f **FLOATING
C873 mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.47539f **FLOATING
C874 mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C875 mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.34045f **FLOATING
C876 mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.34045f **FLOATING
C877 mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.34039f **FLOATING
C878 mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.340337f **FLOATING
C879 mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.340337f **FLOATING
C880 mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.337859f **FLOATING
C881 mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.340337f **FLOATING
C882 mid_4to8_1/8_cap_array_final_1/m1_n130_1630# SUB 6.903774f
C883 mid_4to8_1/8_cap_array_final_1/m1_n130_1750# SUB 2.161829f
C884 mid_4to8_1/8_cap_array_final_1/m1_n130_1870# SUB 2.163925f
C885 mid_4to8_1/8_cap_array_final_1/m1_n130_4220# SUB 2.15064f
C886 mid_4to8_1/8_cap_array_final_1/m1_n130_4340# SUB 2.15295f
C887 mid_4to8_1/8_cap_array_final_1/m1_n130_4460# SUB 6.89743f
C888 mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.340337f **FLOATING
C889 mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# SUB 3.340337f **FLOATING
C890 mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.34039f **FLOATING
C891 mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.34045f **FLOATING
C892 mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.34045f **FLOATING
C893 mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C894 mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.340337f **FLOATING
C895 mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.47539f **FLOATING
C896 phi25 SUB 34.537025f
C897 phi2_n4 SUB 23.24144f
C898 phi2_n5 SUB 28.663544f
C899 mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# SUB 3.340515f **FLOATING
C900 mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# SUB 3.34045f **FLOATING
C901 mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# SUB 3.34045f **FLOATING
C902 mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# SUB 3.34039f **FLOATING
C903 mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# SUB 3.340337f **FLOATING
C904 mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# SUB 3.340337f **FLOATING
C905 mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# SUB 3.337859f **FLOATING
C906 mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# SUB 3.340337f **FLOATING
C907 mid_4to8_0/8_cap_array_final_1/m1_n130_1630# SUB 6.903774f
C908 mid_4to8_0/8_cap_array_final_1/m1_n130_1750# SUB 2.161829f
C909 mid_4to8_0/8_cap_array_final_1/m1_n130_1870# SUB 2.163925f
C910 phi24 SUB 22.777933f
C911 mid_4to8_0/8_cap_array_final_1/m1_n130_4220# SUB 2.15064f
C912 mid_4to8_0/8_cap_array_final_1/m1_n130_4340# SUB 2.15295f
C913 mid_4to8_0/8_cap_array_final_1/m1_n130_4460# SUB 6.89743f
C914 mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# SUB 3.340337f **FLOATING
C915 mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# SUB 3.340337f **FLOATING
C916 phi15 SUB 33.756042f
C917 phi1_n5 SUB 34.770325f
C918 mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# SUB 3.34039f **FLOATING
C919 phi14 SUB 20.096615f
C920 phi1_n4 SUB 22.603916f
C921 mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# SUB 3.34045f **FLOATING
C922 mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# SUB 3.34045f **FLOATING
C923 mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# SUB 3.340515f **FLOATING
C924 mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# SUB 3.340337f **FLOATING
C925 mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# SUB 3.47539f **FLOATING
