magic
tech sky130A
magscale 1 2
timestamp 1730037944
<< error_s >>
rect 3832 28420 3872 28438
rect 3860 28392 3900 28410
<< nwell >>
rect 3310 65820 3878 66552
rect 8300 65820 8868 66552
rect 13290 65820 13858 66552
rect 18280 65820 18848 66552
rect 23270 65820 23838 66552
rect 28260 65820 28828 66552
rect 33250 65820 33818 66552
rect 38240 65820 38808 66552
rect 43230 65820 43798 66552
rect 48220 65820 48788 66552
rect 53210 65820 53778 66552
rect 58200 65820 58768 66552
rect 63190 65820 63758 66552
rect 68180 65820 68748 66552
rect 73170 65820 73738 66552
rect 78160 65820 78728 66552
rect 3310 64110 3878 64842
rect 8300 64110 8868 64842
rect 13290 64110 13858 64842
rect 18280 64110 18848 64842
rect 23270 64110 23838 64842
rect 28260 64110 28828 64842
rect 33250 64110 33818 64842
rect 38240 64110 38808 64842
rect 43230 64110 43798 64842
rect 48220 64110 48788 64842
rect 53210 64110 53778 64842
rect 58200 64110 58768 64842
rect 63190 64110 63758 64842
rect 68180 64110 68748 64842
rect 73170 64110 73738 64842
rect 78160 64110 78728 64842
rect 3310 62400 3878 63132
rect 8300 62400 8868 63132
rect 13290 62400 13858 63132
rect 18280 62400 18848 63132
rect 23270 62400 23838 63132
rect 28260 62400 28828 63132
rect 33250 62400 33818 63132
rect 38240 62400 38808 63132
rect 43230 62400 43798 63132
rect 48220 62400 48788 63132
rect 53210 62400 53778 63132
rect 58200 62400 58768 63132
rect 63190 62400 63758 63132
rect 68180 62400 68748 63132
rect 73170 62400 73738 63132
rect 78160 62400 78728 63132
rect 3310 60690 3878 61422
rect 8300 60690 8868 61422
rect 13290 60690 13858 61422
rect 18280 60690 18848 61422
rect 23270 60690 23838 61422
rect 28260 60690 28828 61422
rect 33250 60690 33818 61422
rect 38240 60690 38808 61422
rect 43230 60690 43798 61422
rect 48220 60690 48788 61422
rect 53210 60690 53778 61422
rect 58200 60690 58768 61422
rect 63190 60690 63758 61422
rect 68180 60690 68748 61422
rect 73170 60690 73738 61422
rect 78160 60690 78728 61422
rect 3310 58980 3878 59712
rect 8300 58980 8868 59712
rect 13290 58980 13858 59712
rect 18280 58980 18848 59712
rect 23270 58980 23838 59712
rect 28260 58980 28828 59712
rect 33250 58980 33818 59712
rect 38240 58980 38808 59712
rect 43230 58980 43798 59712
rect 48220 58980 48788 59712
rect 53210 58980 53778 59712
rect 58200 58980 58768 59712
rect 63190 58980 63758 59712
rect 68180 58980 68748 59712
rect 73170 58980 73738 59712
rect 78160 58980 78728 59712
rect 3310 57270 3878 58002
rect 8300 57270 8868 58002
rect 13290 57270 13858 58002
rect 18280 57270 18848 58002
rect 23270 57270 23838 58002
rect 28260 57270 28828 58002
rect 33250 57270 33818 58002
rect 38240 57270 38808 58002
rect 43230 57270 43798 58002
rect 48220 57270 48788 58002
rect 53210 57270 53778 58002
rect 58200 57270 58768 58002
rect 63190 57270 63758 58002
rect 68180 57270 68748 58002
rect 73170 57270 73738 58002
rect 78160 57270 78728 58002
rect 3310 55560 3878 56292
rect 8300 55560 8868 56292
rect 13290 55560 13858 56292
rect 18280 55560 18848 56292
rect 23270 55560 23838 56292
rect 28260 55560 28828 56292
rect 33250 55560 33818 56292
rect 38240 55560 38808 56292
rect 43230 55560 43798 56292
rect 48220 55560 48788 56292
rect 53210 55560 53778 56292
rect 58200 55560 58768 56292
rect 63190 55560 63758 56292
rect 68180 55560 68748 56292
rect 73170 55560 73738 56292
rect 78160 55560 78728 56292
rect 3310 53850 3878 54582
rect 8300 53850 8868 54582
rect 13290 53850 13858 54582
rect 18280 53850 18848 54582
rect 23270 53850 23838 54582
rect 28260 53850 28828 54582
rect 33250 53850 33818 54582
rect 38240 53850 38808 54582
rect 43230 53850 43798 54582
rect 48220 53850 48788 54582
rect 53210 53850 53778 54582
rect 58200 53850 58768 54582
rect 63190 53850 63758 54582
rect 68180 53850 68748 54582
rect 73170 53850 73738 54582
rect 78160 53850 78728 54582
rect 3310 52140 3878 52872
rect 8300 52140 8868 52872
rect 13290 52140 13858 52872
rect 18280 52140 18848 52872
rect 23270 52140 23838 52872
rect 28260 52140 28828 52872
rect 33250 52140 33818 52872
rect 38240 52140 38808 52872
rect 43230 52140 43798 52872
rect 48220 52140 48788 52872
rect 53210 52140 53778 52872
rect 58200 52140 58768 52872
rect 63190 52140 63758 52872
rect 68180 52140 68748 52872
rect 73170 52140 73738 52872
rect 78160 52140 78728 52872
rect 3310 50430 3878 51162
rect 8300 50430 8868 51162
rect 13290 50430 13858 51162
rect 18280 50430 18848 51162
rect 23270 50430 23838 51162
rect 28260 50430 28828 51162
rect 33250 50430 33818 51162
rect 38240 50430 38808 51162
rect 43230 50430 43798 51162
rect 48220 50430 48788 51162
rect 53210 50430 53778 51162
rect 58200 50430 58768 51162
rect 63190 50430 63758 51162
rect 68180 50430 68748 51162
rect 73170 50430 73738 51162
rect 78160 50430 78728 51162
rect 3310 48720 3878 49452
rect 8300 48720 8868 49452
rect 13290 48720 13858 49452
rect 18280 48720 18848 49452
rect 23270 48720 23838 49452
rect 28260 48720 28828 49452
rect 33250 48720 33818 49452
rect 38240 48720 38808 49452
rect 43230 48720 43798 49452
rect 48220 48720 48788 49452
rect 53210 48720 53778 49452
rect 58200 48720 58768 49452
rect 63190 48720 63758 49452
rect 68180 48720 68748 49452
rect 73170 48720 73738 49452
rect 78160 48720 78728 49452
rect 3310 47010 3878 47742
rect 8300 47010 8868 47742
rect 13290 47010 13858 47742
rect 18280 47010 18848 47742
rect 23270 47010 23838 47742
rect 28260 47010 28828 47742
rect 33250 47010 33818 47742
rect 38240 47010 38808 47742
rect 43230 47010 43798 47742
rect 48220 47010 48788 47742
rect 53210 47010 53778 47742
rect 58200 47010 58768 47742
rect 63190 47010 63758 47742
rect 68180 47010 68748 47742
rect 73170 47010 73738 47742
rect 78160 47010 78728 47742
rect 3310 45300 3878 46032
rect 8300 45300 8868 46032
rect 13290 45300 13858 46032
rect 18280 45300 18848 46032
rect 23270 45300 23838 46032
rect 28260 45300 28828 46032
rect 33250 45300 33818 46032
rect 38240 45300 38808 46032
rect 43230 45300 43798 46032
rect 48220 45300 48788 46032
rect 53210 45300 53778 46032
rect 58200 45300 58768 46032
rect 63190 45300 63758 46032
rect 68180 45300 68748 46032
rect 73170 45300 73738 46032
rect 78160 45300 78728 46032
rect 3310 43590 3878 44322
rect 8300 43590 8868 44322
rect 13290 43590 13858 44322
rect 18280 43590 18848 44322
rect 23270 43590 23838 44322
rect 28260 43590 28828 44322
rect 33250 43590 33818 44322
rect 38240 43590 38808 44322
rect 43230 43590 43798 44322
rect 48220 43590 48788 44322
rect 53210 43590 53778 44322
rect 58200 43590 58768 44322
rect 63190 43590 63758 44322
rect 68180 43590 68748 44322
rect 73170 43590 73738 44322
rect 78160 43590 78728 44322
rect 3310 41880 3878 42612
rect 8300 41880 8868 42612
rect 13290 41880 13858 42612
rect 18280 41880 18848 42612
rect 23270 41880 23838 42612
rect 28260 41880 28828 42612
rect 33250 41880 33818 42612
rect 38240 41880 38808 42612
rect 43230 41880 43798 42612
rect 48220 41880 48788 42612
rect 53210 41880 53778 42612
rect 58200 41880 58768 42612
rect 63190 41880 63758 42612
rect 68180 41880 68748 42612
rect 73170 41880 73738 42612
rect 78160 41880 78728 42612
rect 3310 40170 3878 40902
rect 8300 40170 8868 40902
rect 13290 40170 13858 40902
rect 18280 40170 18848 40902
rect 23270 40170 23838 40902
rect 28260 40170 28828 40902
rect 33250 40170 33818 40902
rect 38240 40170 38808 40902
rect 43230 40170 43798 40902
rect 48220 40170 48788 40902
rect 53210 40170 53778 40902
rect 58200 40170 58768 40902
rect 63190 40170 63758 40902
rect 68180 40170 68748 40902
rect 73170 40170 73738 40902
rect 78160 40170 78728 40902
<< pwell >>
rect 2740 66590 2810 67050
rect 7730 66590 7800 67050
rect 12720 66590 12790 67050
rect 17710 66590 17780 67050
rect 22700 66590 22770 67050
rect 27690 66590 27760 67050
rect 32680 66590 32750 67050
rect 37670 66590 37740 67050
rect 42660 66590 42730 67050
rect 47650 66590 47720 67050
rect 52640 66590 52710 67050
rect 57630 66590 57700 67050
rect 62620 66590 62690 67050
rect 67610 66590 67680 67050
rect 72600 66590 72670 67050
rect 77590 66590 77660 67050
rect 2750 65820 3308 66552
rect 7740 65820 8298 66552
rect 12730 65820 13288 66552
rect 17720 65820 18278 66552
rect 22710 65820 23268 66552
rect 27700 65820 28258 66552
rect 32690 65820 33248 66552
rect 37680 65820 38238 66552
rect 42670 65820 43228 66552
rect 47660 65820 48218 66552
rect 52650 65820 53208 66552
rect 57640 65820 58198 66552
rect 62630 65820 63188 66552
rect 67620 65820 68178 66552
rect 72610 65820 73168 66552
rect 77600 65820 78158 66552
rect 2740 64880 2810 65340
rect 7730 64880 7800 65340
rect 12720 64880 12790 65340
rect 17710 64880 17780 65340
rect 22700 64880 22770 65340
rect 27690 64880 27760 65340
rect 32680 64880 32750 65340
rect 37670 64880 37740 65340
rect 42660 64880 42730 65340
rect 47650 64880 47720 65340
rect 52640 64880 52710 65340
rect 57630 64880 57700 65340
rect 62620 64880 62690 65340
rect 67610 64880 67680 65340
rect 72600 64880 72670 65340
rect 77590 64880 77660 65340
rect 2750 64110 3308 64842
rect 7740 64110 8298 64842
rect 12730 64110 13288 64842
rect 17720 64110 18278 64842
rect 22710 64110 23268 64842
rect 27700 64110 28258 64842
rect 32690 64110 33248 64842
rect 37680 64110 38238 64842
rect 42670 64110 43228 64842
rect 47660 64110 48218 64842
rect 52650 64110 53208 64842
rect 57640 64110 58198 64842
rect 62630 64110 63188 64842
rect 67620 64110 68178 64842
rect 72610 64110 73168 64842
rect 77600 64110 78158 64842
rect 2740 63170 2810 63630
rect 7730 63170 7800 63630
rect 12720 63170 12790 63630
rect 17710 63170 17780 63630
rect 22700 63170 22770 63630
rect 27690 63170 27760 63630
rect 32680 63170 32750 63630
rect 37670 63170 37740 63630
rect 42660 63170 42730 63630
rect 47650 63170 47720 63630
rect 52640 63170 52710 63630
rect 57630 63170 57700 63630
rect 62620 63170 62690 63630
rect 67610 63170 67680 63630
rect 72600 63170 72670 63630
rect 77590 63170 77660 63630
rect 2750 62400 3308 63132
rect 7740 62400 8298 63132
rect 12730 62400 13288 63132
rect 17720 62400 18278 63132
rect 22710 62400 23268 63132
rect 27700 62400 28258 63132
rect 32690 62400 33248 63132
rect 37680 62400 38238 63132
rect 42670 62400 43228 63132
rect 47660 62400 48218 63132
rect 52650 62400 53208 63132
rect 57640 62400 58198 63132
rect 62630 62400 63188 63132
rect 67620 62400 68178 63132
rect 72610 62400 73168 63132
rect 77600 62400 78158 63132
rect 2740 61460 2810 61920
rect 7730 61460 7800 61920
rect 12720 61460 12790 61920
rect 17710 61460 17780 61920
rect 22700 61460 22770 61920
rect 27690 61460 27760 61920
rect 32680 61460 32750 61920
rect 37670 61460 37740 61920
rect 42660 61460 42730 61920
rect 47650 61460 47720 61920
rect 52640 61460 52710 61920
rect 57630 61460 57700 61920
rect 62620 61460 62690 61920
rect 67610 61460 67680 61920
rect 72600 61460 72670 61920
rect 77590 61460 77660 61920
rect 2750 60690 3308 61422
rect 7740 60690 8298 61422
rect 12730 60690 13288 61422
rect 17720 60690 18278 61422
rect 22710 60690 23268 61422
rect 27700 60690 28258 61422
rect 32690 60690 33248 61422
rect 37680 60690 38238 61422
rect 42670 60690 43228 61422
rect 47660 60690 48218 61422
rect 52650 60690 53208 61422
rect 57640 60690 58198 61422
rect 62630 60690 63188 61422
rect 67620 60690 68178 61422
rect 72610 60690 73168 61422
rect 77600 60690 78158 61422
rect 2740 59750 2810 60210
rect 7730 59750 7800 60210
rect 12720 59750 12790 60210
rect 17710 59750 17780 60210
rect 22700 59750 22770 60210
rect 27690 59750 27760 60210
rect 32680 59750 32750 60210
rect 37670 59750 37740 60210
rect 42660 59750 42730 60210
rect 47650 59750 47720 60210
rect 52640 59750 52710 60210
rect 57630 59750 57700 60210
rect 62620 59750 62690 60210
rect 67610 59750 67680 60210
rect 72600 59750 72670 60210
rect 77590 59750 77660 60210
rect 2750 58980 3308 59712
rect 7740 58980 8298 59712
rect 12730 58980 13288 59712
rect 17720 58980 18278 59712
rect 22710 58980 23268 59712
rect 27700 58980 28258 59712
rect 32690 58980 33248 59712
rect 37680 58980 38238 59712
rect 42670 58980 43228 59712
rect 47660 58980 48218 59712
rect 52650 58980 53208 59712
rect 57640 58980 58198 59712
rect 62630 58980 63188 59712
rect 67620 58980 68178 59712
rect 72610 58980 73168 59712
rect 77600 58980 78158 59712
rect 2740 58040 2810 58500
rect 7730 58040 7800 58500
rect 12720 58040 12790 58500
rect 17710 58040 17780 58500
rect 22700 58040 22770 58500
rect 27690 58040 27760 58500
rect 32680 58040 32750 58500
rect 37670 58040 37740 58500
rect 42660 58040 42730 58500
rect 47650 58040 47720 58500
rect 52640 58040 52710 58500
rect 57630 58040 57700 58500
rect 62620 58040 62690 58500
rect 67610 58040 67680 58500
rect 72600 58040 72670 58500
rect 77590 58040 77660 58500
rect 2750 57270 3308 58002
rect 7740 57270 8298 58002
rect 12730 57270 13288 58002
rect 17720 57270 18278 58002
rect 22710 57270 23268 58002
rect 27700 57270 28258 58002
rect 32690 57270 33248 58002
rect 37680 57270 38238 58002
rect 42670 57270 43228 58002
rect 47660 57270 48218 58002
rect 52650 57270 53208 58002
rect 57640 57270 58198 58002
rect 62630 57270 63188 58002
rect 67620 57270 68178 58002
rect 72610 57270 73168 58002
rect 77600 57270 78158 58002
rect 2740 56330 2810 56790
rect 7730 56330 7800 56790
rect 12720 56330 12790 56790
rect 17710 56330 17780 56790
rect 22700 56330 22770 56790
rect 27690 56330 27760 56790
rect 32680 56330 32750 56790
rect 37670 56330 37740 56790
rect 42660 56330 42730 56790
rect 47650 56330 47720 56790
rect 52640 56330 52710 56790
rect 57630 56330 57700 56790
rect 62620 56330 62690 56790
rect 67610 56330 67680 56790
rect 72600 56330 72670 56790
rect 77590 56330 77660 56790
rect 2750 55560 3308 56292
rect 7740 55560 8298 56292
rect 12730 55560 13288 56292
rect 17720 55560 18278 56292
rect 22710 55560 23268 56292
rect 27700 55560 28258 56292
rect 32690 55560 33248 56292
rect 37680 55560 38238 56292
rect 42670 55560 43228 56292
rect 47660 55560 48218 56292
rect 52650 55560 53208 56292
rect 57640 55560 58198 56292
rect 62630 55560 63188 56292
rect 67620 55560 68178 56292
rect 72610 55560 73168 56292
rect 77600 55560 78158 56292
rect 2740 54620 2810 55080
rect 7730 54620 7800 55080
rect 12720 54620 12790 55080
rect 17710 54620 17780 55080
rect 22700 54620 22770 55080
rect 27690 54620 27760 55080
rect 32680 54620 32750 55080
rect 37670 54620 37740 55080
rect 42660 54620 42730 55080
rect 47650 54620 47720 55080
rect 52640 54620 52710 55080
rect 57630 54620 57700 55080
rect 62620 54620 62690 55080
rect 67610 54620 67680 55080
rect 72600 54620 72670 55080
rect 77590 54620 77660 55080
rect 2750 53850 3308 54582
rect 7740 53850 8298 54582
rect 12730 53850 13288 54582
rect 17720 53850 18278 54582
rect 22710 53850 23268 54582
rect 27700 53850 28258 54582
rect 32690 53850 33248 54582
rect 37680 53850 38238 54582
rect 42670 53850 43228 54582
rect 47660 53850 48218 54582
rect 52650 53850 53208 54582
rect 57640 53850 58198 54582
rect 62630 53850 63188 54582
rect 67620 53850 68178 54582
rect 72610 53850 73168 54582
rect 77600 53850 78158 54582
rect 2740 52910 2810 53370
rect 7730 52910 7800 53370
rect 12720 52910 12790 53370
rect 17710 52910 17780 53370
rect 22700 52910 22770 53370
rect 27690 52910 27760 53370
rect 32680 52910 32750 53370
rect 37670 52910 37740 53370
rect 42660 52910 42730 53370
rect 47650 52910 47720 53370
rect 52640 52910 52710 53370
rect 57630 52910 57700 53370
rect 62620 52910 62690 53370
rect 67610 52910 67680 53370
rect 72600 52910 72670 53370
rect 77590 52910 77660 53370
rect 2750 52140 3308 52872
rect 7740 52140 8298 52872
rect 12730 52140 13288 52872
rect 17720 52140 18278 52872
rect 22710 52140 23268 52872
rect 27700 52140 28258 52872
rect 32690 52140 33248 52872
rect 37680 52140 38238 52872
rect 42670 52140 43228 52872
rect 47660 52140 48218 52872
rect 52650 52140 53208 52872
rect 57640 52140 58198 52872
rect 62630 52140 63188 52872
rect 67620 52140 68178 52872
rect 72610 52140 73168 52872
rect 77600 52140 78158 52872
rect 2740 51200 2810 51660
rect 7730 51200 7800 51660
rect 12720 51200 12790 51660
rect 17710 51200 17780 51660
rect 22700 51200 22770 51660
rect 27690 51200 27760 51660
rect 32680 51200 32750 51660
rect 37670 51200 37740 51660
rect 42660 51200 42730 51660
rect 47650 51200 47720 51660
rect 52640 51200 52710 51660
rect 57630 51200 57700 51660
rect 62620 51200 62690 51660
rect 67610 51200 67680 51660
rect 72600 51200 72670 51660
rect 77590 51200 77660 51660
rect 2750 50430 3308 51162
rect 7740 50430 8298 51162
rect 12730 50430 13288 51162
rect 17720 50430 18278 51162
rect 22710 50430 23268 51162
rect 27700 50430 28258 51162
rect 32690 50430 33248 51162
rect 37680 50430 38238 51162
rect 42670 50430 43228 51162
rect 47660 50430 48218 51162
rect 52650 50430 53208 51162
rect 57640 50430 58198 51162
rect 62630 50430 63188 51162
rect 67620 50430 68178 51162
rect 72610 50430 73168 51162
rect 77600 50430 78158 51162
rect 2740 49490 2810 49950
rect 7730 49490 7800 49950
rect 12720 49490 12790 49950
rect 17710 49490 17780 49950
rect 22700 49490 22770 49950
rect 27690 49490 27760 49950
rect 32680 49490 32750 49950
rect 37670 49490 37740 49950
rect 42660 49490 42730 49950
rect 47650 49490 47720 49950
rect 52640 49490 52710 49950
rect 57630 49490 57700 49950
rect 62620 49490 62690 49950
rect 67610 49490 67680 49950
rect 72600 49490 72670 49950
rect 77590 49490 77660 49950
rect 2750 48720 3308 49452
rect 7740 48720 8298 49452
rect 12730 48720 13288 49452
rect 17720 48720 18278 49452
rect 22710 48720 23268 49452
rect 27700 48720 28258 49452
rect 32690 48720 33248 49452
rect 37680 48720 38238 49452
rect 42670 48720 43228 49452
rect 47660 48720 48218 49452
rect 52650 48720 53208 49452
rect 57640 48720 58198 49452
rect 62630 48720 63188 49452
rect 67620 48720 68178 49452
rect 72610 48720 73168 49452
rect 77600 48720 78158 49452
rect 2740 47780 2810 48240
rect 7730 47780 7800 48240
rect 12720 47780 12790 48240
rect 17710 47780 17780 48240
rect 22700 47780 22770 48240
rect 27690 47780 27760 48240
rect 32680 47780 32750 48240
rect 37670 47780 37740 48240
rect 42660 47780 42730 48240
rect 47650 47780 47720 48240
rect 52640 47780 52710 48240
rect 57630 47780 57700 48240
rect 62620 47780 62690 48240
rect 67610 47780 67680 48240
rect 72600 47780 72670 48240
rect 77590 47780 77660 48240
rect 2750 47010 3308 47742
rect 7740 47010 8298 47742
rect 12730 47010 13288 47742
rect 17720 47010 18278 47742
rect 22710 47010 23268 47742
rect 27700 47010 28258 47742
rect 32690 47010 33248 47742
rect 37680 47010 38238 47742
rect 42670 47010 43228 47742
rect 47660 47010 48218 47742
rect 52650 47010 53208 47742
rect 57640 47010 58198 47742
rect 62630 47010 63188 47742
rect 67620 47010 68178 47742
rect 72610 47010 73168 47742
rect 77600 47010 78158 47742
rect 2740 46070 2810 46530
rect 7730 46070 7800 46530
rect 12720 46070 12790 46530
rect 17710 46070 17780 46530
rect 22700 46070 22770 46530
rect 27690 46070 27760 46530
rect 32680 46070 32750 46530
rect 37670 46070 37740 46530
rect 42660 46070 42730 46530
rect 47650 46070 47720 46530
rect 52640 46070 52710 46530
rect 57630 46070 57700 46530
rect 62620 46070 62690 46530
rect 67610 46070 67680 46530
rect 72600 46070 72670 46530
rect 77590 46070 77660 46530
rect 2750 45300 3308 46032
rect 7740 45300 8298 46032
rect 12730 45300 13288 46032
rect 17720 45300 18278 46032
rect 22710 45300 23268 46032
rect 27700 45300 28258 46032
rect 32690 45300 33248 46032
rect 37680 45300 38238 46032
rect 42670 45300 43228 46032
rect 47660 45300 48218 46032
rect 52650 45300 53208 46032
rect 57640 45300 58198 46032
rect 62630 45300 63188 46032
rect 67620 45300 68178 46032
rect 72610 45300 73168 46032
rect 77600 45300 78158 46032
rect 2740 44360 2810 44820
rect 7730 44360 7800 44820
rect 12720 44360 12790 44820
rect 17710 44360 17780 44820
rect 22700 44360 22770 44820
rect 27690 44360 27760 44820
rect 32680 44360 32750 44820
rect 37670 44360 37740 44820
rect 42660 44360 42730 44820
rect 47650 44360 47720 44820
rect 52640 44360 52710 44820
rect 57630 44360 57700 44820
rect 62620 44360 62690 44820
rect 67610 44360 67680 44820
rect 72600 44360 72670 44820
rect 77590 44360 77660 44820
rect 2750 43590 3308 44322
rect 7740 43590 8298 44322
rect 12730 43590 13288 44322
rect 17720 43590 18278 44322
rect 22710 43590 23268 44322
rect 27700 43590 28258 44322
rect 32690 43590 33248 44322
rect 37680 43590 38238 44322
rect 42670 43590 43228 44322
rect 47660 43590 48218 44322
rect 52650 43590 53208 44322
rect 57640 43590 58198 44322
rect 62630 43590 63188 44322
rect 67620 43590 68178 44322
rect 72610 43590 73168 44322
rect 77600 43590 78158 44322
rect 2740 42650 2810 43110
rect 7730 42650 7800 43110
rect 12720 42650 12790 43110
rect 17710 42650 17780 43110
rect 22700 42650 22770 43110
rect 27690 42650 27760 43110
rect 32680 42650 32750 43110
rect 37670 42650 37740 43110
rect 42660 42650 42730 43110
rect 47650 42650 47720 43110
rect 52640 42650 52710 43110
rect 57630 42650 57700 43110
rect 62620 42650 62690 43110
rect 67610 42650 67680 43110
rect 72600 42650 72670 43110
rect 77590 42650 77660 43110
rect 2750 41880 3308 42612
rect 7740 41880 8298 42612
rect 12730 41880 13288 42612
rect 17720 41880 18278 42612
rect 22710 41880 23268 42612
rect 27700 41880 28258 42612
rect 32690 41880 33248 42612
rect 37680 41880 38238 42612
rect 42670 41880 43228 42612
rect 47660 41880 48218 42612
rect 52650 41880 53208 42612
rect 57640 41880 58198 42612
rect 62630 41880 63188 42612
rect 67620 41880 68178 42612
rect 72610 41880 73168 42612
rect 77600 41880 78158 42612
rect 2740 40940 2810 41400
rect 7730 40940 7800 41400
rect 12720 40940 12790 41400
rect 17710 40940 17780 41400
rect 22700 40940 22770 41400
rect 27690 40940 27760 41400
rect 32680 40940 32750 41400
rect 37670 40940 37740 41400
rect 42660 40940 42730 41400
rect 47650 40940 47720 41400
rect 52640 40940 52710 41400
rect 57630 40940 57700 41400
rect 62620 40940 62690 41400
rect 67610 40940 67680 41400
rect 72600 40940 72670 41400
rect 77590 40940 77660 41400
rect 2750 40170 3308 40902
rect 7740 40170 8298 40902
rect 12730 40170 13288 40902
rect 17720 40170 18278 40902
rect 22710 40170 23268 40902
rect 27700 40170 28258 40902
rect 32690 40170 33248 40902
rect 37680 40170 38238 40902
rect 42670 40170 43228 40902
rect 47660 40170 48218 40902
rect 52650 40170 53208 40902
rect 57640 40170 58198 40902
rect 62630 40170 63188 40902
rect 67620 40170 68178 40902
rect 72610 40170 73168 40902
rect 77600 40170 78158 40902
<< nmos >>
rect 2960 66326 3160 66356
rect 2960 66016 3160 66046
rect 7950 66326 8150 66356
rect 7950 66016 8150 66046
rect 12940 66326 13140 66356
rect 12940 66016 13140 66046
rect 17930 66326 18130 66356
rect 17930 66016 18130 66046
rect 22920 66326 23120 66356
rect 22920 66016 23120 66046
rect 27910 66326 28110 66356
rect 27910 66016 28110 66046
rect 32900 66326 33100 66356
rect 32900 66016 33100 66046
rect 37890 66326 38090 66356
rect 37890 66016 38090 66046
rect 42880 66326 43080 66356
rect 42880 66016 43080 66046
rect 47870 66326 48070 66356
rect 47870 66016 48070 66046
rect 52860 66326 53060 66356
rect 52860 66016 53060 66046
rect 57850 66326 58050 66356
rect 57850 66016 58050 66046
rect 62840 66326 63040 66356
rect 62840 66016 63040 66046
rect 67830 66326 68030 66356
rect 67830 66016 68030 66046
rect 72820 66326 73020 66356
rect 72820 66016 73020 66046
rect 77810 66326 78010 66356
rect 77810 66016 78010 66046
rect 2960 64616 3160 64646
rect 2960 64306 3160 64336
rect 7950 64616 8150 64646
rect 7950 64306 8150 64336
rect 12940 64616 13140 64646
rect 12940 64306 13140 64336
rect 17930 64616 18130 64646
rect 17930 64306 18130 64336
rect 22920 64616 23120 64646
rect 22920 64306 23120 64336
rect 27910 64616 28110 64646
rect 27910 64306 28110 64336
rect 32900 64616 33100 64646
rect 32900 64306 33100 64336
rect 37890 64616 38090 64646
rect 37890 64306 38090 64336
rect 42880 64616 43080 64646
rect 42880 64306 43080 64336
rect 47870 64616 48070 64646
rect 47870 64306 48070 64336
rect 52860 64616 53060 64646
rect 52860 64306 53060 64336
rect 57850 64616 58050 64646
rect 57850 64306 58050 64336
rect 62840 64616 63040 64646
rect 62840 64306 63040 64336
rect 67830 64616 68030 64646
rect 67830 64306 68030 64336
rect 72820 64616 73020 64646
rect 72820 64306 73020 64336
rect 77810 64616 78010 64646
rect 77810 64306 78010 64336
rect 2960 62906 3160 62936
rect 2960 62596 3160 62626
rect 7950 62906 8150 62936
rect 7950 62596 8150 62626
rect 12940 62906 13140 62936
rect 12940 62596 13140 62626
rect 17930 62906 18130 62936
rect 17930 62596 18130 62626
rect 22920 62906 23120 62936
rect 22920 62596 23120 62626
rect 27910 62906 28110 62936
rect 27910 62596 28110 62626
rect 32900 62906 33100 62936
rect 32900 62596 33100 62626
rect 37890 62906 38090 62936
rect 37890 62596 38090 62626
rect 42880 62906 43080 62936
rect 42880 62596 43080 62626
rect 47870 62906 48070 62936
rect 47870 62596 48070 62626
rect 52860 62906 53060 62936
rect 52860 62596 53060 62626
rect 57850 62906 58050 62936
rect 57850 62596 58050 62626
rect 62840 62906 63040 62936
rect 62840 62596 63040 62626
rect 67830 62906 68030 62936
rect 67830 62596 68030 62626
rect 72820 62906 73020 62936
rect 72820 62596 73020 62626
rect 77810 62906 78010 62936
rect 77810 62596 78010 62626
rect 2960 61196 3160 61226
rect 2960 60886 3160 60916
rect 7950 61196 8150 61226
rect 7950 60886 8150 60916
rect 12940 61196 13140 61226
rect 12940 60886 13140 60916
rect 17930 61196 18130 61226
rect 17930 60886 18130 60916
rect 22920 61196 23120 61226
rect 22920 60886 23120 60916
rect 27910 61196 28110 61226
rect 27910 60886 28110 60916
rect 32900 61196 33100 61226
rect 32900 60886 33100 60916
rect 37890 61196 38090 61226
rect 37890 60886 38090 60916
rect 42880 61196 43080 61226
rect 42880 60886 43080 60916
rect 47870 61196 48070 61226
rect 47870 60886 48070 60916
rect 52860 61196 53060 61226
rect 52860 60886 53060 60916
rect 57850 61196 58050 61226
rect 57850 60886 58050 60916
rect 62840 61196 63040 61226
rect 62840 60886 63040 60916
rect 67830 61196 68030 61226
rect 67830 60886 68030 60916
rect 72820 61196 73020 61226
rect 72820 60886 73020 60916
rect 77810 61196 78010 61226
rect 77810 60886 78010 60916
rect 2960 59486 3160 59516
rect 2960 59176 3160 59206
rect 7950 59486 8150 59516
rect 7950 59176 8150 59206
rect 12940 59486 13140 59516
rect 12940 59176 13140 59206
rect 17930 59486 18130 59516
rect 17930 59176 18130 59206
rect 22920 59486 23120 59516
rect 22920 59176 23120 59206
rect 27910 59486 28110 59516
rect 27910 59176 28110 59206
rect 32900 59486 33100 59516
rect 32900 59176 33100 59206
rect 37890 59486 38090 59516
rect 37890 59176 38090 59206
rect 42880 59486 43080 59516
rect 42880 59176 43080 59206
rect 47870 59486 48070 59516
rect 47870 59176 48070 59206
rect 52860 59486 53060 59516
rect 52860 59176 53060 59206
rect 57850 59486 58050 59516
rect 57850 59176 58050 59206
rect 62840 59486 63040 59516
rect 62840 59176 63040 59206
rect 67830 59486 68030 59516
rect 67830 59176 68030 59206
rect 72820 59486 73020 59516
rect 72820 59176 73020 59206
rect 77810 59486 78010 59516
rect 77810 59176 78010 59206
rect 2960 57776 3160 57806
rect 2960 57466 3160 57496
rect 7950 57776 8150 57806
rect 7950 57466 8150 57496
rect 12940 57776 13140 57806
rect 12940 57466 13140 57496
rect 17930 57776 18130 57806
rect 17930 57466 18130 57496
rect 22920 57776 23120 57806
rect 22920 57466 23120 57496
rect 27910 57776 28110 57806
rect 27910 57466 28110 57496
rect 32900 57776 33100 57806
rect 32900 57466 33100 57496
rect 37890 57776 38090 57806
rect 37890 57466 38090 57496
rect 42880 57776 43080 57806
rect 42880 57466 43080 57496
rect 47870 57776 48070 57806
rect 47870 57466 48070 57496
rect 52860 57776 53060 57806
rect 52860 57466 53060 57496
rect 57850 57776 58050 57806
rect 57850 57466 58050 57496
rect 62840 57776 63040 57806
rect 62840 57466 63040 57496
rect 67830 57776 68030 57806
rect 67830 57466 68030 57496
rect 72820 57776 73020 57806
rect 72820 57466 73020 57496
rect 77810 57776 78010 57806
rect 77810 57466 78010 57496
rect 2960 56066 3160 56096
rect 2960 55756 3160 55786
rect 7950 56066 8150 56096
rect 7950 55756 8150 55786
rect 12940 56066 13140 56096
rect 12940 55756 13140 55786
rect 17930 56066 18130 56096
rect 17930 55756 18130 55786
rect 22920 56066 23120 56096
rect 22920 55756 23120 55786
rect 27910 56066 28110 56096
rect 27910 55756 28110 55786
rect 32900 56066 33100 56096
rect 32900 55756 33100 55786
rect 37890 56066 38090 56096
rect 37890 55756 38090 55786
rect 42880 56066 43080 56096
rect 42880 55756 43080 55786
rect 47870 56066 48070 56096
rect 47870 55756 48070 55786
rect 52860 56066 53060 56096
rect 52860 55756 53060 55786
rect 57850 56066 58050 56096
rect 57850 55756 58050 55786
rect 62840 56066 63040 56096
rect 62840 55756 63040 55786
rect 67830 56066 68030 56096
rect 67830 55756 68030 55786
rect 72820 56066 73020 56096
rect 72820 55756 73020 55786
rect 77810 56066 78010 56096
rect 77810 55756 78010 55786
rect 2960 54356 3160 54386
rect 2960 54046 3160 54076
rect 7950 54356 8150 54386
rect 7950 54046 8150 54076
rect 12940 54356 13140 54386
rect 12940 54046 13140 54076
rect 17930 54356 18130 54386
rect 17930 54046 18130 54076
rect 22920 54356 23120 54386
rect 22920 54046 23120 54076
rect 27910 54356 28110 54386
rect 27910 54046 28110 54076
rect 32900 54356 33100 54386
rect 32900 54046 33100 54076
rect 37890 54356 38090 54386
rect 37890 54046 38090 54076
rect 42880 54356 43080 54386
rect 42880 54046 43080 54076
rect 47870 54356 48070 54386
rect 47870 54046 48070 54076
rect 52860 54356 53060 54386
rect 52860 54046 53060 54076
rect 57850 54356 58050 54386
rect 57850 54046 58050 54076
rect 62840 54356 63040 54386
rect 62840 54046 63040 54076
rect 67830 54356 68030 54386
rect 67830 54046 68030 54076
rect 72820 54356 73020 54386
rect 72820 54046 73020 54076
rect 77810 54356 78010 54386
rect 77810 54046 78010 54076
rect 2960 52646 3160 52676
rect 2960 52336 3160 52366
rect 7950 52646 8150 52676
rect 7950 52336 8150 52366
rect 12940 52646 13140 52676
rect 12940 52336 13140 52366
rect 17930 52646 18130 52676
rect 17930 52336 18130 52366
rect 22920 52646 23120 52676
rect 22920 52336 23120 52366
rect 27910 52646 28110 52676
rect 27910 52336 28110 52366
rect 32900 52646 33100 52676
rect 32900 52336 33100 52366
rect 37890 52646 38090 52676
rect 37890 52336 38090 52366
rect 42880 52646 43080 52676
rect 42880 52336 43080 52366
rect 47870 52646 48070 52676
rect 47870 52336 48070 52366
rect 52860 52646 53060 52676
rect 52860 52336 53060 52366
rect 57850 52646 58050 52676
rect 57850 52336 58050 52366
rect 62840 52646 63040 52676
rect 62840 52336 63040 52366
rect 67830 52646 68030 52676
rect 67830 52336 68030 52366
rect 72820 52646 73020 52676
rect 72820 52336 73020 52366
rect 77810 52646 78010 52676
rect 77810 52336 78010 52366
rect 2960 50936 3160 50966
rect 2960 50626 3160 50656
rect 7950 50936 8150 50966
rect 7950 50626 8150 50656
rect 12940 50936 13140 50966
rect 12940 50626 13140 50656
rect 17930 50936 18130 50966
rect 17930 50626 18130 50656
rect 22920 50936 23120 50966
rect 22920 50626 23120 50656
rect 27910 50936 28110 50966
rect 27910 50626 28110 50656
rect 32900 50936 33100 50966
rect 32900 50626 33100 50656
rect 37890 50936 38090 50966
rect 37890 50626 38090 50656
rect 42880 50936 43080 50966
rect 42880 50626 43080 50656
rect 47870 50936 48070 50966
rect 47870 50626 48070 50656
rect 52860 50936 53060 50966
rect 52860 50626 53060 50656
rect 57850 50936 58050 50966
rect 57850 50626 58050 50656
rect 62840 50936 63040 50966
rect 62840 50626 63040 50656
rect 67830 50936 68030 50966
rect 67830 50626 68030 50656
rect 72820 50936 73020 50966
rect 72820 50626 73020 50656
rect 77810 50936 78010 50966
rect 77810 50626 78010 50656
rect 2960 49226 3160 49256
rect 2960 48916 3160 48946
rect 7950 49226 8150 49256
rect 7950 48916 8150 48946
rect 12940 49226 13140 49256
rect 12940 48916 13140 48946
rect 17930 49226 18130 49256
rect 17930 48916 18130 48946
rect 22920 49226 23120 49256
rect 22920 48916 23120 48946
rect 27910 49226 28110 49256
rect 27910 48916 28110 48946
rect 32900 49226 33100 49256
rect 32900 48916 33100 48946
rect 37890 49226 38090 49256
rect 37890 48916 38090 48946
rect 42880 49226 43080 49256
rect 42880 48916 43080 48946
rect 47870 49226 48070 49256
rect 47870 48916 48070 48946
rect 52860 49226 53060 49256
rect 52860 48916 53060 48946
rect 57850 49226 58050 49256
rect 57850 48916 58050 48946
rect 62840 49226 63040 49256
rect 62840 48916 63040 48946
rect 67830 49226 68030 49256
rect 67830 48916 68030 48946
rect 72820 49226 73020 49256
rect 72820 48916 73020 48946
rect 77810 49226 78010 49256
rect 77810 48916 78010 48946
rect 2960 47516 3160 47546
rect 2960 47206 3160 47236
rect 7950 47516 8150 47546
rect 7950 47206 8150 47236
rect 12940 47516 13140 47546
rect 12940 47206 13140 47236
rect 17930 47516 18130 47546
rect 17930 47206 18130 47236
rect 22920 47516 23120 47546
rect 22920 47206 23120 47236
rect 27910 47516 28110 47546
rect 27910 47206 28110 47236
rect 32900 47516 33100 47546
rect 32900 47206 33100 47236
rect 37890 47516 38090 47546
rect 37890 47206 38090 47236
rect 42880 47516 43080 47546
rect 42880 47206 43080 47236
rect 47870 47516 48070 47546
rect 47870 47206 48070 47236
rect 52860 47516 53060 47546
rect 52860 47206 53060 47236
rect 57850 47516 58050 47546
rect 57850 47206 58050 47236
rect 62840 47516 63040 47546
rect 62840 47206 63040 47236
rect 67830 47516 68030 47546
rect 67830 47206 68030 47236
rect 72820 47516 73020 47546
rect 72820 47206 73020 47236
rect 77810 47516 78010 47546
rect 77810 47206 78010 47236
rect 2960 45806 3160 45836
rect 2960 45496 3160 45526
rect 7950 45806 8150 45836
rect 7950 45496 8150 45526
rect 12940 45806 13140 45836
rect 12940 45496 13140 45526
rect 17930 45806 18130 45836
rect 17930 45496 18130 45526
rect 22920 45806 23120 45836
rect 22920 45496 23120 45526
rect 27910 45806 28110 45836
rect 27910 45496 28110 45526
rect 32900 45806 33100 45836
rect 32900 45496 33100 45526
rect 37890 45806 38090 45836
rect 37890 45496 38090 45526
rect 42880 45806 43080 45836
rect 42880 45496 43080 45526
rect 47870 45806 48070 45836
rect 47870 45496 48070 45526
rect 52860 45806 53060 45836
rect 52860 45496 53060 45526
rect 57850 45806 58050 45836
rect 57850 45496 58050 45526
rect 62840 45806 63040 45836
rect 62840 45496 63040 45526
rect 67830 45806 68030 45836
rect 67830 45496 68030 45526
rect 72820 45806 73020 45836
rect 72820 45496 73020 45526
rect 77810 45806 78010 45836
rect 77810 45496 78010 45526
rect 2960 44096 3160 44126
rect 2960 43786 3160 43816
rect 7950 44096 8150 44126
rect 7950 43786 8150 43816
rect 12940 44096 13140 44126
rect 12940 43786 13140 43816
rect 17930 44096 18130 44126
rect 17930 43786 18130 43816
rect 22920 44096 23120 44126
rect 22920 43786 23120 43816
rect 27910 44096 28110 44126
rect 27910 43786 28110 43816
rect 32900 44096 33100 44126
rect 32900 43786 33100 43816
rect 37890 44096 38090 44126
rect 37890 43786 38090 43816
rect 42880 44096 43080 44126
rect 42880 43786 43080 43816
rect 47870 44096 48070 44126
rect 47870 43786 48070 43816
rect 52860 44096 53060 44126
rect 52860 43786 53060 43816
rect 57850 44096 58050 44126
rect 57850 43786 58050 43816
rect 62840 44096 63040 44126
rect 62840 43786 63040 43816
rect 67830 44096 68030 44126
rect 67830 43786 68030 43816
rect 72820 44096 73020 44126
rect 72820 43786 73020 43816
rect 77810 44096 78010 44126
rect 77810 43786 78010 43816
rect 2960 42386 3160 42416
rect 2960 42076 3160 42106
rect 7950 42386 8150 42416
rect 7950 42076 8150 42106
rect 12940 42386 13140 42416
rect 12940 42076 13140 42106
rect 17930 42386 18130 42416
rect 17930 42076 18130 42106
rect 22920 42386 23120 42416
rect 22920 42076 23120 42106
rect 27910 42386 28110 42416
rect 27910 42076 28110 42106
rect 32900 42386 33100 42416
rect 32900 42076 33100 42106
rect 37890 42386 38090 42416
rect 37890 42076 38090 42106
rect 42880 42386 43080 42416
rect 42880 42076 43080 42106
rect 47870 42386 48070 42416
rect 47870 42076 48070 42106
rect 52860 42386 53060 42416
rect 52860 42076 53060 42106
rect 57850 42386 58050 42416
rect 57850 42076 58050 42106
rect 62840 42386 63040 42416
rect 62840 42076 63040 42106
rect 67830 42386 68030 42416
rect 67830 42076 68030 42106
rect 72820 42386 73020 42416
rect 72820 42076 73020 42106
rect 77810 42386 78010 42416
rect 77810 42076 78010 42106
rect 2960 40676 3160 40706
rect 2960 40366 3160 40396
rect 7950 40676 8150 40706
rect 7950 40366 8150 40396
rect 12940 40676 13140 40706
rect 12940 40366 13140 40396
rect 17930 40676 18130 40706
rect 17930 40366 18130 40396
rect 22920 40676 23120 40706
rect 22920 40366 23120 40396
rect 27910 40676 28110 40706
rect 27910 40366 28110 40396
rect 32900 40676 33100 40706
rect 32900 40366 33100 40396
rect 37890 40676 38090 40706
rect 37890 40366 38090 40396
rect 42880 40676 43080 40706
rect 42880 40366 43080 40396
rect 47870 40676 48070 40706
rect 47870 40366 48070 40396
rect 52860 40676 53060 40706
rect 52860 40366 53060 40396
rect 57850 40676 58050 40706
rect 57850 40366 58050 40396
rect 62840 40676 63040 40706
rect 62840 40366 63040 40396
rect 67830 40676 68030 40706
rect 67830 40366 68030 40396
rect 72820 40676 73020 40706
rect 72820 40366 73020 40396
rect 77810 40676 78010 40706
rect 77810 40366 78010 40396
<< pmos >>
rect 3458 66326 3658 66356
rect 3458 66016 3658 66046
rect 8448 66326 8648 66356
rect 8448 66016 8648 66046
rect 13438 66326 13638 66356
rect 13438 66016 13638 66046
rect 18428 66326 18628 66356
rect 18428 66016 18628 66046
rect 23418 66326 23618 66356
rect 23418 66016 23618 66046
rect 28408 66326 28608 66356
rect 28408 66016 28608 66046
rect 33398 66326 33598 66356
rect 33398 66016 33598 66046
rect 38388 66326 38588 66356
rect 38388 66016 38588 66046
rect 43378 66326 43578 66356
rect 43378 66016 43578 66046
rect 48368 66326 48568 66356
rect 48368 66016 48568 66046
rect 53358 66326 53558 66356
rect 53358 66016 53558 66046
rect 58348 66326 58548 66356
rect 58348 66016 58548 66046
rect 63338 66326 63538 66356
rect 63338 66016 63538 66046
rect 68328 66326 68528 66356
rect 68328 66016 68528 66046
rect 73318 66326 73518 66356
rect 73318 66016 73518 66046
rect 78308 66326 78508 66356
rect 78308 66016 78508 66046
rect 3458 64616 3658 64646
rect 3458 64306 3658 64336
rect 8448 64616 8648 64646
rect 8448 64306 8648 64336
rect 13438 64616 13638 64646
rect 13438 64306 13638 64336
rect 18428 64616 18628 64646
rect 18428 64306 18628 64336
rect 23418 64616 23618 64646
rect 23418 64306 23618 64336
rect 28408 64616 28608 64646
rect 28408 64306 28608 64336
rect 33398 64616 33598 64646
rect 33398 64306 33598 64336
rect 38388 64616 38588 64646
rect 38388 64306 38588 64336
rect 43378 64616 43578 64646
rect 43378 64306 43578 64336
rect 48368 64616 48568 64646
rect 48368 64306 48568 64336
rect 53358 64616 53558 64646
rect 53358 64306 53558 64336
rect 58348 64616 58548 64646
rect 58348 64306 58548 64336
rect 63338 64616 63538 64646
rect 63338 64306 63538 64336
rect 68328 64616 68528 64646
rect 68328 64306 68528 64336
rect 73318 64616 73518 64646
rect 73318 64306 73518 64336
rect 78308 64616 78508 64646
rect 78308 64306 78508 64336
rect 3458 62906 3658 62936
rect 3458 62596 3658 62626
rect 8448 62906 8648 62936
rect 8448 62596 8648 62626
rect 13438 62906 13638 62936
rect 13438 62596 13638 62626
rect 18428 62906 18628 62936
rect 18428 62596 18628 62626
rect 23418 62906 23618 62936
rect 23418 62596 23618 62626
rect 28408 62906 28608 62936
rect 28408 62596 28608 62626
rect 33398 62906 33598 62936
rect 33398 62596 33598 62626
rect 38388 62906 38588 62936
rect 38388 62596 38588 62626
rect 43378 62906 43578 62936
rect 43378 62596 43578 62626
rect 48368 62906 48568 62936
rect 48368 62596 48568 62626
rect 53358 62906 53558 62936
rect 53358 62596 53558 62626
rect 58348 62906 58548 62936
rect 58348 62596 58548 62626
rect 63338 62906 63538 62936
rect 63338 62596 63538 62626
rect 68328 62906 68528 62936
rect 68328 62596 68528 62626
rect 73318 62906 73518 62936
rect 73318 62596 73518 62626
rect 78308 62906 78508 62936
rect 78308 62596 78508 62626
rect 3458 61196 3658 61226
rect 3458 60886 3658 60916
rect 8448 61196 8648 61226
rect 8448 60886 8648 60916
rect 13438 61196 13638 61226
rect 13438 60886 13638 60916
rect 18428 61196 18628 61226
rect 18428 60886 18628 60916
rect 23418 61196 23618 61226
rect 23418 60886 23618 60916
rect 28408 61196 28608 61226
rect 28408 60886 28608 60916
rect 33398 61196 33598 61226
rect 33398 60886 33598 60916
rect 38388 61196 38588 61226
rect 38388 60886 38588 60916
rect 43378 61196 43578 61226
rect 43378 60886 43578 60916
rect 48368 61196 48568 61226
rect 48368 60886 48568 60916
rect 53358 61196 53558 61226
rect 53358 60886 53558 60916
rect 58348 61196 58548 61226
rect 58348 60886 58548 60916
rect 63338 61196 63538 61226
rect 63338 60886 63538 60916
rect 68328 61196 68528 61226
rect 68328 60886 68528 60916
rect 73318 61196 73518 61226
rect 73318 60886 73518 60916
rect 78308 61196 78508 61226
rect 78308 60886 78508 60916
rect 3458 59486 3658 59516
rect 3458 59176 3658 59206
rect 8448 59486 8648 59516
rect 8448 59176 8648 59206
rect 13438 59486 13638 59516
rect 13438 59176 13638 59206
rect 18428 59486 18628 59516
rect 18428 59176 18628 59206
rect 23418 59486 23618 59516
rect 23418 59176 23618 59206
rect 28408 59486 28608 59516
rect 28408 59176 28608 59206
rect 33398 59486 33598 59516
rect 33398 59176 33598 59206
rect 38388 59486 38588 59516
rect 38388 59176 38588 59206
rect 43378 59486 43578 59516
rect 43378 59176 43578 59206
rect 48368 59486 48568 59516
rect 48368 59176 48568 59206
rect 53358 59486 53558 59516
rect 53358 59176 53558 59206
rect 58348 59486 58548 59516
rect 58348 59176 58548 59206
rect 63338 59486 63538 59516
rect 63338 59176 63538 59206
rect 68328 59486 68528 59516
rect 68328 59176 68528 59206
rect 73318 59486 73518 59516
rect 73318 59176 73518 59206
rect 78308 59486 78508 59516
rect 78308 59176 78508 59206
rect 3458 57776 3658 57806
rect 3458 57466 3658 57496
rect 8448 57776 8648 57806
rect 8448 57466 8648 57496
rect 13438 57776 13638 57806
rect 13438 57466 13638 57496
rect 18428 57776 18628 57806
rect 18428 57466 18628 57496
rect 23418 57776 23618 57806
rect 23418 57466 23618 57496
rect 28408 57776 28608 57806
rect 28408 57466 28608 57496
rect 33398 57776 33598 57806
rect 33398 57466 33598 57496
rect 38388 57776 38588 57806
rect 38388 57466 38588 57496
rect 43378 57776 43578 57806
rect 43378 57466 43578 57496
rect 48368 57776 48568 57806
rect 48368 57466 48568 57496
rect 53358 57776 53558 57806
rect 53358 57466 53558 57496
rect 58348 57776 58548 57806
rect 58348 57466 58548 57496
rect 63338 57776 63538 57806
rect 63338 57466 63538 57496
rect 68328 57776 68528 57806
rect 68328 57466 68528 57496
rect 73318 57776 73518 57806
rect 73318 57466 73518 57496
rect 78308 57776 78508 57806
rect 78308 57466 78508 57496
rect 3458 56066 3658 56096
rect 3458 55756 3658 55786
rect 8448 56066 8648 56096
rect 8448 55756 8648 55786
rect 13438 56066 13638 56096
rect 13438 55756 13638 55786
rect 18428 56066 18628 56096
rect 18428 55756 18628 55786
rect 23418 56066 23618 56096
rect 23418 55756 23618 55786
rect 28408 56066 28608 56096
rect 28408 55756 28608 55786
rect 33398 56066 33598 56096
rect 33398 55756 33598 55786
rect 38388 56066 38588 56096
rect 38388 55756 38588 55786
rect 43378 56066 43578 56096
rect 43378 55756 43578 55786
rect 48368 56066 48568 56096
rect 48368 55756 48568 55786
rect 53358 56066 53558 56096
rect 53358 55756 53558 55786
rect 58348 56066 58548 56096
rect 58348 55756 58548 55786
rect 63338 56066 63538 56096
rect 63338 55756 63538 55786
rect 68328 56066 68528 56096
rect 68328 55756 68528 55786
rect 73318 56066 73518 56096
rect 73318 55756 73518 55786
rect 78308 56066 78508 56096
rect 78308 55756 78508 55786
rect 3458 54356 3658 54386
rect 3458 54046 3658 54076
rect 8448 54356 8648 54386
rect 8448 54046 8648 54076
rect 13438 54356 13638 54386
rect 13438 54046 13638 54076
rect 18428 54356 18628 54386
rect 18428 54046 18628 54076
rect 23418 54356 23618 54386
rect 23418 54046 23618 54076
rect 28408 54356 28608 54386
rect 28408 54046 28608 54076
rect 33398 54356 33598 54386
rect 33398 54046 33598 54076
rect 38388 54356 38588 54386
rect 38388 54046 38588 54076
rect 43378 54356 43578 54386
rect 43378 54046 43578 54076
rect 48368 54356 48568 54386
rect 48368 54046 48568 54076
rect 53358 54356 53558 54386
rect 53358 54046 53558 54076
rect 58348 54356 58548 54386
rect 58348 54046 58548 54076
rect 63338 54356 63538 54386
rect 63338 54046 63538 54076
rect 68328 54356 68528 54386
rect 68328 54046 68528 54076
rect 73318 54356 73518 54386
rect 73318 54046 73518 54076
rect 78308 54356 78508 54386
rect 78308 54046 78508 54076
rect 3458 52646 3658 52676
rect 3458 52336 3658 52366
rect 8448 52646 8648 52676
rect 8448 52336 8648 52366
rect 13438 52646 13638 52676
rect 13438 52336 13638 52366
rect 18428 52646 18628 52676
rect 18428 52336 18628 52366
rect 23418 52646 23618 52676
rect 23418 52336 23618 52366
rect 28408 52646 28608 52676
rect 28408 52336 28608 52366
rect 33398 52646 33598 52676
rect 33398 52336 33598 52366
rect 38388 52646 38588 52676
rect 38388 52336 38588 52366
rect 43378 52646 43578 52676
rect 43378 52336 43578 52366
rect 48368 52646 48568 52676
rect 48368 52336 48568 52366
rect 53358 52646 53558 52676
rect 53358 52336 53558 52366
rect 58348 52646 58548 52676
rect 58348 52336 58548 52366
rect 63338 52646 63538 52676
rect 63338 52336 63538 52366
rect 68328 52646 68528 52676
rect 68328 52336 68528 52366
rect 73318 52646 73518 52676
rect 73318 52336 73518 52366
rect 78308 52646 78508 52676
rect 78308 52336 78508 52366
rect 3458 50936 3658 50966
rect 3458 50626 3658 50656
rect 8448 50936 8648 50966
rect 8448 50626 8648 50656
rect 13438 50936 13638 50966
rect 13438 50626 13638 50656
rect 18428 50936 18628 50966
rect 18428 50626 18628 50656
rect 23418 50936 23618 50966
rect 23418 50626 23618 50656
rect 28408 50936 28608 50966
rect 28408 50626 28608 50656
rect 33398 50936 33598 50966
rect 33398 50626 33598 50656
rect 38388 50936 38588 50966
rect 38388 50626 38588 50656
rect 43378 50936 43578 50966
rect 43378 50626 43578 50656
rect 48368 50936 48568 50966
rect 48368 50626 48568 50656
rect 53358 50936 53558 50966
rect 53358 50626 53558 50656
rect 58348 50936 58548 50966
rect 58348 50626 58548 50656
rect 63338 50936 63538 50966
rect 63338 50626 63538 50656
rect 68328 50936 68528 50966
rect 68328 50626 68528 50656
rect 73318 50936 73518 50966
rect 73318 50626 73518 50656
rect 78308 50936 78508 50966
rect 78308 50626 78508 50656
rect 3458 49226 3658 49256
rect 3458 48916 3658 48946
rect 8448 49226 8648 49256
rect 8448 48916 8648 48946
rect 13438 49226 13638 49256
rect 13438 48916 13638 48946
rect 18428 49226 18628 49256
rect 18428 48916 18628 48946
rect 23418 49226 23618 49256
rect 23418 48916 23618 48946
rect 28408 49226 28608 49256
rect 28408 48916 28608 48946
rect 33398 49226 33598 49256
rect 33398 48916 33598 48946
rect 38388 49226 38588 49256
rect 38388 48916 38588 48946
rect 43378 49226 43578 49256
rect 43378 48916 43578 48946
rect 48368 49226 48568 49256
rect 48368 48916 48568 48946
rect 53358 49226 53558 49256
rect 53358 48916 53558 48946
rect 58348 49226 58548 49256
rect 58348 48916 58548 48946
rect 63338 49226 63538 49256
rect 63338 48916 63538 48946
rect 68328 49226 68528 49256
rect 68328 48916 68528 48946
rect 73318 49226 73518 49256
rect 73318 48916 73518 48946
rect 78308 49226 78508 49256
rect 78308 48916 78508 48946
rect 3458 47516 3658 47546
rect 3458 47206 3658 47236
rect 8448 47516 8648 47546
rect 8448 47206 8648 47236
rect 13438 47516 13638 47546
rect 13438 47206 13638 47236
rect 18428 47516 18628 47546
rect 18428 47206 18628 47236
rect 23418 47516 23618 47546
rect 23418 47206 23618 47236
rect 28408 47516 28608 47546
rect 28408 47206 28608 47236
rect 33398 47516 33598 47546
rect 33398 47206 33598 47236
rect 38388 47516 38588 47546
rect 38388 47206 38588 47236
rect 43378 47516 43578 47546
rect 43378 47206 43578 47236
rect 48368 47516 48568 47546
rect 48368 47206 48568 47236
rect 53358 47516 53558 47546
rect 53358 47206 53558 47236
rect 58348 47516 58548 47546
rect 58348 47206 58548 47236
rect 63338 47516 63538 47546
rect 63338 47206 63538 47236
rect 68328 47516 68528 47546
rect 68328 47206 68528 47236
rect 73318 47516 73518 47546
rect 73318 47206 73518 47236
rect 78308 47516 78508 47546
rect 78308 47206 78508 47236
rect 3458 45806 3658 45836
rect 3458 45496 3658 45526
rect 8448 45806 8648 45836
rect 8448 45496 8648 45526
rect 13438 45806 13638 45836
rect 13438 45496 13638 45526
rect 18428 45806 18628 45836
rect 18428 45496 18628 45526
rect 23418 45806 23618 45836
rect 23418 45496 23618 45526
rect 28408 45806 28608 45836
rect 28408 45496 28608 45526
rect 33398 45806 33598 45836
rect 33398 45496 33598 45526
rect 38388 45806 38588 45836
rect 38388 45496 38588 45526
rect 43378 45806 43578 45836
rect 43378 45496 43578 45526
rect 48368 45806 48568 45836
rect 48368 45496 48568 45526
rect 53358 45806 53558 45836
rect 53358 45496 53558 45526
rect 58348 45806 58548 45836
rect 58348 45496 58548 45526
rect 63338 45806 63538 45836
rect 63338 45496 63538 45526
rect 68328 45806 68528 45836
rect 68328 45496 68528 45526
rect 73318 45806 73518 45836
rect 73318 45496 73518 45526
rect 78308 45806 78508 45836
rect 78308 45496 78508 45526
rect 3458 44096 3658 44126
rect 3458 43786 3658 43816
rect 8448 44096 8648 44126
rect 8448 43786 8648 43816
rect 13438 44096 13638 44126
rect 13438 43786 13638 43816
rect 18428 44096 18628 44126
rect 18428 43786 18628 43816
rect 23418 44096 23618 44126
rect 23418 43786 23618 43816
rect 28408 44096 28608 44126
rect 28408 43786 28608 43816
rect 33398 44096 33598 44126
rect 33398 43786 33598 43816
rect 38388 44096 38588 44126
rect 38388 43786 38588 43816
rect 43378 44096 43578 44126
rect 43378 43786 43578 43816
rect 48368 44096 48568 44126
rect 48368 43786 48568 43816
rect 53358 44096 53558 44126
rect 53358 43786 53558 43816
rect 58348 44096 58548 44126
rect 58348 43786 58548 43816
rect 63338 44096 63538 44126
rect 63338 43786 63538 43816
rect 68328 44096 68528 44126
rect 68328 43786 68528 43816
rect 73318 44096 73518 44126
rect 73318 43786 73518 43816
rect 78308 44096 78508 44126
rect 78308 43786 78508 43816
rect 3458 42386 3658 42416
rect 3458 42076 3658 42106
rect 8448 42386 8648 42416
rect 8448 42076 8648 42106
rect 13438 42386 13638 42416
rect 13438 42076 13638 42106
rect 18428 42386 18628 42416
rect 18428 42076 18628 42106
rect 23418 42386 23618 42416
rect 23418 42076 23618 42106
rect 28408 42386 28608 42416
rect 28408 42076 28608 42106
rect 33398 42386 33598 42416
rect 33398 42076 33598 42106
rect 38388 42386 38588 42416
rect 38388 42076 38588 42106
rect 43378 42386 43578 42416
rect 43378 42076 43578 42106
rect 48368 42386 48568 42416
rect 48368 42076 48568 42106
rect 53358 42386 53558 42416
rect 53358 42076 53558 42106
rect 58348 42386 58548 42416
rect 58348 42076 58548 42106
rect 63338 42386 63538 42416
rect 63338 42076 63538 42106
rect 68328 42386 68528 42416
rect 68328 42076 68528 42106
rect 73318 42386 73518 42416
rect 73318 42076 73518 42106
rect 78308 42386 78508 42416
rect 78308 42076 78508 42106
rect 3458 40676 3658 40706
rect 3458 40366 3658 40396
rect 8448 40676 8648 40706
rect 8448 40366 8648 40396
rect 13438 40676 13638 40706
rect 13438 40366 13638 40396
rect 18428 40676 18628 40706
rect 18428 40366 18628 40396
rect 23418 40676 23618 40706
rect 23418 40366 23618 40396
rect 28408 40676 28608 40706
rect 28408 40366 28608 40396
rect 33398 40676 33598 40706
rect 33398 40366 33598 40396
rect 38388 40676 38588 40706
rect 38388 40366 38588 40396
rect 43378 40676 43578 40706
rect 43378 40366 43578 40396
rect 48368 40676 48568 40706
rect 48368 40366 48568 40396
rect 53358 40676 53558 40706
rect 53358 40366 53558 40396
rect 58348 40676 58548 40706
rect 58348 40366 58548 40396
rect 63338 40676 63538 40706
rect 63338 40366 63538 40396
rect 68328 40676 68528 40706
rect 68328 40366 68528 40396
rect 73318 40676 73518 40706
rect 73318 40366 73518 40396
rect 78308 40676 78508 40706
rect 78308 40366 78508 40396
<< ndiff >>
rect 2960 66402 3160 66414
rect 2960 66368 2972 66402
rect 3148 66368 3160 66402
rect 2960 66356 3160 66368
rect 2960 66314 3160 66326
rect 2960 66280 2972 66314
rect 3148 66280 3160 66314
rect 2960 66268 3160 66280
rect 2960 66092 3160 66104
rect 2960 66058 2972 66092
rect 3148 66058 3160 66092
rect 2960 66046 3160 66058
rect 2960 66004 3160 66016
rect 2960 65970 2972 66004
rect 3148 65970 3160 66004
rect 2960 65958 3160 65970
rect 7950 66402 8150 66414
rect 7950 66368 7962 66402
rect 8138 66368 8150 66402
rect 7950 66356 8150 66368
rect 7950 66314 8150 66326
rect 7950 66280 7962 66314
rect 8138 66280 8150 66314
rect 7950 66268 8150 66280
rect 7950 66092 8150 66104
rect 7950 66058 7962 66092
rect 8138 66058 8150 66092
rect 7950 66046 8150 66058
rect 7950 66004 8150 66016
rect 7950 65970 7962 66004
rect 8138 65970 8150 66004
rect 7950 65958 8150 65970
rect 12940 66402 13140 66414
rect 12940 66368 12952 66402
rect 13128 66368 13140 66402
rect 12940 66356 13140 66368
rect 12940 66314 13140 66326
rect 12940 66280 12952 66314
rect 13128 66280 13140 66314
rect 12940 66268 13140 66280
rect 12940 66092 13140 66104
rect 12940 66058 12952 66092
rect 13128 66058 13140 66092
rect 12940 66046 13140 66058
rect 12940 66004 13140 66016
rect 12940 65970 12952 66004
rect 13128 65970 13140 66004
rect 12940 65958 13140 65970
rect 17930 66402 18130 66414
rect 17930 66368 17942 66402
rect 18118 66368 18130 66402
rect 17930 66356 18130 66368
rect 17930 66314 18130 66326
rect 17930 66280 17942 66314
rect 18118 66280 18130 66314
rect 17930 66268 18130 66280
rect 17930 66092 18130 66104
rect 17930 66058 17942 66092
rect 18118 66058 18130 66092
rect 17930 66046 18130 66058
rect 17930 66004 18130 66016
rect 17930 65970 17942 66004
rect 18118 65970 18130 66004
rect 17930 65958 18130 65970
rect 22920 66402 23120 66414
rect 22920 66368 22932 66402
rect 23108 66368 23120 66402
rect 22920 66356 23120 66368
rect 22920 66314 23120 66326
rect 22920 66280 22932 66314
rect 23108 66280 23120 66314
rect 22920 66268 23120 66280
rect 22920 66092 23120 66104
rect 22920 66058 22932 66092
rect 23108 66058 23120 66092
rect 22920 66046 23120 66058
rect 22920 66004 23120 66016
rect 22920 65970 22932 66004
rect 23108 65970 23120 66004
rect 22920 65958 23120 65970
rect 27910 66402 28110 66414
rect 27910 66368 27922 66402
rect 28098 66368 28110 66402
rect 27910 66356 28110 66368
rect 27910 66314 28110 66326
rect 27910 66280 27922 66314
rect 28098 66280 28110 66314
rect 27910 66268 28110 66280
rect 27910 66092 28110 66104
rect 27910 66058 27922 66092
rect 28098 66058 28110 66092
rect 27910 66046 28110 66058
rect 27910 66004 28110 66016
rect 27910 65970 27922 66004
rect 28098 65970 28110 66004
rect 27910 65958 28110 65970
rect 32900 66402 33100 66414
rect 32900 66368 32912 66402
rect 33088 66368 33100 66402
rect 32900 66356 33100 66368
rect 32900 66314 33100 66326
rect 32900 66280 32912 66314
rect 33088 66280 33100 66314
rect 32900 66268 33100 66280
rect 32900 66092 33100 66104
rect 32900 66058 32912 66092
rect 33088 66058 33100 66092
rect 32900 66046 33100 66058
rect 32900 66004 33100 66016
rect 32900 65970 32912 66004
rect 33088 65970 33100 66004
rect 32900 65958 33100 65970
rect 37890 66402 38090 66414
rect 37890 66368 37902 66402
rect 38078 66368 38090 66402
rect 37890 66356 38090 66368
rect 37890 66314 38090 66326
rect 37890 66280 37902 66314
rect 38078 66280 38090 66314
rect 37890 66268 38090 66280
rect 37890 66092 38090 66104
rect 37890 66058 37902 66092
rect 38078 66058 38090 66092
rect 37890 66046 38090 66058
rect 37890 66004 38090 66016
rect 37890 65970 37902 66004
rect 38078 65970 38090 66004
rect 37890 65958 38090 65970
rect 42880 66402 43080 66414
rect 42880 66368 42892 66402
rect 43068 66368 43080 66402
rect 42880 66356 43080 66368
rect 42880 66314 43080 66326
rect 42880 66280 42892 66314
rect 43068 66280 43080 66314
rect 42880 66268 43080 66280
rect 42880 66092 43080 66104
rect 42880 66058 42892 66092
rect 43068 66058 43080 66092
rect 42880 66046 43080 66058
rect 42880 66004 43080 66016
rect 42880 65970 42892 66004
rect 43068 65970 43080 66004
rect 42880 65958 43080 65970
rect 47870 66402 48070 66414
rect 47870 66368 47882 66402
rect 48058 66368 48070 66402
rect 47870 66356 48070 66368
rect 47870 66314 48070 66326
rect 47870 66280 47882 66314
rect 48058 66280 48070 66314
rect 47870 66268 48070 66280
rect 47870 66092 48070 66104
rect 47870 66058 47882 66092
rect 48058 66058 48070 66092
rect 47870 66046 48070 66058
rect 47870 66004 48070 66016
rect 47870 65970 47882 66004
rect 48058 65970 48070 66004
rect 47870 65958 48070 65970
rect 52860 66402 53060 66414
rect 52860 66368 52872 66402
rect 53048 66368 53060 66402
rect 52860 66356 53060 66368
rect 52860 66314 53060 66326
rect 52860 66280 52872 66314
rect 53048 66280 53060 66314
rect 52860 66268 53060 66280
rect 52860 66092 53060 66104
rect 52860 66058 52872 66092
rect 53048 66058 53060 66092
rect 52860 66046 53060 66058
rect 52860 66004 53060 66016
rect 52860 65970 52872 66004
rect 53048 65970 53060 66004
rect 52860 65958 53060 65970
rect 57850 66402 58050 66414
rect 57850 66368 57862 66402
rect 58038 66368 58050 66402
rect 57850 66356 58050 66368
rect 57850 66314 58050 66326
rect 57850 66280 57862 66314
rect 58038 66280 58050 66314
rect 57850 66268 58050 66280
rect 57850 66092 58050 66104
rect 57850 66058 57862 66092
rect 58038 66058 58050 66092
rect 57850 66046 58050 66058
rect 57850 66004 58050 66016
rect 57850 65970 57862 66004
rect 58038 65970 58050 66004
rect 57850 65958 58050 65970
rect 62840 66402 63040 66414
rect 62840 66368 62852 66402
rect 63028 66368 63040 66402
rect 62840 66356 63040 66368
rect 62840 66314 63040 66326
rect 62840 66280 62852 66314
rect 63028 66280 63040 66314
rect 62840 66268 63040 66280
rect 62840 66092 63040 66104
rect 62840 66058 62852 66092
rect 63028 66058 63040 66092
rect 62840 66046 63040 66058
rect 62840 66004 63040 66016
rect 62840 65970 62852 66004
rect 63028 65970 63040 66004
rect 62840 65958 63040 65970
rect 67830 66402 68030 66414
rect 67830 66368 67842 66402
rect 68018 66368 68030 66402
rect 67830 66356 68030 66368
rect 67830 66314 68030 66326
rect 67830 66280 67842 66314
rect 68018 66280 68030 66314
rect 67830 66268 68030 66280
rect 67830 66092 68030 66104
rect 67830 66058 67842 66092
rect 68018 66058 68030 66092
rect 67830 66046 68030 66058
rect 67830 66004 68030 66016
rect 67830 65970 67842 66004
rect 68018 65970 68030 66004
rect 67830 65958 68030 65970
rect 72820 66402 73020 66414
rect 72820 66368 72832 66402
rect 73008 66368 73020 66402
rect 72820 66356 73020 66368
rect 72820 66314 73020 66326
rect 72820 66280 72832 66314
rect 73008 66280 73020 66314
rect 72820 66268 73020 66280
rect 72820 66092 73020 66104
rect 72820 66058 72832 66092
rect 73008 66058 73020 66092
rect 72820 66046 73020 66058
rect 72820 66004 73020 66016
rect 72820 65970 72832 66004
rect 73008 65970 73020 66004
rect 72820 65958 73020 65970
rect 77810 66402 78010 66414
rect 77810 66368 77822 66402
rect 77998 66368 78010 66402
rect 77810 66356 78010 66368
rect 77810 66314 78010 66326
rect 77810 66280 77822 66314
rect 77998 66280 78010 66314
rect 77810 66268 78010 66280
rect 77810 66092 78010 66104
rect 77810 66058 77822 66092
rect 77998 66058 78010 66092
rect 77810 66046 78010 66058
rect 77810 66004 78010 66016
rect 77810 65970 77822 66004
rect 77998 65970 78010 66004
rect 77810 65958 78010 65970
rect 2960 64692 3160 64704
rect 2960 64658 2972 64692
rect 3148 64658 3160 64692
rect 2960 64646 3160 64658
rect 2960 64604 3160 64616
rect 2960 64570 2972 64604
rect 3148 64570 3160 64604
rect 2960 64558 3160 64570
rect 2960 64382 3160 64394
rect 2960 64348 2972 64382
rect 3148 64348 3160 64382
rect 2960 64336 3160 64348
rect 2960 64294 3160 64306
rect 2960 64260 2972 64294
rect 3148 64260 3160 64294
rect 2960 64248 3160 64260
rect 7950 64692 8150 64704
rect 7950 64658 7962 64692
rect 8138 64658 8150 64692
rect 7950 64646 8150 64658
rect 7950 64604 8150 64616
rect 7950 64570 7962 64604
rect 8138 64570 8150 64604
rect 7950 64558 8150 64570
rect 7950 64382 8150 64394
rect 7950 64348 7962 64382
rect 8138 64348 8150 64382
rect 7950 64336 8150 64348
rect 7950 64294 8150 64306
rect 7950 64260 7962 64294
rect 8138 64260 8150 64294
rect 7950 64248 8150 64260
rect 12940 64692 13140 64704
rect 12940 64658 12952 64692
rect 13128 64658 13140 64692
rect 12940 64646 13140 64658
rect 12940 64604 13140 64616
rect 12940 64570 12952 64604
rect 13128 64570 13140 64604
rect 12940 64558 13140 64570
rect 12940 64382 13140 64394
rect 12940 64348 12952 64382
rect 13128 64348 13140 64382
rect 12940 64336 13140 64348
rect 12940 64294 13140 64306
rect 12940 64260 12952 64294
rect 13128 64260 13140 64294
rect 12940 64248 13140 64260
rect 17930 64692 18130 64704
rect 17930 64658 17942 64692
rect 18118 64658 18130 64692
rect 17930 64646 18130 64658
rect 17930 64604 18130 64616
rect 17930 64570 17942 64604
rect 18118 64570 18130 64604
rect 17930 64558 18130 64570
rect 17930 64382 18130 64394
rect 17930 64348 17942 64382
rect 18118 64348 18130 64382
rect 17930 64336 18130 64348
rect 17930 64294 18130 64306
rect 17930 64260 17942 64294
rect 18118 64260 18130 64294
rect 17930 64248 18130 64260
rect 22920 64692 23120 64704
rect 22920 64658 22932 64692
rect 23108 64658 23120 64692
rect 22920 64646 23120 64658
rect 22920 64604 23120 64616
rect 22920 64570 22932 64604
rect 23108 64570 23120 64604
rect 22920 64558 23120 64570
rect 22920 64382 23120 64394
rect 22920 64348 22932 64382
rect 23108 64348 23120 64382
rect 22920 64336 23120 64348
rect 22920 64294 23120 64306
rect 22920 64260 22932 64294
rect 23108 64260 23120 64294
rect 22920 64248 23120 64260
rect 27910 64692 28110 64704
rect 27910 64658 27922 64692
rect 28098 64658 28110 64692
rect 27910 64646 28110 64658
rect 27910 64604 28110 64616
rect 27910 64570 27922 64604
rect 28098 64570 28110 64604
rect 27910 64558 28110 64570
rect 27910 64382 28110 64394
rect 27910 64348 27922 64382
rect 28098 64348 28110 64382
rect 27910 64336 28110 64348
rect 27910 64294 28110 64306
rect 27910 64260 27922 64294
rect 28098 64260 28110 64294
rect 27910 64248 28110 64260
rect 32900 64692 33100 64704
rect 32900 64658 32912 64692
rect 33088 64658 33100 64692
rect 32900 64646 33100 64658
rect 32900 64604 33100 64616
rect 32900 64570 32912 64604
rect 33088 64570 33100 64604
rect 32900 64558 33100 64570
rect 32900 64382 33100 64394
rect 32900 64348 32912 64382
rect 33088 64348 33100 64382
rect 32900 64336 33100 64348
rect 32900 64294 33100 64306
rect 32900 64260 32912 64294
rect 33088 64260 33100 64294
rect 32900 64248 33100 64260
rect 37890 64692 38090 64704
rect 37890 64658 37902 64692
rect 38078 64658 38090 64692
rect 37890 64646 38090 64658
rect 37890 64604 38090 64616
rect 37890 64570 37902 64604
rect 38078 64570 38090 64604
rect 37890 64558 38090 64570
rect 37890 64382 38090 64394
rect 37890 64348 37902 64382
rect 38078 64348 38090 64382
rect 37890 64336 38090 64348
rect 37890 64294 38090 64306
rect 37890 64260 37902 64294
rect 38078 64260 38090 64294
rect 37890 64248 38090 64260
rect 42880 64692 43080 64704
rect 42880 64658 42892 64692
rect 43068 64658 43080 64692
rect 42880 64646 43080 64658
rect 42880 64604 43080 64616
rect 42880 64570 42892 64604
rect 43068 64570 43080 64604
rect 42880 64558 43080 64570
rect 42880 64382 43080 64394
rect 42880 64348 42892 64382
rect 43068 64348 43080 64382
rect 42880 64336 43080 64348
rect 42880 64294 43080 64306
rect 42880 64260 42892 64294
rect 43068 64260 43080 64294
rect 42880 64248 43080 64260
rect 47870 64692 48070 64704
rect 47870 64658 47882 64692
rect 48058 64658 48070 64692
rect 47870 64646 48070 64658
rect 47870 64604 48070 64616
rect 47870 64570 47882 64604
rect 48058 64570 48070 64604
rect 47870 64558 48070 64570
rect 47870 64382 48070 64394
rect 47870 64348 47882 64382
rect 48058 64348 48070 64382
rect 47870 64336 48070 64348
rect 47870 64294 48070 64306
rect 47870 64260 47882 64294
rect 48058 64260 48070 64294
rect 47870 64248 48070 64260
rect 52860 64692 53060 64704
rect 52860 64658 52872 64692
rect 53048 64658 53060 64692
rect 52860 64646 53060 64658
rect 52860 64604 53060 64616
rect 52860 64570 52872 64604
rect 53048 64570 53060 64604
rect 52860 64558 53060 64570
rect 52860 64382 53060 64394
rect 52860 64348 52872 64382
rect 53048 64348 53060 64382
rect 52860 64336 53060 64348
rect 52860 64294 53060 64306
rect 52860 64260 52872 64294
rect 53048 64260 53060 64294
rect 52860 64248 53060 64260
rect 57850 64692 58050 64704
rect 57850 64658 57862 64692
rect 58038 64658 58050 64692
rect 57850 64646 58050 64658
rect 57850 64604 58050 64616
rect 57850 64570 57862 64604
rect 58038 64570 58050 64604
rect 57850 64558 58050 64570
rect 57850 64382 58050 64394
rect 57850 64348 57862 64382
rect 58038 64348 58050 64382
rect 57850 64336 58050 64348
rect 57850 64294 58050 64306
rect 57850 64260 57862 64294
rect 58038 64260 58050 64294
rect 57850 64248 58050 64260
rect 62840 64692 63040 64704
rect 62840 64658 62852 64692
rect 63028 64658 63040 64692
rect 62840 64646 63040 64658
rect 62840 64604 63040 64616
rect 62840 64570 62852 64604
rect 63028 64570 63040 64604
rect 62840 64558 63040 64570
rect 62840 64382 63040 64394
rect 62840 64348 62852 64382
rect 63028 64348 63040 64382
rect 62840 64336 63040 64348
rect 62840 64294 63040 64306
rect 62840 64260 62852 64294
rect 63028 64260 63040 64294
rect 62840 64248 63040 64260
rect 67830 64692 68030 64704
rect 67830 64658 67842 64692
rect 68018 64658 68030 64692
rect 67830 64646 68030 64658
rect 67830 64604 68030 64616
rect 67830 64570 67842 64604
rect 68018 64570 68030 64604
rect 67830 64558 68030 64570
rect 67830 64382 68030 64394
rect 67830 64348 67842 64382
rect 68018 64348 68030 64382
rect 67830 64336 68030 64348
rect 67830 64294 68030 64306
rect 67830 64260 67842 64294
rect 68018 64260 68030 64294
rect 67830 64248 68030 64260
rect 72820 64692 73020 64704
rect 72820 64658 72832 64692
rect 73008 64658 73020 64692
rect 72820 64646 73020 64658
rect 72820 64604 73020 64616
rect 72820 64570 72832 64604
rect 73008 64570 73020 64604
rect 72820 64558 73020 64570
rect 72820 64382 73020 64394
rect 72820 64348 72832 64382
rect 73008 64348 73020 64382
rect 72820 64336 73020 64348
rect 72820 64294 73020 64306
rect 72820 64260 72832 64294
rect 73008 64260 73020 64294
rect 72820 64248 73020 64260
rect 77810 64692 78010 64704
rect 77810 64658 77822 64692
rect 77998 64658 78010 64692
rect 77810 64646 78010 64658
rect 77810 64604 78010 64616
rect 77810 64570 77822 64604
rect 77998 64570 78010 64604
rect 77810 64558 78010 64570
rect 77810 64382 78010 64394
rect 77810 64348 77822 64382
rect 77998 64348 78010 64382
rect 77810 64336 78010 64348
rect 77810 64294 78010 64306
rect 77810 64260 77822 64294
rect 77998 64260 78010 64294
rect 77810 64248 78010 64260
rect 2960 62982 3160 62994
rect 2960 62948 2972 62982
rect 3148 62948 3160 62982
rect 2960 62936 3160 62948
rect 2960 62894 3160 62906
rect 2960 62860 2972 62894
rect 3148 62860 3160 62894
rect 2960 62848 3160 62860
rect 2960 62672 3160 62684
rect 2960 62638 2972 62672
rect 3148 62638 3160 62672
rect 2960 62626 3160 62638
rect 2960 62584 3160 62596
rect 2960 62550 2972 62584
rect 3148 62550 3160 62584
rect 2960 62538 3160 62550
rect 7950 62982 8150 62994
rect 7950 62948 7962 62982
rect 8138 62948 8150 62982
rect 7950 62936 8150 62948
rect 7950 62894 8150 62906
rect 7950 62860 7962 62894
rect 8138 62860 8150 62894
rect 7950 62848 8150 62860
rect 7950 62672 8150 62684
rect 7950 62638 7962 62672
rect 8138 62638 8150 62672
rect 7950 62626 8150 62638
rect 7950 62584 8150 62596
rect 7950 62550 7962 62584
rect 8138 62550 8150 62584
rect 7950 62538 8150 62550
rect 12940 62982 13140 62994
rect 12940 62948 12952 62982
rect 13128 62948 13140 62982
rect 12940 62936 13140 62948
rect 12940 62894 13140 62906
rect 12940 62860 12952 62894
rect 13128 62860 13140 62894
rect 12940 62848 13140 62860
rect 12940 62672 13140 62684
rect 12940 62638 12952 62672
rect 13128 62638 13140 62672
rect 12940 62626 13140 62638
rect 12940 62584 13140 62596
rect 12940 62550 12952 62584
rect 13128 62550 13140 62584
rect 12940 62538 13140 62550
rect 17930 62982 18130 62994
rect 17930 62948 17942 62982
rect 18118 62948 18130 62982
rect 17930 62936 18130 62948
rect 17930 62894 18130 62906
rect 17930 62860 17942 62894
rect 18118 62860 18130 62894
rect 17930 62848 18130 62860
rect 17930 62672 18130 62684
rect 17930 62638 17942 62672
rect 18118 62638 18130 62672
rect 17930 62626 18130 62638
rect 17930 62584 18130 62596
rect 17930 62550 17942 62584
rect 18118 62550 18130 62584
rect 17930 62538 18130 62550
rect 22920 62982 23120 62994
rect 22920 62948 22932 62982
rect 23108 62948 23120 62982
rect 22920 62936 23120 62948
rect 22920 62894 23120 62906
rect 22920 62860 22932 62894
rect 23108 62860 23120 62894
rect 22920 62848 23120 62860
rect 22920 62672 23120 62684
rect 22920 62638 22932 62672
rect 23108 62638 23120 62672
rect 22920 62626 23120 62638
rect 22920 62584 23120 62596
rect 22920 62550 22932 62584
rect 23108 62550 23120 62584
rect 22920 62538 23120 62550
rect 27910 62982 28110 62994
rect 27910 62948 27922 62982
rect 28098 62948 28110 62982
rect 27910 62936 28110 62948
rect 27910 62894 28110 62906
rect 27910 62860 27922 62894
rect 28098 62860 28110 62894
rect 27910 62848 28110 62860
rect 27910 62672 28110 62684
rect 27910 62638 27922 62672
rect 28098 62638 28110 62672
rect 27910 62626 28110 62638
rect 27910 62584 28110 62596
rect 27910 62550 27922 62584
rect 28098 62550 28110 62584
rect 27910 62538 28110 62550
rect 32900 62982 33100 62994
rect 32900 62948 32912 62982
rect 33088 62948 33100 62982
rect 32900 62936 33100 62948
rect 32900 62894 33100 62906
rect 32900 62860 32912 62894
rect 33088 62860 33100 62894
rect 32900 62848 33100 62860
rect 32900 62672 33100 62684
rect 32900 62638 32912 62672
rect 33088 62638 33100 62672
rect 32900 62626 33100 62638
rect 32900 62584 33100 62596
rect 32900 62550 32912 62584
rect 33088 62550 33100 62584
rect 32900 62538 33100 62550
rect 37890 62982 38090 62994
rect 37890 62948 37902 62982
rect 38078 62948 38090 62982
rect 37890 62936 38090 62948
rect 37890 62894 38090 62906
rect 37890 62860 37902 62894
rect 38078 62860 38090 62894
rect 37890 62848 38090 62860
rect 37890 62672 38090 62684
rect 37890 62638 37902 62672
rect 38078 62638 38090 62672
rect 37890 62626 38090 62638
rect 37890 62584 38090 62596
rect 37890 62550 37902 62584
rect 38078 62550 38090 62584
rect 37890 62538 38090 62550
rect 42880 62982 43080 62994
rect 42880 62948 42892 62982
rect 43068 62948 43080 62982
rect 42880 62936 43080 62948
rect 42880 62894 43080 62906
rect 42880 62860 42892 62894
rect 43068 62860 43080 62894
rect 42880 62848 43080 62860
rect 42880 62672 43080 62684
rect 42880 62638 42892 62672
rect 43068 62638 43080 62672
rect 42880 62626 43080 62638
rect 42880 62584 43080 62596
rect 42880 62550 42892 62584
rect 43068 62550 43080 62584
rect 42880 62538 43080 62550
rect 47870 62982 48070 62994
rect 47870 62948 47882 62982
rect 48058 62948 48070 62982
rect 47870 62936 48070 62948
rect 47870 62894 48070 62906
rect 47870 62860 47882 62894
rect 48058 62860 48070 62894
rect 47870 62848 48070 62860
rect 47870 62672 48070 62684
rect 47870 62638 47882 62672
rect 48058 62638 48070 62672
rect 47870 62626 48070 62638
rect 47870 62584 48070 62596
rect 47870 62550 47882 62584
rect 48058 62550 48070 62584
rect 47870 62538 48070 62550
rect 52860 62982 53060 62994
rect 52860 62948 52872 62982
rect 53048 62948 53060 62982
rect 52860 62936 53060 62948
rect 52860 62894 53060 62906
rect 52860 62860 52872 62894
rect 53048 62860 53060 62894
rect 52860 62848 53060 62860
rect 52860 62672 53060 62684
rect 52860 62638 52872 62672
rect 53048 62638 53060 62672
rect 52860 62626 53060 62638
rect 52860 62584 53060 62596
rect 52860 62550 52872 62584
rect 53048 62550 53060 62584
rect 52860 62538 53060 62550
rect 57850 62982 58050 62994
rect 57850 62948 57862 62982
rect 58038 62948 58050 62982
rect 57850 62936 58050 62948
rect 57850 62894 58050 62906
rect 57850 62860 57862 62894
rect 58038 62860 58050 62894
rect 57850 62848 58050 62860
rect 57850 62672 58050 62684
rect 57850 62638 57862 62672
rect 58038 62638 58050 62672
rect 57850 62626 58050 62638
rect 57850 62584 58050 62596
rect 57850 62550 57862 62584
rect 58038 62550 58050 62584
rect 57850 62538 58050 62550
rect 62840 62982 63040 62994
rect 62840 62948 62852 62982
rect 63028 62948 63040 62982
rect 62840 62936 63040 62948
rect 62840 62894 63040 62906
rect 62840 62860 62852 62894
rect 63028 62860 63040 62894
rect 62840 62848 63040 62860
rect 62840 62672 63040 62684
rect 62840 62638 62852 62672
rect 63028 62638 63040 62672
rect 62840 62626 63040 62638
rect 62840 62584 63040 62596
rect 62840 62550 62852 62584
rect 63028 62550 63040 62584
rect 62840 62538 63040 62550
rect 67830 62982 68030 62994
rect 67830 62948 67842 62982
rect 68018 62948 68030 62982
rect 67830 62936 68030 62948
rect 67830 62894 68030 62906
rect 67830 62860 67842 62894
rect 68018 62860 68030 62894
rect 67830 62848 68030 62860
rect 67830 62672 68030 62684
rect 67830 62638 67842 62672
rect 68018 62638 68030 62672
rect 67830 62626 68030 62638
rect 67830 62584 68030 62596
rect 67830 62550 67842 62584
rect 68018 62550 68030 62584
rect 67830 62538 68030 62550
rect 72820 62982 73020 62994
rect 72820 62948 72832 62982
rect 73008 62948 73020 62982
rect 72820 62936 73020 62948
rect 72820 62894 73020 62906
rect 72820 62860 72832 62894
rect 73008 62860 73020 62894
rect 72820 62848 73020 62860
rect 72820 62672 73020 62684
rect 72820 62638 72832 62672
rect 73008 62638 73020 62672
rect 72820 62626 73020 62638
rect 72820 62584 73020 62596
rect 72820 62550 72832 62584
rect 73008 62550 73020 62584
rect 72820 62538 73020 62550
rect 77810 62982 78010 62994
rect 77810 62948 77822 62982
rect 77998 62948 78010 62982
rect 77810 62936 78010 62948
rect 77810 62894 78010 62906
rect 77810 62860 77822 62894
rect 77998 62860 78010 62894
rect 77810 62848 78010 62860
rect 77810 62672 78010 62684
rect 77810 62638 77822 62672
rect 77998 62638 78010 62672
rect 77810 62626 78010 62638
rect 77810 62584 78010 62596
rect 77810 62550 77822 62584
rect 77998 62550 78010 62584
rect 77810 62538 78010 62550
rect 2960 61272 3160 61284
rect 2960 61238 2972 61272
rect 3148 61238 3160 61272
rect 2960 61226 3160 61238
rect 2960 61184 3160 61196
rect 2960 61150 2972 61184
rect 3148 61150 3160 61184
rect 2960 61138 3160 61150
rect 2960 60962 3160 60974
rect 2960 60928 2972 60962
rect 3148 60928 3160 60962
rect 2960 60916 3160 60928
rect 2960 60874 3160 60886
rect 2960 60840 2972 60874
rect 3148 60840 3160 60874
rect 2960 60828 3160 60840
rect 7950 61272 8150 61284
rect 7950 61238 7962 61272
rect 8138 61238 8150 61272
rect 7950 61226 8150 61238
rect 7950 61184 8150 61196
rect 7950 61150 7962 61184
rect 8138 61150 8150 61184
rect 7950 61138 8150 61150
rect 7950 60962 8150 60974
rect 7950 60928 7962 60962
rect 8138 60928 8150 60962
rect 7950 60916 8150 60928
rect 7950 60874 8150 60886
rect 7950 60840 7962 60874
rect 8138 60840 8150 60874
rect 7950 60828 8150 60840
rect 12940 61272 13140 61284
rect 12940 61238 12952 61272
rect 13128 61238 13140 61272
rect 12940 61226 13140 61238
rect 12940 61184 13140 61196
rect 12940 61150 12952 61184
rect 13128 61150 13140 61184
rect 12940 61138 13140 61150
rect 12940 60962 13140 60974
rect 12940 60928 12952 60962
rect 13128 60928 13140 60962
rect 12940 60916 13140 60928
rect 12940 60874 13140 60886
rect 12940 60840 12952 60874
rect 13128 60840 13140 60874
rect 12940 60828 13140 60840
rect 17930 61272 18130 61284
rect 17930 61238 17942 61272
rect 18118 61238 18130 61272
rect 17930 61226 18130 61238
rect 17930 61184 18130 61196
rect 17930 61150 17942 61184
rect 18118 61150 18130 61184
rect 17930 61138 18130 61150
rect 17930 60962 18130 60974
rect 17930 60928 17942 60962
rect 18118 60928 18130 60962
rect 17930 60916 18130 60928
rect 17930 60874 18130 60886
rect 17930 60840 17942 60874
rect 18118 60840 18130 60874
rect 17930 60828 18130 60840
rect 22920 61272 23120 61284
rect 22920 61238 22932 61272
rect 23108 61238 23120 61272
rect 22920 61226 23120 61238
rect 22920 61184 23120 61196
rect 22920 61150 22932 61184
rect 23108 61150 23120 61184
rect 22920 61138 23120 61150
rect 22920 60962 23120 60974
rect 22920 60928 22932 60962
rect 23108 60928 23120 60962
rect 22920 60916 23120 60928
rect 22920 60874 23120 60886
rect 22920 60840 22932 60874
rect 23108 60840 23120 60874
rect 22920 60828 23120 60840
rect 27910 61272 28110 61284
rect 27910 61238 27922 61272
rect 28098 61238 28110 61272
rect 27910 61226 28110 61238
rect 27910 61184 28110 61196
rect 27910 61150 27922 61184
rect 28098 61150 28110 61184
rect 27910 61138 28110 61150
rect 27910 60962 28110 60974
rect 27910 60928 27922 60962
rect 28098 60928 28110 60962
rect 27910 60916 28110 60928
rect 27910 60874 28110 60886
rect 27910 60840 27922 60874
rect 28098 60840 28110 60874
rect 27910 60828 28110 60840
rect 32900 61272 33100 61284
rect 32900 61238 32912 61272
rect 33088 61238 33100 61272
rect 32900 61226 33100 61238
rect 32900 61184 33100 61196
rect 32900 61150 32912 61184
rect 33088 61150 33100 61184
rect 32900 61138 33100 61150
rect 32900 60962 33100 60974
rect 32900 60928 32912 60962
rect 33088 60928 33100 60962
rect 32900 60916 33100 60928
rect 32900 60874 33100 60886
rect 32900 60840 32912 60874
rect 33088 60840 33100 60874
rect 32900 60828 33100 60840
rect 37890 61272 38090 61284
rect 37890 61238 37902 61272
rect 38078 61238 38090 61272
rect 37890 61226 38090 61238
rect 37890 61184 38090 61196
rect 37890 61150 37902 61184
rect 38078 61150 38090 61184
rect 37890 61138 38090 61150
rect 37890 60962 38090 60974
rect 37890 60928 37902 60962
rect 38078 60928 38090 60962
rect 37890 60916 38090 60928
rect 37890 60874 38090 60886
rect 37890 60840 37902 60874
rect 38078 60840 38090 60874
rect 37890 60828 38090 60840
rect 42880 61272 43080 61284
rect 42880 61238 42892 61272
rect 43068 61238 43080 61272
rect 42880 61226 43080 61238
rect 42880 61184 43080 61196
rect 42880 61150 42892 61184
rect 43068 61150 43080 61184
rect 42880 61138 43080 61150
rect 42880 60962 43080 60974
rect 42880 60928 42892 60962
rect 43068 60928 43080 60962
rect 42880 60916 43080 60928
rect 42880 60874 43080 60886
rect 42880 60840 42892 60874
rect 43068 60840 43080 60874
rect 42880 60828 43080 60840
rect 47870 61272 48070 61284
rect 47870 61238 47882 61272
rect 48058 61238 48070 61272
rect 47870 61226 48070 61238
rect 47870 61184 48070 61196
rect 47870 61150 47882 61184
rect 48058 61150 48070 61184
rect 47870 61138 48070 61150
rect 47870 60962 48070 60974
rect 47870 60928 47882 60962
rect 48058 60928 48070 60962
rect 47870 60916 48070 60928
rect 47870 60874 48070 60886
rect 47870 60840 47882 60874
rect 48058 60840 48070 60874
rect 47870 60828 48070 60840
rect 52860 61272 53060 61284
rect 52860 61238 52872 61272
rect 53048 61238 53060 61272
rect 52860 61226 53060 61238
rect 52860 61184 53060 61196
rect 52860 61150 52872 61184
rect 53048 61150 53060 61184
rect 52860 61138 53060 61150
rect 52860 60962 53060 60974
rect 52860 60928 52872 60962
rect 53048 60928 53060 60962
rect 52860 60916 53060 60928
rect 52860 60874 53060 60886
rect 52860 60840 52872 60874
rect 53048 60840 53060 60874
rect 52860 60828 53060 60840
rect 57850 61272 58050 61284
rect 57850 61238 57862 61272
rect 58038 61238 58050 61272
rect 57850 61226 58050 61238
rect 57850 61184 58050 61196
rect 57850 61150 57862 61184
rect 58038 61150 58050 61184
rect 57850 61138 58050 61150
rect 57850 60962 58050 60974
rect 57850 60928 57862 60962
rect 58038 60928 58050 60962
rect 57850 60916 58050 60928
rect 57850 60874 58050 60886
rect 57850 60840 57862 60874
rect 58038 60840 58050 60874
rect 57850 60828 58050 60840
rect 62840 61272 63040 61284
rect 62840 61238 62852 61272
rect 63028 61238 63040 61272
rect 62840 61226 63040 61238
rect 62840 61184 63040 61196
rect 62840 61150 62852 61184
rect 63028 61150 63040 61184
rect 62840 61138 63040 61150
rect 62840 60962 63040 60974
rect 62840 60928 62852 60962
rect 63028 60928 63040 60962
rect 62840 60916 63040 60928
rect 62840 60874 63040 60886
rect 62840 60840 62852 60874
rect 63028 60840 63040 60874
rect 62840 60828 63040 60840
rect 67830 61272 68030 61284
rect 67830 61238 67842 61272
rect 68018 61238 68030 61272
rect 67830 61226 68030 61238
rect 67830 61184 68030 61196
rect 67830 61150 67842 61184
rect 68018 61150 68030 61184
rect 67830 61138 68030 61150
rect 67830 60962 68030 60974
rect 67830 60928 67842 60962
rect 68018 60928 68030 60962
rect 67830 60916 68030 60928
rect 67830 60874 68030 60886
rect 67830 60840 67842 60874
rect 68018 60840 68030 60874
rect 67830 60828 68030 60840
rect 72820 61272 73020 61284
rect 72820 61238 72832 61272
rect 73008 61238 73020 61272
rect 72820 61226 73020 61238
rect 72820 61184 73020 61196
rect 72820 61150 72832 61184
rect 73008 61150 73020 61184
rect 72820 61138 73020 61150
rect 72820 60962 73020 60974
rect 72820 60928 72832 60962
rect 73008 60928 73020 60962
rect 72820 60916 73020 60928
rect 72820 60874 73020 60886
rect 72820 60840 72832 60874
rect 73008 60840 73020 60874
rect 72820 60828 73020 60840
rect 77810 61272 78010 61284
rect 77810 61238 77822 61272
rect 77998 61238 78010 61272
rect 77810 61226 78010 61238
rect 77810 61184 78010 61196
rect 77810 61150 77822 61184
rect 77998 61150 78010 61184
rect 77810 61138 78010 61150
rect 77810 60962 78010 60974
rect 77810 60928 77822 60962
rect 77998 60928 78010 60962
rect 77810 60916 78010 60928
rect 77810 60874 78010 60886
rect 77810 60840 77822 60874
rect 77998 60840 78010 60874
rect 77810 60828 78010 60840
rect 2960 59562 3160 59574
rect 2960 59528 2972 59562
rect 3148 59528 3160 59562
rect 2960 59516 3160 59528
rect 2960 59474 3160 59486
rect 2960 59440 2972 59474
rect 3148 59440 3160 59474
rect 2960 59428 3160 59440
rect 2960 59252 3160 59264
rect 2960 59218 2972 59252
rect 3148 59218 3160 59252
rect 2960 59206 3160 59218
rect 2960 59164 3160 59176
rect 2960 59130 2972 59164
rect 3148 59130 3160 59164
rect 2960 59118 3160 59130
rect 7950 59562 8150 59574
rect 7950 59528 7962 59562
rect 8138 59528 8150 59562
rect 7950 59516 8150 59528
rect 7950 59474 8150 59486
rect 7950 59440 7962 59474
rect 8138 59440 8150 59474
rect 7950 59428 8150 59440
rect 7950 59252 8150 59264
rect 7950 59218 7962 59252
rect 8138 59218 8150 59252
rect 7950 59206 8150 59218
rect 7950 59164 8150 59176
rect 7950 59130 7962 59164
rect 8138 59130 8150 59164
rect 7950 59118 8150 59130
rect 12940 59562 13140 59574
rect 12940 59528 12952 59562
rect 13128 59528 13140 59562
rect 12940 59516 13140 59528
rect 12940 59474 13140 59486
rect 12940 59440 12952 59474
rect 13128 59440 13140 59474
rect 12940 59428 13140 59440
rect 12940 59252 13140 59264
rect 12940 59218 12952 59252
rect 13128 59218 13140 59252
rect 12940 59206 13140 59218
rect 12940 59164 13140 59176
rect 12940 59130 12952 59164
rect 13128 59130 13140 59164
rect 12940 59118 13140 59130
rect 17930 59562 18130 59574
rect 17930 59528 17942 59562
rect 18118 59528 18130 59562
rect 17930 59516 18130 59528
rect 17930 59474 18130 59486
rect 17930 59440 17942 59474
rect 18118 59440 18130 59474
rect 17930 59428 18130 59440
rect 17930 59252 18130 59264
rect 17930 59218 17942 59252
rect 18118 59218 18130 59252
rect 17930 59206 18130 59218
rect 17930 59164 18130 59176
rect 17930 59130 17942 59164
rect 18118 59130 18130 59164
rect 17930 59118 18130 59130
rect 22920 59562 23120 59574
rect 22920 59528 22932 59562
rect 23108 59528 23120 59562
rect 22920 59516 23120 59528
rect 22920 59474 23120 59486
rect 22920 59440 22932 59474
rect 23108 59440 23120 59474
rect 22920 59428 23120 59440
rect 22920 59252 23120 59264
rect 22920 59218 22932 59252
rect 23108 59218 23120 59252
rect 22920 59206 23120 59218
rect 22920 59164 23120 59176
rect 22920 59130 22932 59164
rect 23108 59130 23120 59164
rect 22920 59118 23120 59130
rect 27910 59562 28110 59574
rect 27910 59528 27922 59562
rect 28098 59528 28110 59562
rect 27910 59516 28110 59528
rect 27910 59474 28110 59486
rect 27910 59440 27922 59474
rect 28098 59440 28110 59474
rect 27910 59428 28110 59440
rect 27910 59252 28110 59264
rect 27910 59218 27922 59252
rect 28098 59218 28110 59252
rect 27910 59206 28110 59218
rect 27910 59164 28110 59176
rect 27910 59130 27922 59164
rect 28098 59130 28110 59164
rect 27910 59118 28110 59130
rect 32900 59562 33100 59574
rect 32900 59528 32912 59562
rect 33088 59528 33100 59562
rect 32900 59516 33100 59528
rect 32900 59474 33100 59486
rect 32900 59440 32912 59474
rect 33088 59440 33100 59474
rect 32900 59428 33100 59440
rect 32900 59252 33100 59264
rect 32900 59218 32912 59252
rect 33088 59218 33100 59252
rect 32900 59206 33100 59218
rect 32900 59164 33100 59176
rect 32900 59130 32912 59164
rect 33088 59130 33100 59164
rect 32900 59118 33100 59130
rect 37890 59562 38090 59574
rect 37890 59528 37902 59562
rect 38078 59528 38090 59562
rect 37890 59516 38090 59528
rect 37890 59474 38090 59486
rect 37890 59440 37902 59474
rect 38078 59440 38090 59474
rect 37890 59428 38090 59440
rect 37890 59252 38090 59264
rect 37890 59218 37902 59252
rect 38078 59218 38090 59252
rect 37890 59206 38090 59218
rect 37890 59164 38090 59176
rect 37890 59130 37902 59164
rect 38078 59130 38090 59164
rect 37890 59118 38090 59130
rect 42880 59562 43080 59574
rect 42880 59528 42892 59562
rect 43068 59528 43080 59562
rect 42880 59516 43080 59528
rect 42880 59474 43080 59486
rect 42880 59440 42892 59474
rect 43068 59440 43080 59474
rect 42880 59428 43080 59440
rect 42880 59252 43080 59264
rect 42880 59218 42892 59252
rect 43068 59218 43080 59252
rect 42880 59206 43080 59218
rect 42880 59164 43080 59176
rect 42880 59130 42892 59164
rect 43068 59130 43080 59164
rect 42880 59118 43080 59130
rect 47870 59562 48070 59574
rect 47870 59528 47882 59562
rect 48058 59528 48070 59562
rect 47870 59516 48070 59528
rect 47870 59474 48070 59486
rect 47870 59440 47882 59474
rect 48058 59440 48070 59474
rect 47870 59428 48070 59440
rect 47870 59252 48070 59264
rect 47870 59218 47882 59252
rect 48058 59218 48070 59252
rect 47870 59206 48070 59218
rect 47870 59164 48070 59176
rect 47870 59130 47882 59164
rect 48058 59130 48070 59164
rect 47870 59118 48070 59130
rect 52860 59562 53060 59574
rect 52860 59528 52872 59562
rect 53048 59528 53060 59562
rect 52860 59516 53060 59528
rect 52860 59474 53060 59486
rect 52860 59440 52872 59474
rect 53048 59440 53060 59474
rect 52860 59428 53060 59440
rect 52860 59252 53060 59264
rect 52860 59218 52872 59252
rect 53048 59218 53060 59252
rect 52860 59206 53060 59218
rect 52860 59164 53060 59176
rect 52860 59130 52872 59164
rect 53048 59130 53060 59164
rect 52860 59118 53060 59130
rect 57850 59562 58050 59574
rect 57850 59528 57862 59562
rect 58038 59528 58050 59562
rect 57850 59516 58050 59528
rect 57850 59474 58050 59486
rect 57850 59440 57862 59474
rect 58038 59440 58050 59474
rect 57850 59428 58050 59440
rect 57850 59252 58050 59264
rect 57850 59218 57862 59252
rect 58038 59218 58050 59252
rect 57850 59206 58050 59218
rect 57850 59164 58050 59176
rect 57850 59130 57862 59164
rect 58038 59130 58050 59164
rect 57850 59118 58050 59130
rect 62840 59562 63040 59574
rect 62840 59528 62852 59562
rect 63028 59528 63040 59562
rect 62840 59516 63040 59528
rect 62840 59474 63040 59486
rect 62840 59440 62852 59474
rect 63028 59440 63040 59474
rect 62840 59428 63040 59440
rect 62840 59252 63040 59264
rect 62840 59218 62852 59252
rect 63028 59218 63040 59252
rect 62840 59206 63040 59218
rect 62840 59164 63040 59176
rect 62840 59130 62852 59164
rect 63028 59130 63040 59164
rect 62840 59118 63040 59130
rect 67830 59562 68030 59574
rect 67830 59528 67842 59562
rect 68018 59528 68030 59562
rect 67830 59516 68030 59528
rect 67830 59474 68030 59486
rect 67830 59440 67842 59474
rect 68018 59440 68030 59474
rect 67830 59428 68030 59440
rect 67830 59252 68030 59264
rect 67830 59218 67842 59252
rect 68018 59218 68030 59252
rect 67830 59206 68030 59218
rect 67830 59164 68030 59176
rect 67830 59130 67842 59164
rect 68018 59130 68030 59164
rect 67830 59118 68030 59130
rect 72820 59562 73020 59574
rect 72820 59528 72832 59562
rect 73008 59528 73020 59562
rect 72820 59516 73020 59528
rect 72820 59474 73020 59486
rect 72820 59440 72832 59474
rect 73008 59440 73020 59474
rect 72820 59428 73020 59440
rect 72820 59252 73020 59264
rect 72820 59218 72832 59252
rect 73008 59218 73020 59252
rect 72820 59206 73020 59218
rect 72820 59164 73020 59176
rect 72820 59130 72832 59164
rect 73008 59130 73020 59164
rect 72820 59118 73020 59130
rect 77810 59562 78010 59574
rect 77810 59528 77822 59562
rect 77998 59528 78010 59562
rect 77810 59516 78010 59528
rect 77810 59474 78010 59486
rect 77810 59440 77822 59474
rect 77998 59440 78010 59474
rect 77810 59428 78010 59440
rect 77810 59252 78010 59264
rect 77810 59218 77822 59252
rect 77998 59218 78010 59252
rect 77810 59206 78010 59218
rect 77810 59164 78010 59176
rect 77810 59130 77822 59164
rect 77998 59130 78010 59164
rect 77810 59118 78010 59130
rect 2960 57852 3160 57864
rect 2960 57818 2972 57852
rect 3148 57818 3160 57852
rect 2960 57806 3160 57818
rect 2960 57764 3160 57776
rect 2960 57730 2972 57764
rect 3148 57730 3160 57764
rect 2960 57718 3160 57730
rect 2960 57542 3160 57554
rect 2960 57508 2972 57542
rect 3148 57508 3160 57542
rect 2960 57496 3160 57508
rect 2960 57454 3160 57466
rect 2960 57420 2972 57454
rect 3148 57420 3160 57454
rect 2960 57408 3160 57420
rect 7950 57852 8150 57864
rect 7950 57818 7962 57852
rect 8138 57818 8150 57852
rect 7950 57806 8150 57818
rect 7950 57764 8150 57776
rect 7950 57730 7962 57764
rect 8138 57730 8150 57764
rect 7950 57718 8150 57730
rect 7950 57542 8150 57554
rect 7950 57508 7962 57542
rect 8138 57508 8150 57542
rect 7950 57496 8150 57508
rect 7950 57454 8150 57466
rect 7950 57420 7962 57454
rect 8138 57420 8150 57454
rect 7950 57408 8150 57420
rect 12940 57852 13140 57864
rect 12940 57818 12952 57852
rect 13128 57818 13140 57852
rect 12940 57806 13140 57818
rect 12940 57764 13140 57776
rect 12940 57730 12952 57764
rect 13128 57730 13140 57764
rect 12940 57718 13140 57730
rect 12940 57542 13140 57554
rect 12940 57508 12952 57542
rect 13128 57508 13140 57542
rect 12940 57496 13140 57508
rect 12940 57454 13140 57466
rect 12940 57420 12952 57454
rect 13128 57420 13140 57454
rect 12940 57408 13140 57420
rect 17930 57852 18130 57864
rect 17930 57818 17942 57852
rect 18118 57818 18130 57852
rect 17930 57806 18130 57818
rect 17930 57764 18130 57776
rect 17930 57730 17942 57764
rect 18118 57730 18130 57764
rect 17930 57718 18130 57730
rect 17930 57542 18130 57554
rect 17930 57508 17942 57542
rect 18118 57508 18130 57542
rect 17930 57496 18130 57508
rect 17930 57454 18130 57466
rect 17930 57420 17942 57454
rect 18118 57420 18130 57454
rect 17930 57408 18130 57420
rect 22920 57852 23120 57864
rect 22920 57818 22932 57852
rect 23108 57818 23120 57852
rect 22920 57806 23120 57818
rect 22920 57764 23120 57776
rect 22920 57730 22932 57764
rect 23108 57730 23120 57764
rect 22920 57718 23120 57730
rect 22920 57542 23120 57554
rect 22920 57508 22932 57542
rect 23108 57508 23120 57542
rect 22920 57496 23120 57508
rect 22920 57454 23120 57466
rect 22920 57420 22932 57454
rect 23108 57420 23120 57454
rect 22920 57408 23120 57420
rect 27910 57852 28110 57864
rect 27910 57818 27922 57852
rect 28098 57818 28110 57852
rect 27910 57806 28110 57818
rect 27910 57764 28110 57776
rect 27910 57730 27922 57764
rect 28098 57730 28110 57764
rect 27910 57718 28110 57730
rect 27910 57542 28110 57554
rect 27910 57508 27922 57542
rect 28098 57508 28110 57542
rect 27910 57496 28110 57508
rect 27910 57454 28110 57466
rect 27910 57420 27922 57454
rect 28098 57420 28110 57454
rect 27910 57408 28110 57420
rect 32900 57852 33100 57864
rect 32900 57818 32912 57852
rect 33088 57818 33100 57852
rect 32900 57806 33100 57818
rect 32900 57764 33100 57776
rect 32900 57730 32912 57764
rect 33088 57730 33100 57764
rect 32900 57718 33100 57730
rect 32900 57542 33100 57554
rect 32900 57508 32912 57542
rect 33088 57508 33100 57542
rect 32900 57496 33100 57508
rect 32900 57454 33100 57466
rect 32900 57420 32912 57454
rect 33088 57420 33100 57454
rect 32900 57408 33100 57420
rect 37890 57852 38090 57864
rect 37890 57818 37902 57852
rect 38078 57818 38090 57852
rect 37890 57806 38090 57818
rect 37890 57764 38090 57776
rect 37890 57730 37902 57764
rect 38078 57730 38090 57764
rect 37890 57718 38090 57730
rect 37890 57542 38090 57554
rect 37890 57508 37902 57542
rect 38078 57508 38090 57542
rect 37890 57496 38090 57508
rect 37890 57454 38090 57466
rect 37890 57420 37902 57454
rect 38078 57420 38090 57454
rect 37890 57408 38090 57420
rect 42880 57852 43080 57864
rect 42880 57818 42892 57852
rect 43068 57818 43080 57852
rect 42880 57806 43080 57818
rect 42880 57764 43080 57776
rect 42880 57730 42892 57764
rect 43068 57730 43080 57764
rect 42880 57718 43080 57730
rect 42880 57542 43080 57554
rect 42880 57508 42892 57542
rect 43068 57508 43080 57542
rect 42880 57496 43080 57508
rect 42880 57454 43080 57466
rect 42880 57420 42892 57454
rect 43068 57420 43080 57454
rect 42880 57408 43080 57420
rect 47870 57852 48070 57864
rect 47870 57818 47882 57852
rect 48058 57818 48070 57852
rect 47870 57806 48070 57818
rect 47870 57764 48070 57776
rect 47870 57730 47882 57764
rect 48058 57730 48070 57764
rect 47870 57718 48070 57730
rect 47870 57542 48070 57554
rect 47870 57508 47882 57542
rect 48058 57508 48070 57542
rect 47870 57496 48070 57508
rect 47870 57454 48070 57466
rect 47870 57420 47882 57454
rect 48058 57420 48070 57454
rect 47870 57408 48070 57420
rect 52860 57852 53060 57864
rect 52860 57818 52872 57852
rect 53048 57818 53060 57852
rect 52860 57806 53060 57818
rect 52860 57764 53060 57776
rect 52860 57730 52872 57764
rect 53048 57730 53060 57764
rect 52860 57718 53060 57730
rect 52860 57542 53060 57554
rect 52860 57508 52872 57542
rect 53048 57508 53060 57542
rect 52860 57496 53060 57508
rect 52860 57454 53060 57466
rect 52860 57420 52872 57454
rect 53048 57420 53060 57454
rect 52860 57408 53060 57420
rect 57850 57852 58050 57864
rect 57850 57818 57862 57852
rect 58038 57818 58050 57852
rect 57850 57806 58050 57818
rect 57850 57764 58050 57776
rect 57850 57730 57862 57764
rect 58038 57730 58050 57764
rect 57850 57718 58050 57730
rect 57850 57542 58050 57554
rect 57850 57508 57862 57542
rect 58038 57508 58050 57542
rect 57850 57496 58050 57508
rect 57850 57454 58050 57466
rect 57850 57420 57862 57454
rect 58038 57420 58050 57454
rect 57850 57408 58050 57420
rect 62840 57852 63040 57864
rect 62840 57818 62852 57852
rect 63028 57818 63040 57852
rect 62840 57806 63040 57818
rect 62840 57764 63040 57776
rect 62840 57730 62852 57764
rect 63028 57730 63040 57764
rect 62840 57718 63040 57730
rect 62840 57542 63040 57554
rect 62840 57508 62852 57542
rect 63028 57508 63040 57542
rect 62840 57496 63040 57508
rect 62840 57454 63040 57466
rect 62840 57420 62852 57454
rect 63028 57420 63040 57454
rect 62840 57408 63040 57420
rect 67830 57852 68030 57864
rect 67830 57818 67842 57852
rect 68018 57818 68030 57852
rect 67830 57806 68030 57818
rect 67830 57764 68030 57776
rect 67830 57730 67842 57764
rect 68018 57730 68030 57764
rect 67830 57718 68030 57730
rect 67830 57542 68030 57554
rect 67830 57508 67842 57542
rect 68018 57508 68030 57542
rect 67830 57496 68030 57508
rect 67830 57454 68030 57466
rect 67830 57420 67842 57454
rect 68018 57420 68030 57454
rect 67830 57408 68030 57420
rect 72820 57852 73020 57864
rect 72820 57818 72832 57852
rect 73008 57818 73020 57852
rect 72820 57806 73020 57818
rect 72820 57764 73020 57776
rect 72820 57730 72832 57764
rect 73008 57730 73020 57764
rect 72820 57718 73020 57730
rect 72820 57542 73020 57554
rect 72820 57508 72832 57542
rect 73008 57508 73020 57542
rect 72820 57496 73020 57508
rect 72820 57454 73020 57466
rect 72820 57420 72832 57454
rect 73008 57420 73020 57454
rect 72820 57408 73020 57420
rect 77810 57852 78010 57864
rect 77810 57818 77822 57852
rect 77998 57818 78010 57852
rect 77810 57806 78010 57818
rect 77810 57764 78010 57776
rect 77810 57730 77822 57764
rect 77998 57730 78010 57764
rect 77810 57718 78010 57730
rect 77810 57542 78010 57554
rect 77810 57508 77822 57542
rect 77998 57508 78010 57542
rect 77810 57496 78010 57508
rect 77810 57454 78010 57466
rect 77810 57420 77822 57454
rect 77998 57420 78010 57454
rect 77810 57408 78010 57420
rect 2960 56142 3160 56154
rect 2960 56108 2972 56142
rect 3148 56108 3160 56142
rect 2960 56096 3160 56108
rect 2960 56054 3160 56066
rect 2960 56020 2972 56054
rect 3148 56020 3160 56054
rect 2960 56008 3160 56020
rect 2960 55832 3160 55844
rect 2960 55798 2972 55832
rect 3148 55798 3160 55832
rect 2960 55786 3160 55798
rect 2960 55744 3160 55756
rect 2960 55710 2972 55744
rect 3148 55710 3160 55744
rect 2960 55698 3160 55710
rect 7950 56142 8150 56154
rect 7950 56108 7962 56142
rect 8138 56108 8150 56142
rect 7950 56096 8150 56108
rect 7950 56054 8150 56066
rect 7950 56020 7962 56054
rect 8138 56020 8150 56054
rect 7950 56008 8150 56020
rect 7950 55832 8150 55844
rect 7950 55798 7962 55832
rect 8138 55798 8150 55832
rect 7950 55786 8150 55798
rect 7950 55744 8150 55756
rect 7950 55710 7962 55744
rect 8138 55710 8150 55744
rect 7950 55698 8150 55710
rect 12940 56142 13140 56154
rect 12940 56108 12952 56142
rect 13128 56108 13140 56142
rect 12940 56096 13140 56108
rect 12940 56054 13140 56066
rect 12940 56020 12952 56054
rect 13128 56020 13140 56054
rect 12940 56008 13140 56020
rect 12940 55832 13140 55844
rect 12940 55798 12952 55832
rect 13128 55798 13140 55832
rect 12940 55786 13140 55798
rect 12940 55744 13140 55756
rect 12940 55710 12952 55744
rect 13128 55710 13140 55744
rect 12940 55698 13140 55710
rect 17930 56142 18130 56154
rect 17930 56108 17942 56142
rect 18118 56108 18130 56142
rect 17930 56096 18130 56108
rect 17930 56054 18130 56066
rect 17930 56020 17942 56054
rect 18118 56020 18130 56054
rect 17930 56008 18130 56020
rect 17930 55832 18130 55844
rect 17930 55798 17942 55832
rect 18118 55798 18130 55832
rect 17930 55786 18130 55798
rect 17930 55744 18130 55756
rect 17930 55710 17942 55744
rect 18118 55710 18130 55744
rect 17930 55698 18130 55710
rect 22920 56142 23120 56154
rect 22920 56108 22932 56142
rect 23108 56108 23120 56142
rect 22920 56096 23120 56108
rect 22920 56054 23120 56066
rect 22920 56020 22932 56054
rect 23108 56020 23120 56054
rect 22920 56008 23120 56020
rect 22920 55832 23120 55844
rect 22920 55798 22932 55832
rect 23108 55798 23120 55832
rect 22920 55786 23120 55798
rect 22920 55744 23120 55756
rect 22920 55710 22932 55744
rect 23108 55710 23120 55744
rect 22920 55698 23120 55710
rect 27910 56142 28110 56154
rect 27910 56108 27922 56142
rect 28098 56108 28110 56142
rect 27910 56096 28110 56108
rect 27910 56054 28110 56066
rect 27910 56020 27922 56054
rect 28098 56020 28110 56054
rect 27910 56008 28110 56020
rect 27910 55832 28110 55844
rect 27910 55798 27922 55832
rect 28098 55798 28110 55832
rect 27910 55786 28110 55798
rect 27910 55744 28110 55756
rect 27910 55710 27922 55744
rect 28098 55710 28110 55744
rect 27910 55698 28110 55710
rect 32900 56142 33100 56154
rect 32900 56108 32912 56142
rect 33088 56108 33100 56142
rect 32900 56096 33100 56108
rect 32900 56054 33100 56066
rect 32900 56020 32912 56054
rect 33088 56020 33100 56054
rect 32900 56008 33100 56020
rect 32900 55832 33100 55844
rect 32900 55798 32912 55832
rect 33088 55798 33100 55832
rect 32900 55786 33100 55798
rect 32900 55744 33100 55756
rect 32900 55710 32912 55744
rect 33088 55710 33100 55744
rect 32900 55698 33100 55710
rect 37890 56142 38090 56154
rect 37890 56108 37902 56142
rect 38078 56108 38090 56142
rect 37890 56096 38090 56108
rect 37890 56054 38090 56066
rect 37890 56020 37902 56054
rect 38078 56020 38090 56054
rect 37890 56008 38090 56020
rect 37890 55832 38090 55844
rect 37890 55798 37902 55832
rect 38078 55798 38090 55832
rect 37890 55786 38090 55798
rect 37890 55744 38090 55756
rect 37890 55710 37902 55744
rect 38078 55710 38090 55744
rect 37890 55698 38090 55710
rect 42880 56142 43080 56154
rect 42880 56108 42892 56142
rect 43068 56108 43080 56142
rect 42880 56096 43080 56108
rect 42880 56054 43080 56066
rect 42880 56020 42892 56054
rect 43068 56020 43080 56054
rect 42880 56008 43080 56020
rect 42880 55832 43080 55844
rect 42880 55798 42892 55832
rect 43068 55798 43080 55832
rect 42880 55786 43080 55798
rect 42880 55744 43080 55756
rect 42880 55710 42892 55744
rect 43068 55710 43080 55744
rect 42880 55698 43080 55710
rect 47870 56142 48070 56154
rect 47870 56108 47882 56142
rect 48058 56108 48070 56142
rect 47870 56096 48070 56108
rect 47870 56054 48070 56066
rect 47870 56020 47882 56054
rect 48058 56020 48070 56054
rect 47870 56008 48070 56020
rect 47870 55832 48070 55844
rect 47870 55798 47882 55832
rect 48058 55798 48070 55832
rect 47870 55786 48070 55798
rect 47870 55744 48070 55756
rect 47870 55710 47882 55744
rect 48058 55710 48070 55744
rect 47870 55698 48070 55710
rect 52860 56142 53060 56154
rect 52860 56108 52872 56142
rect 53048 56108 53060 56142
rect 52860 56096 53060 56108
rect 52860 56054 53060 56066
rect 52860 56020 52872 56054
rect 53048 56020 53060 56054
rect 52860 56008 53060 56020
rect 52860 55832 53060 55844
rect 52860 55798 52872 55832
rect 53048 55798 53060 55832
rect 52860 55786 53060 55798
rect 52860 55744 53060 55756
rect 52860 55710 52872 55744
rect 53048 55710 53060 55744
rect 52860 55698 53060 55710
rect 57850 56142 58050 56154
rect 57850 56108 57862 56142
rect 58038 56108 58050 56142
rect 57850 56096 58050 56108
rect 57850 56054 58050 56066
rect 57850 56020 57862 56054
rect 58038 56020 58050 56054
rect 57850 56008 58050 56020
rect 57850 55832 58050 55844
rect 57850 55798 57862 55832
rect 58038 55798 58050 55832
rect 57850 55786 58050 55798
rect 57850 55744 58050 55756
rect 57850 55710 57862 55744
rect 58038 55710 58050 55744
rect 57850 55698 58050 55710
rect 62840 56142 63040 56154
rect 62840 56108 62852 56142
rect 63028 56108 63040 56142
rect 62840 56096 63040 56108
rect 62840 56054 63040 56066
rect 62840 56020 62852 56054
rect 63028 56020 63040 56054
rect 62840 56008 63040 56020
rect 62840 55832 63040 55844
rect 62840 55798 62852 55832
rect 63028 55798 63040 55832
rect 62840 55786 63040 55798
rect 62840 55744 63040 55756
rect 62840 55710 62852 55744
rect 63028 55710 63040 55744
rect 62840 55698 63040 55710
rect 67830 56142 68030 56154
rect 67830 56108 67842 56142
rect 68018 56108 68030 56142
rect 67830 56096 68030 56108
rect 67830 56054 68030 56066
rect 67830 56020 67842 56054
rect 68018 56020 68030 56054
rect 67830 56008 68030 56020
rect 67830 55832 68030 55844
rect 67830 55798 67842 55832
rect 68018 55798 68030 55832
rect 67830 55786 68030 55798
rect 67830 55744 68030 55756
rect 67830 55710 67842 55744
rect 68018 55710 68030 55744
rect 67830 55698 68030 55710
rect 72820 56142 73020 56154
rect 72820 56108 72832 56142
rect 73008 56108 73020 56142
rect 72820 56096 73020 56108
rect 72820 56054 73020 56066
rect 72820 56020 72832 56054
rect 73008 56020 73020 56054
rect 72820 56008 73020 56020
rect 72820 55832 73020 55844
rect 72820 55798 72832 55832
rect 73008 55798 73020 55832
rect 72820 55786 73020 55798
rect 72820 55744 73020 55756
rect 72820 55710 72832 55744
rect 73008 55710 73020 55744
rect 72820 55698 73020 55710
rect 77810 56142 78010 56154
rect 77810 56108 77822 56142
rect 77998 56108 78010 56142
rect 77810 56096 78010 56108
rect 77810 56054 78010 56066
rect 77810 56020 77822 56054
rect 77998 56020 78010 56054
rect 77810 56008 78010 56020
rect 77810 55832 78010 55844
rect 77810 55798 77822 55832
rect 77998 55798 78010 55832
rect 77810 55786 78010 55798
rect 77810 55744 78010 55756
rect 77810 55710 77822 55744
rect 77998 55710 78010 55744
rect 77810 55698 78010 55710
rect 2960 54432 3160 54444
rect 2960 54398 2972 54432
rect 3148 54398 3160 54432
rect 2960 54386 3160 54398
rect 2960 54344 3160 54356
rect 2960 54310 2972 54344
rect 3148 54310 3160 54344
rect 2960 54298 3160 54310
rect 2960 54122 3160 54134
rect 2960 54088 2972 54122
rect 3148 54088 3160 54122
rect 2960 54076 3160 54088
rect 2960 54034 3160 54046
rect 2960 54000 2972 54034
rect 3148 54000 3160 54034
rect 2960 53988 3160 54000
rect 7950 54432 8150 54444
rect 7950 54398 7962 54432
rect 8138 54398 8150 54432
rect 7950 54386 8150 54398
rect 7950 54344 8150 54356
rect 7950 54310 7962 54344
rect 8138 54310 8150 54344
rect 7950 54298 8150 54310
rect 7950 54122 8150 54134
rect 7950 54088 7962 54122
rect 8138 54088 8150 54122
rect 7950 54076 8150 54088
rect 7950 54034 8150 54046
rect 7950 54000 7962 54034
rect 8138 54000 8150 54034
rect 7950 53988 8150 54000
rect 12940 54432 13140 54444
rect 12940 54398 12952 54432
rect 13128 54398 13140 54432
rect 12940 54386 13140 54398
rect 12940 54344 13140 54356
rect 12940 54310 12952 54344
rect 13128 54310 13140 54344
rect 12940 54298 13140 54310
rect 12940 54122 13140 54134
rect 12940 54088 12952 54122
rect 13128 54088 13140 54122
rect 12940 54076 13140 54088
rect 12940 54034 13140 54046
rect 12940 54000 12952 54034
rect 13128 54000 13140 54034
rect 12940 53988 13140 54000
rect 17930 54432 18130 54444
rect 17930 54398 17942 54432
rect 18118 54398 18130 54432
rect 17930 54386 18130 54398
rect 17930 54344 18130 54356
rect 17930 54310 17942 54344
rect 18118 54310 18130 54344
rect 17930 54298 18130 54310
rect 17930 54122 18130 54134
rect 17930 54088 17942 54122
rect 18118 54088 18130 54122
rect 17930 54076 18130 54088
rect 17930 54034 18130 54046
rect 17930 54000 17942 54034
rect 18118 54000 18130 54034
rect 17930 53988 18130 54000
rect 22920 54432 23120 54444
rect 22920 54398 22932 54432
rect 23108 54398 23120 54432
rect 22920 54386 23120 54398
rect 22920 54344 23120 54356
rect 22920 54310 22932 54344
rect 23108 54310 23120 54344
rect 22920 54298 23120 54310
rect 22920 54122 23120 54134
rect 22920 54088 22932 54122
rect 23108 54088 23120 54122
rect 22920 54076 23120 54088
rect 22920 54034 23120 54046
rect 22920 54000 22932 54034
rect 23108 54000 23120 54034
rect 22920 53988 23120 54000
rect 27910 54432 28110 54444
rect 27910 54398 27922 54432
rect 28098 54398 28110 54432
rect 27910 54386 28110 54398
rect 27910 54344 28110 54356
rect 27910 54310 27922 54344
rect 28098 54310 28110 54344
rect 27910 54298 28110 54310
rect 27910 54122 28110 54134
rect 27910 54088 27922 54122
rect 28098 54088 28110 54122
rect 27910 54076 28110 54088
rect 27910 54034 28110 54046
rect 27910 54000 27922 54034
rect 28098 54000 28110 54034
rect 27910 53988 28110 54000
rect 32900 54432 33100 54444
rect 32900 54398 32912 54432
rect 33088 54398 33100 54432
rect 32900 54386 33100 54398
rect 32900 54344 33100 54356
rect 32900 54310 32912 54344
rect 33088 54310 33100 54344
rect 32900 54298 33100 54310
rect 32900 54122 33100 54134
rect 32900 54088 32912 54122
rect 33088 54088 33100 54122
rect 32900 54076 33100 54088
rect 32900 54034 33100 54046
rect 32900 54000 32912 54034
rect 33088 54000 33100 54034
rect 32900 53988 33100 54000
rect 37890 54432 38090 54444
rect 37890 54398 37902 54432
rect 38078 54398 38090 54432
rect 37890 54386 38090 54398
rect 37890 54344 38090 54356
rect 37890 54310 37902 54344
rect 38078 54310 38090 54344
rect 37890 54298 38090 54310
rect 37890 54122 38090 54134
rect 37890 54088 37902 54122
rect 38078 54088 38090 54122
rect 37890 54076 38090 54088
rect 37890 54034 38090 54046
rect 37890 54000 37902 54034
rect 38078 54000 38090 54034
rect 37890 53988 38090 54000
rect 42880 54432 43080 54444
rect 42880 54398 42892 54432
rect 43068 54398 43080 54432
rect 42880 54386 43080 54398
rect 42880 54344 43080 54356
rect 42880 54310 42892 54344
rect 43068 54310 43080 54344
rect 42880 54298 43080 54310
rect 42880 54122 43080 54134
rect 42880 54088 42892 54122
rect 43068 54088 43080 54122
rect 42880 54076 43080 54088
rect 42880 54034 43080 54046
rect 42880 54000 42892 54034
rect 43068 54000 43080 54034
rect 42880 53988 43080 54000
rect 47870 54432 48070 54444
rect 47870 54398 47882 54432
rect 48058 54398 48070 54432
rect 47870 54386 48070 54398
rect 47870 54344 48070 54356
rect 47870 54310 47882 54344
rect 48058 54310 48070 54344
rect 47870 54298 48070 54310
rect 47870 54122 48070 54134
rect 47870 54088 47882 54122
rect 48058 54088 48070 54122
rect 47870 54076 48070 54088
rect 47870 54034 48070 54046
rect 47870 54000 47882 54034
rect 48058 54000 48070 54034
rect 47870 53988 48070 54000
rect 52860 54432 53060 54444
rect 52860 54398 52872 54432
rect 53048 54398 53060 54432
rect 52860 54386 53060 54398
rect 52860 54344 53060 54356
rect 52860 54310 52872 54344
rect 53048 54310 53060 54344
rect 52860 54298 53060 54310
rect 52860 54122 53060 54134
rect 52860 54088 52872 54122
rect 53048 54088 53060 54122
rect 52860 54076 53060 54088
rect 52860 54034 53060 54046
rect 52860 54000 52872 54034
rect 53048 54000 53060 54034
rect 52860 53988 53060 54000
rect 57850 54432 58050 54444
rect 57850 54398 57862 54432
rect 58038 54398 58050 54432
rect 57850 54386 58050 54398
rect 57850 54344 58050 54356
rect 57850 54310 57862 54344
rect 58038 54310 58050 54344
rect 57850 54298 58050 54310
rect 57850 54122 58050 54134
rect 57850 54088 57862 54122
rect 58038 54088 58050 54122
rect 57850 54076 58050 54088
rect 57850 54034 58050 54046
rect 57850 54000 57862 54034
rect 58038 54000 58050 54034
rect 57850 53988 58050 54000
rect 62840 54432 63040 54444
rect 62840 54398 62852 54432
rect 63028 54398 63040 54432
rect 62840 54386 63040 54398
rect 62840 54344 63040 54356
rect 62840 54310 62852 54344
rect 63028 54310 63040 54344
rect 62840 54298 63040 54310
rect 62840 54122 63040 54134
rect 62840 54088 62852 54122
rect 63028 54088 63040 54122
rect 62840 54076 63040 54088
rect 62840 54034 63040 54046
rect 62840 54000 62852 54034
rect 63028 54000 63040 54034
rect 62840 53988 63040 54000
rect 67830 54432 68030 54444
rect 67830 54398 67842 54432
rect 68018 54398 68030 54432
rect 67830 54386 68030 54398
rect 67830 54344 68030 54356
rect 67830 54310 67842 54344
rect 68018 54310 68030 54344
rect 67830 54298 68030 54310
rect 67830 54122 68030 54134
rect 67830 54088 67842 54122
rect 68018 54088 68030 54122
rect 67830 54076 68030 54088
rect 67830 54034 68030 54046
rect 67830 54000 67842 54034
rect 68018 54000 68030 54034
rect 67830 53988 68030 54000
rect 72820 54432 73020 54444
rect 72820 54398 72832 54432
rect 73008 54398 73020 54432
rect 72820 54386 73020 54398
rect 72820 54344 73020 54356
rect 72820 54310 72832 54344
rect 73008 54310 73020 54344
rect 72820 54298 73020 54310
rect 72820 54122 73020 54134
rect 72820 54088 72832 54122
rect 73008 54088 73020 54122
rect 72820 54076 73020 54088
rect 72820 54034 73020 54046
rect 72820 54000 72832 54034
rect 73008 54000 73020 54034
rect 72820 53988 73020 54000
rect 77810 54432 78010 54444
rect 77810 54398 77822 54432
rect 77998 54398 78010 54432
rect 77810 54386 78010 54398
rect 77810 54344 78010 54356
rect 77810 54310 77822 54344
rect 77998 54310 78010 54344
rect 77810 54298 78010 54310
rect 77810 54122 78010 54134
rect 77810 54088 77822 54122
rect 77998 54088 78010 54122
rect 77810 54076 78010 54088
rect 77810 54034 78010 54046
rect 77810 54000 77822 54034
rect 77998 54000 78010 54034
rect 77810 53988 78010 54000
rect 2960 52722 3160 52734
rect 2960 52688 2972 52722
rect 3148 52688 3160 52722
rect 2960 52676 3160 52688
rect 2960 52634 3160 52646
rect 2960 52600 2972 52634
rect 3148 52600 3160 52634
rect 2960 52588 3160 52600
rect 2960 52412 3160 52424
rect 2960 52378 2972 52412
rect 3148 52378 3160 52412
rect 2960 52366 3160 52378
rect 2960 52324 3160 52336
rect 2960 52290 2972 52324
rect 3148 52290 3160 52324
rect 2960 52278 3160 52290
rect 7950 52722 8150 52734
rect 7950 52688 7962 52722
rect 8138 52688 8150 52722
rect 7950 52676 8150 52688
rect 7950 52634 8150 52646
rect 7950 52600 7962 52634
rect 8138 52600 8150 52634
rect 7950 52588 8150 52600
rect 7950 52412 8150 52424
rect 7950 52378 7962 52412
rect 8138 52378 8150 52412
rect 7950 52366 8150 52378
rect 7950 52324 8150 52336
rect 7950 52290 7962 52324
rect 8138 52290 8150 52324
rect 7950 52278 8150 52290
rect 12940 52722 13140 52734
rect 12940 52688 12952 52722
rect 13128 52688 13140 52722
rect 12940 52676 13140 52688
rect 12940 52634 13140 52646
rect 12940 52600 12952 52634
rect 13128 52600 13140 52634
rect 12940 52588 13140 52600
rect 12940 52412 13140 52424
rect 12940 52378 12952 52412
rect 13128 52378 13140 52412
rect 12940 52366 13140 52378
rect 12940 52324 13140 52336
rect 12940 52290 12952 52324
rect 13128 52290 13140 52324
rect 12940 52278 13140 52290
rect 17930 52722 18130 52734
rect 17930 52688 17942 52722
rect 18118 52688 18130 52722
rect 17930 52676 18130 52688
rect 17930 52634 18130 52646
rect 17930 52600 17942 52634
rect 18118 52600 18130 52634
rect 17930 52588 18130 52600
rect 17930 52412 18130 52424
rect 17930 52378 17942 52412
rect 18118 52378 18130 52412
rect 17930 52366 18130 52378
rect 17930 52324 18130 52336
rect 17930 52290 17942 52324
rect 18118 52290 18130 52324
rect 17930 52278 18130 52290
rect 22920 52722 23120 52734
rect 22920 52688 22932 52722
rect 23108 52688 23120 52722
rect 22920 52676 23120 52688
rect 22920 52634 23120 52646
rect 22920 52600 22932 52634
rect 23108 52600 23120 52634
rect 22920 52588 23120 52600
rect 22920 52412 23120 52424
rect 22920 52378 22932 52412
rect 23108 52378 23120 52412
rect 22920 52366 23120 52378
rect 22920 52324 23120 52336
rect 22920 52290 22932 52324
rect 23108 52290 23120 52324
rect 22920 52278 23120 52290
rect 27910 52722 28110 52734
rect 27910 52688 27922 52722
rect 28098 52688 28110 52722
rect 27910 52676 28110 52688
rect 27910 52634 28110 52646
rect 27910 52600 27922 52634
rect 28098 52600 28110 52634
rect 27910 52588 28110 52600
rect 27910 52412 28110 52424
rect 27910 52378 27922 52412
rect 28098 52378 28110 52412
rect 27910 52366 28110 52378
rect 27910 52324 28110 52336
rect 27910 52290 27922 52324
rect 28098 52290 28110 52324
rect 27910 52278 28110 52290
rect 32900 52722 33100 52734
rect 32900 52688 32912 52722
rect 33088 52688 33100 52722
rect 32900 52676 33100 52688
rect 32900 52634 33100 52646
rect 32900 52600 32912 52634
rect 33088 52600 33100 52634
rect 32900 52588 33100 52600
rect 32900 52412 33100 52424
rect 32900 52378 32912 52412
rect 33088 52378 33100 52412
rect 32900 52366 33100 52378
rect 32900 52324 33100 52336
rect 32900 52290 32912 52324
rect 33088 52290 33100 52324
rect 32900 52278 33100 52290
rect 37890 52722 38090 52734
rect 37890 52688 37902 52722
rect 38078 52688 38090 52722
rect 37890 52676 38090 52688
rect 37890 52634 38090 52646
rect 37890 52600 37902 52634
rect 38078 52600 38090 52634
rect 37890 52588 38090 52600
rect 37890 52412 38090 52424
rect 37890 52378 37902 52412
rect 38078 52378 38090 52412
rect 37890 52366 38090 52378
rect 37890 52324 38090 52336
rect 37890 52290 37902 52324
rect 38078 52290 38090 52324
rect 37890 52278 38090 52290
rect 42880 52722 43080 52734
rect 42880 52688 42892 52722
rect 43068 52688 43080 52722
rect 42880 52676 43080 52688
rect 42880 52634 43080 52646
rect 42880 52600 42892 52634
rect 43068 52600 43080 52634
rect 42880 52588 43080 52600
rect 42880 52412 43080 52424
rect 42880 52378 42892 52412
rect 43068 52378 43080 52412
rect 42880 52366 43080 52378
rect 42880 52324 43080 52336
rect 42880 52290 42892 52324
rect 43068 52290 43080 52324
rect 42880 52278 43080 52290
rect 47870 52722 48070 52734
rect 47870 52688 47882 52722
rect 48058 52688 48070 52722
rect 47870 52676 48070 52688
rect 47870 52634 48070 52646
rect 47870 52600 47882 52634
rect 48058 52600 48070 52634
rect 47870 52588 48070 52600
rect 47870 52412 48070 52424
rect 47870 52378 47882 52412
rect 48058 52378 48070 52412
rect 47870 52366 48070 52378
rect 47870 52324 48070 52336
rect 47870 52290 47882 52324
rect 48058 52290 48070 52324
rect 47870 52278 48070 52290
rect 52860 52722 53060 52734
rect 52860 52688 52872 52722
rect 53048 52688 53060 52722
rect 52860 52676 53060 52688
rect 52860 52634 53060 52646
rect 52860 52600 52872 52634
rect 53048 52600 53060 52634
rect 52860 52588 53060 52600
rect 52860 52412 53060 52424
rect 52860 52378 52872 52412
rect 53048 52378 53060 52412
rect 52860 52366 53060 52378
rect 52860 52324 53060 52336
rect 52860 52290 52872 52324
rect 53048 52290 53060 52324
rect 52860 52278 53060 52290
rect 57850 52722 58050 52734
rect 57850 52688 57862 52722
rect 58038 52688 58050 52722
rect 57850 52676 58050 52688
rect 57850 52634 58050 52646
rect 57850 52600 57862 52634
rect 58038 52600 58050 52634
rect 57850 52588 58050 52600
rect 57850 52412 58050 52424
rect 57850 52378 57862 52412
rect 58038 52378 58050 52412
rect 57850 52366 58050 52378
rect 57850 52324 58050 52336
rect 57850 52290 57862 52324
rect 58038 52290 58050 52324
rect 57850 52278 58050 52290
rect 62840 52722 63040 52734
rect 62840 52688 62852 52722
rect 63028 52688 63040 52722
rect 62840 52676 63040 52688
rect 62840 52634 63040 52646
rect 62840 52600 62852 52634
rect 63028 52600 63040 52634
rect 62840 52588 63040 52600
rect 62840 52412 63040 52424
rect 62840 52378 62852 52412
rect 63028 52378 63040 52412
rect 62840 52366 63040 52378
rect 62840 52324 63040 52336
rect 62840 52290 62852 52324
rect 63028 52290 63040 52324
rect 62840 52278 63040 52290
rect 67830 52722 68030 52734
rect 67830 52688 67842 52722
rect 68018 52688 68030 52722
rect 67830 52676 68030 52688
rect 67830 52634 68030 52646
rect 67830 52600 67842 52634
rect 68018 52600 68030 52634
rect 67830 52588 68030 52600
rect 67830 52412 68030 52424
rect 67830 52378 67842 52412
rect 68018 52378 68030 52412
rect 67830 52366 68030 52378
rect 67830 52324 68030 52336
rect 67830 52290 67842 52324
rect 68018 52290 68030 52324
rect 67830 52278 68030 52290
rect 72820 52722 73020 52734
rect 72820 52688 72832 52722
rect 73008 52688 73020 52722
rect 72820 52676 73020 52688
rect 72820 52634 73020 52646
rect 72820 52600 72832 52634
rect 73008 52600 73020 52634
rect 72820 52588 73020 52600
rect 72820 52412 73020 52424
rect 72820 52378 72832 52412
rect 73008 52378 73020 52412
rect 72820 52366 73020 52378
rect 72820 52324 73020 52336
rect 72820 52290 72832 52324
rect 73008 52290 73020 52324
rect 72820 52278 73020 52290
rect 77810 52722 78010 52734
rect 77810 52688 77822 52722
rect 77998 52688 78010 52722
rect 77810 52676 78010 52688
rect 77810 52634 78010 52646
rect 77810 52600 77822 52634
rect 77998 52600 78010 52634
rect 77810 52588 78010 52600
rect 77810 52412 78010 52424
rect 77810 52378 77822 52412
rect 77998 52378 78010 52412
rect 77810 52366 78010 52378
rect 77810 52324 78010 52336
rect 77810 52290 77822 52324
rect 77998 52290 78010 52324
rect 77810 52278 78010 52290
rect 2960 51012 3160 51024
rect 2960 50978 2972 51012
rect 3148 50978 3160 51012
rect 2960 50966 3160 50978
rect 2960 50924 3160 50936
rect 2960 50890 2972 50924
rect 3148 50890 3160 50924
rect 2960 50878 3160 50890
rect 2960 50702 3160 50714
rect 2960 50668 2972 50702
rect 3148 50668 3160 50702
rect 2960 50656 3160 50668
rect 2960 50614 3160 50626
rect 2960 50580 2972 50614
rect 3148 50580 3160 50614
rect 2960 50568 3160 50580
rect 7950 51012 8150 51024
rect 7950 50978 7962 51012
rect 8138 50978 8150 51012
rect 7950 50966 8150 50978
rect 7950 50924 8150 50936
rect 7950 50890 7962 50924
rect 8138 50890 8150 50924
rect 7950 50878 8150 50890
rect 7950 50702 8150 50714
rect 7950 50668 7962 50702
rect 8138 50668 8150 50702
rect 7950 50656 8150 50668
rect 7950 50614 8150 50626
rect 7950 50580 7962 50614
rect 8138 50580 8150 50614
rect 7950 50568 8150 50580
rect 12940 51012 13140 51024
rect 12940 50978 12952 51012
rect 13128 50978 13140 51012
rect 12940 50966 13140 50978
rect 12940 50924 13140 50936
rect 12940 50890 12952 50924
rect 13128 50890 13140 50924
rect 12940 50878 13140 50890
rect 12940 50702 13140 50714
rect 12940 50668 12952 50702
rect 13128 50668 13140 50702
rect 12940 50656 13140 50668
rect 12940 50614 13140 50626
rect 12940 50580 12952 50614
rect 13128 50580 13140 50614
rect 12940 50568 13140 50580
rect 17930 51012 18130 51024
rect 17930 50978 17942 51012
rect 18118 50978 18130 51012
rect 17930 50966 18130 50978
rect 17930 50924 18130 50936
rect 17930 50890 17942 50924
rect 18118 50890 18130 50924
rect 17930 50878 18130 50890
rect 17930 50702 18130 50714
rect 17930 50668 17942 50702
rect 18118 50668 18130 50702
rect 17930 50656 18130 50668
rect 17930 50614 18130 50626
rect 17930 50580 17942 50614
rect 18118 50580 18130 50614
rect 17930 50568 18130 50580
rect 22920 51012 23120 51024
rect 22920 50978 22932 51012
rect 23108 50978 23120 51012
rect 22920 50966 23120 50978
rect 22920 50924 23120 50936
rect 22920 50890 22932 50924
rect 23108 50890 23120 50924
rect 22920 50878 23120 50890
rect 22920 50702 23120 50714
rect 22920 50668 22932 50702
rect 23108 50668 23120 50702
rect 22920 50656 23120 50668
rect 22920 50614 23120 50626
rect 22920 50580 22932 50614
rect 23108 50580 23120 50614
rect 22920 50568 23120 50580
rect 27910 51012 28110 51024
rect 27910 50978 27922 51012
rect 28098 50978 28110 51012
rect 27910 50966 28110 50978
rect 27910 50924 28110 50936
rect 27910 50890 27922 50924
rect 28098 50890 28110 50924
rect 27910 50878 28110 50890
rect 27910 50702 28110 50714
rect 27910 50668 27922 50702
rect 28098 50668 28110 50702
rect 27910 50656 28110 50668
rect 27910 50614 28110 50626
rect 27910 50580 27922 50614
rect 28098 50580 28110 50614
rect 27910 50568 28110 50580
rect 32900 51012 33100 51024
rect 32900 50978 32912 51012
rect 33088 50978 33100 51012
rect 32900 50966 33100 50978
rect 32900 50924 33100 50936
rect 32900 50890 32912 50924
rect 33088 50890 33100 50924
rect 32900 50878 33100 50890
rect 32900 50702 33100 50714
rect 32900 50668 32912 50702
rect 33088 50668 33100 50702
rect 32900 50656 33100 50668
rect 32900 50614 33100 50626
rect 32900 50580 32912 50614
rect 33088 50580 33100 50614
rect 32900 50568 33100 50580
rect 37890 51012 38090 51024
rect 37890 50978 37902 51012
rect 38078 50978 38090 51012
rect 37890 50966 38090 50978
rect 37890 50924 38090 50936
rect 37890 50890 37902 50924
rect 38078 50890 38090 50924
rect 37890 50878 38090 50890
rect 37890 50702 38090 50714
rect 37890 50668 37902 50702
rect 38078 50668 38090 50702
rect 37890 50656 38090 50668
rect 37890 50614 38090 50626
rect 37890 50580 37902 50614
rect 38078 50580 38090 50614
rect 37890 50568 38090 50580
rect 42880 51012 43080 51024
rect 42880 50978 42892 51012
rect 43068 50978 43080 51012
rect 42880 50966 43080 50978
rect 42880 50924 43080 50936
rect 42880 50890 42892 50924
rect 43068 50890 43080 50924
rect 42880 50878 43080 50890
rect 42880 50702 43080 50714
rect 42880 50668 42892 50702
rect 43068 50668 43080 50702
rect 42880 50656 43080 50668
rect 42880 50614 43080 50626
rect 42880 50580 42892 50614
rect 43068 50580 43080 50614
rect 42880 50568 43080 50580
rect 47870 51012 48070 51024
rect 47870 50978 47882 51012
rect 48058 50978 48070 51012
rect 47870 50966 48070 50978
rect 47870 50924 48070 50936
rect 47870 50890 47882 50924
rect 48058 50890 48070 50924
rect 47870 50878 48070 50890
rect 47870 50702 48070 50714
rect 47870 50668 47882 50702
rect 48058 50668 48070 50702
rect 47870 50656 48070 50668
rect 47870 50614 48070 50626
rect 47870 50580 47882 50614
rect 48058 50580 48070 50614
rect 47870 50568 48070 50580
rect 52860 51012 53060 51024
rect 52860 50978 52872 51012
rect 53048 50978 53060 51012
rect 52860 50966 53060 50978
rect 52860 50924 53060 50936
rect 52860 50890 52872 50924
rect 53048 50890 53060 50924
rect 52860 50878 53060 50890
rect 52860 50702 53060 50714
rect 52860 50668 52872 50702
rect 53048 50668 53060 50702
rect 52860 50656 53060 50668
rect 52860 50614 53060 50626
rect 52860 50580 52872 50614
rect 53048 50580 53060 50614
rect 52860 50568 53060 50580
rect 57850 51012 58050 51024
rect 57850 50978 57862 51012
rect 58038 50978 58050 51012
rect 57850 50966 58050 50978
rect 57850 50924 58050 50936
rect 57850 50890 57862 50924
rect 58038 50890 58050 50924
rect 57850 50878 58050 50890
rect 57850 50702 58050 50714
rect 57850 50668 57862 50702
rect 58038 50668 58050 50702
rect 57850 50656 58050 50668
rect 57850 50614 58050 50626
rect 57850 50580 57862 50614
rect 58038 50580 58050 50614
rect 57850 50568 58050 50580
rect 62840 51012 63040 51024
rect 62840 50978 62852 51012
rect 63028 50978 63040 51012
rect 62840 50966 63040 50978
rect 62840 50924 63040 50936
rect 62840 50890 62852 50924
rect 63028 50890 63040 50924
rect 62840 50878 63040 50890
rect 62840 50702 63040 50714
rect 62840 50668 62852 50702
rect 63028 50668 63040 50702
rect 62840 50656 63040 50668
rect 62840 50614 63040 50626
rect 62840 50580 62852 50614
rect 63028 50580 63040 50614
rect 62840 50568 63040 50580
rect 67830 51012 68030 51024
rect 67830 50978 67842 51012
rect 68018 50978 68030 51012
rect 67830 50966 68030 50978
rect 67830 50924 68030 50936
rect 67830 50890 67842 50924
rect 68018 50890 68030 50924
rect 67830 50878 68030 50890
rect 67830 50702 68030 50714
rect 67830 50668 67842 50702
rect 68018 50668 68030 50702
rect 67830 50656 68030 50668
rect 67830 50614 68030 50626
rect 67830 50580 67842 50614
rect 68018 50580 68030 50614
rect 67830 50568 68030 50580
rect 72820 51012 73020 51024
rect 72820 50978 72832 51012
rect 73008 50978 73020 51012
rect 72820 50966 73020 50978
rect 72820 50924 73020 50936
rect 72820 50890 72832 50924
rect 73008 50890 73020 50924
rect 72820 50878 73020 50890
rect 72820 50702 73020 50714
rect 72820 50668 72832 50702
rect 73008 50668 73020 50702
rect 72820 50656 73020 50668
rect 72820 50614 73020 50626
rect 72820 50580 72832 50614
rect 73008 50580 73020 50614
rect 72820 50568 73020 50580
rect 77810 51012 78010 51024
rect 77810 50978 77822 51012
rect 77998 50978 78010 51012
rect 77810 50966 78010 50978
rect 77810 50924 78010 50936
rect 77810 50890 77822 50924
rect 77998 50890 78010 50924
rect 77810 50878 78010 50890
rect 77810 50702 78010 50714
rect 77810 50668 77822 50702
rect 77998 50668 78010 50702
rect 77810 50656 78010 50668
rect 77810 50614 78010 50626
rect 77810 50580 77822 50614
rect 77998 50580 78010 50614
rect 77810 50568 78010 50580
rect 2960 49302 3160 49314
rect 2960 49268 2972 49302
rect 3148 49268 3160 49302
rect 2960 49256 3160 49268
rect 2960 49214 3160 49226
rect 2960 49180 2972 49214
rect 3148 49180 3160 49214
rect 2960 49168 3160 49180
rect 2960 48992 3160 49004
rect 2960 48958 2972 48992
rect 3148 48958 3160 48992
rect 2960 48946 3160 48958
rect 2960 48904 3160 48916
rect 2960 48870 2972 48904
rect 3148 48870 3160 48904
rect 2960 48858 3160 48870
rect 7950 49302 8150 49314
rect 7950 49268 7962 49302
rect 8138 49268 8150 49302
rect 7950 49256 8150 49268
rect 7950 49214 8150 49226
rect 7950 49180 7962 49214
rect 8138 49180 8150 49214
rect 7950 49168 8150 49180
rect 7950 48992 8150 49004
rect 7950 48958 7962 48992
rect 8138 48958 8150 48992
rect 7950 48946 8150 48958
rect 7950 48904 8150 48916
rect 7950 48870 7962 48904
rect 8138 48870 8150 48904
rect 7950 48858 8150 48870
rect 12940 49302 13140 49314
rect 12940 49268 12952 49302
rect 13128 49268 13140 49302
rect 12940 49256 13140 49268
rect 12940 49214 13140 49226
rect 12940 49180 12952 49214
rect 13128 49180 13140 49214
rect 12940 49168 13140 49180
rect 12940 48992 13140 49004
rect 12940 48958 12952 48992
rect 13128 48958 13140 48992
rect 12940 48946 13140 48958
rect 12940 48904 13140 48916
rect 12940 48870 12952 48904
rect 13128 48870 13140 48904
rect 12940 48858 13140 48870
rect 17930 49302 18130 49314
rect 17930 49268 17942 49302
rect 18118 49268 18130 49302
rect 17930 49256 18130 49268
rect 17930 49214 18130 49226
rect 17930 49180 17942 49214
rect 18118 49180 18130 49214
rect 17930 49168 18130 49180
rect 17930 48992 18130 49004
rect 17930 48958 17942 48992
rect 18118 48958 18130 48992
rect 17930 48946 18130 48958
rect 17930 48904 18130 48916
rect 17930 48870 17942 48904
rect 18118 48870 18130 48904
rect 17930 48858 18130 48870
rect 22920 49302 23120 49314
rect 22920 49268 22932 49302
rect 23108 49268 23120 49302
rect 22920 49256 23120 49268
rect 22920 49214 23120 49226
rect 22920 49180 22932 49214
rect 23108 49180 23120 49214
rect 22920 49168 23120 49180
rect 22920 48992 23120 49004
rect 22920 48958 22932 48992
rect 23108 48958 23120 48992
rect 22920 48946 23120 48958
rect 22920 48904 23120 48916
rect 22920 48870 22932 48904
rect 23108 48870 23120 48904
rect 22920 48858 23120 48870
rect 27910 49302 28110 49314
rect 27910 49268 27922 49302
rect 28098 49268 28110 49302
rect 27910 49256 28110 49268
rect 27910 49214 28110 49226
rect 27910 49180 27922 49214
rect 28098 49180 28110 49214
rect 27910 49168 28110 49180
rect 27910 48992 28110 49004
rect 27910 48958 27922 48992
rect 28098 48958 28110 48992
rect 27910 48946 28110 48958
rect 27910 48904 28110 48916
rect 27910 48870 27922 48904
rect 28098 48870 28110 48904
rect 27910 48858 28110 48870
rect 32900 49302 33100 49314
rect 32900 49268 32912 49302
rect 33088 49268 33100 49302
rect 32900 49256 33100 49268
rect 32900 49214 33100 49226
rect 32900 49180 32912 49214
rect 33088 49180 33100 49214
rect 32900 49168 33100 49180
rect 32900 48992 33100 49004
rect 32900 48958 32912 48992
rect 33088 48958 33100 48992
rect 32900 48946 33100 48958
rect 32900 48904 33100 48916
rect 32900 48870 32912 48904
rect 33088 48870 33100 48904
rect 32900 48858 33100 48870
rect 37890 49302 38090 49314
rect 37890 49268 37902 49302
rect 38078 49268 38090 49302
rect 37890 49256 38090 49268
rect 37890 49214 38090 49226
rect 37890 49180 37902 49214
rect 38078 49180 38090 49214
rect 37890 49168 38090 49180
rect 37890 48992 38090 49004
rect 37890 48958 37902 48992
rect 38078 48958 38090 48992
rect 37890 48946 38090 48958
rect 37890 48904 38090 48916
rect 37890 48870 37902 48904
rect 38078 48870 38090 48904
rect 37890 48858 38090 48870
rect 42880 49302 43080 49314
rect 42880 49268 42892 49302
rect 43068 49268 43080 49302
rect 42880 49256 43080 49268
rect 42880 49214 43080 49226
rect 42880 49180 42892 49214
rect 43068 49180 43080 49214
rect 42880 49168 43080 49180
rect 42880 48992 43080 49004
rect 42880 48958 42892 48992
rect 43068 48958 43080 48992
rect 42880 48946 43080 48958
rect 42880 48904 43080 48916
rect 42880 48870 42892 48904
rect 43068 48870 43080 48904
rect 42880 48858 43080 48870
rect 47870 49302 48070 49314
rect 47870 49268 47882 49302
rect 48058 49268 48070 49302
rect 47870 49256 48070 49268
rect 47870 49214 48070 49226
rect 47870 49180 47882 49214
rect 48058 49180 48070 49214
rect 47870 49168 48070 49180
rect 47870 48992 48070 49004
rect 47870 48958 47882 48992
rect 48058 48958 48070 48992
rect 47870 48946 48070 48958
rect 47870 48904 48070 48916
rect 47870 48870 47882 48904
rect 48058 48870 48070 48904
rect 47870 48858 48070 48870
rect 52860 49302 53060 49314
rect 52860 49268 52872 49302
rect 53048 49268 53060 49302
rect 52860 49256 53060 49268
rect 52860 49214 53060 49226
rect 52860 49180 52872 49214
rect 53048 49180 53060 49214
rect 52860 49168 53060 49180
rect 52860 48992 53060 49004
rect 52860 48958 52872 48992
rect 53048 48958 53060 48992
rect 52860 48946 53060 48958
rect 52860 48904 53060 48916
rect 52860 48870 52872 48904
rect 53048 48870 53060 48904
rect 52860 48858 53060 48870
rect 57850 49302 58050 49314
rect 57850 49268 57862 49302
rect 58038 49268 58050 49302
rect 57850 49256 58050 49268
rect 57850 49214 58050 49226
rect 57850 49180 57862 49214
rect 58038 49180 58050 49214
rect 57850 49168 58050 49180
rect 57850 48992 58050 49004
rect 57850 48958 57862 48992
rect 58038 48958 58050 48992
rect 57850 48946 58050 48958
rect 57850 48904 58050 48916
rect 57850 48870 57862 48904
rect 58038 48870 58050 48904
rect 57850 48858 58050 48870
rect 62840 49302 63040 49314
rect 62840 49268 62852 49302
rect 63028 49268 63040 49302
rect 62840 49256 63040 49268
rect 62840 49214 63040 49226
rect 62840 49180 62852 49214
rect 63028 49180 63040 49214
rect 62840 49168 63040 49180
rect 62840 48992 63040 49004
rect 62840 48958 62852 48992
rect 63028 48958 63040 48992
rect 62840 48946 63040 48958
rect 62840 48904 63040 48916
rect 62840 48870 62852 48904
rect 63028 48870 63040 48904
rect 62840 48858 63040 48870
rect 67830 49302 68030 49314
rect 67830 49268 67842 49302
rect 68018 49268 68030 49302
rect 67830 49256 68030 49268
rect 67830 49214 68030 49226
rect 67830 49180 67842 49214
rect 68018 49180 68030 49214
rect 67830 49168 68030 49180
rect 67830 48992 68030 49004
rect 67830 48958 67842 48992
rect 68018 48958 68030 48992
rect 67830 48946 68030 48958
rect 67830 48904 68030 48916
rect 67830 48870 67842 48904
rect 68018 48870 68030 48904
rect 67830 48858 68030 48870
rect 72820 49302 73020 49314
rect 72820 49268 72832 49302
rect 73008 49268 73020 49302
rect 72820 49256 73020 49268
rect 72820 49214 73020 49226
rect 72820 49180 72832 49214
rect 73008 49180 73020 49214
rect 72820 49168 73020 49180
rect 72820 48992 73020 49004
rect 72820 48958 72832 48992
rect 73008 48958 73020 48992
rect 72820 48946 73020 48958
rect 72820 48904 73020 48916
rect 72820 48870 72832 48904
rect 73008 48870 73020 48904
rect 72820 48858 73020 48870
rect 77810 49302 78010 49314
rect 77810 49268 77822 49302
rect 77998 49268 78010 49302
rect 77810 49256 78010 49268
rect 77810 49214 78010 49226
rect 77810 49180 77822 49214
rect 77998 49180 78010 49214
rect 77810 49168 78010 49180
rect 77810 48992 78010 49004
rect 77810 48958 77822 48992
rect 77998 48958 78010 48992
rect 77810 48946 78010 48958
rect 77810 48904 78010 48916
rect 77810 48870 77822 48904
rect 77998 48870 78010 48904
rect 77810 48858 78010 48870
rect 2960 47592 3160 47604
rect 2960 47558 2972 47592
rect 3148 47558 3160 47592
rect 2960 47546 3160 47558
rect 2960 47504 3160 47516
rect 2960 47470 2972 47504
rect 3148 47470 3160 47504
rect 2960 47458 3160 47470
rect 2960 47282 3160 47294
rect 2960 47248 2972 47282
rect 3148 47248 3160 47282
rect 2960 47236 3160 47248
rect 2960 47194 3160 47206
rect 2960 47160 2972 47194
rect 3148 47160 3160 47194
rect 2960 47148 3160 47160
rect 7950 47592 8150 47604
rect 7950 47558 7962 47592
rect 8138 47558 8150 47592
rect 7950 47546 8150 47558
rect 7950 47504 8150 47516
rect 7950 47470 7962 47504
rect 8138 47470 8150 47504
rect 7950 47458 8150 47470
rect 7950 47282 8150 47294
rect 7950 47248 7962 47282
rect 8138 47248 8150 47282
rect 7950 47236 8150 47248
rect 7950 47194 8150 47206
rect 7950 47160 7962 47194
rect 8138 47160 8150 47194
rect 7950 47148 8150 47160
rect 12940 47592 13140 47604
rect 12940 47558 12952 47592
rect 13128 47558 13140 47592
rect 12940 47546 13140 47558
rect 12940 47504 13140 47516
rect 12940 47470 12952 47504
rect 13128 47470 13140 47504
rect 12940 47458 13140 47470
rect 12940 47282 13140 47294
rect 12940 47248 12952 47282
rect 13128 47248 13140 47282
rect 12940 47236 13140 47248
rect 12940 47194 13140 47206
rect 12940 47160 12952 47194
rect 13128 47160 13140 47194
rect 12940 47148 13140 47160
rect 17930 47592 18130 47604
rect 17930 47558 17942 47592
rect 18118 47558 18130 47592
rect 17930 47546 18130 47558
rect 17930 47504 18130 47516
rect 17930 47470 17942 47504
rect 18118 47470 18130 47504
rect 17930 47458 18130 47470
rect 17930 47282 18130 47294
rect 17930 47248 17942 47282
rect 18118 47248 18130 47282
rect 17930 47236 18130 47248
rect 17930 47194 18130 47206
rect 17930 47160 17942 47194
rect 18118 47160 18130 47194
rect 17930 47148 18130 47160
rect 22920 47592 23120 47604
rect 22920 47558 22932 47592
rect 23108 47558 23120 47592
rect 22920 47546 23120 47558
rect 22920 47504 23120 47516
rect 22920 47470 22932 47504
rect 23108 47470 23120 47504
rect 22920 47458 23120 47470
rect 22920 47282 23120 47294
rect 22920 47248 22932 47282
rect 23108 47248 23120 47282
rect 22920 47236 23120 47248
rect 22920 47194 23120 47206
rect 22920 47160 22932 47194
rect 23108 47160 23120 47194
rect 22920 47148 23120 47160
rect 27910 47592 28110 47604
rect 27910 47558 27922 47592
rect 28098 47558 28110 47592
rect 27910 47546 28110 47558
rect 27910 47504 28110 47516
rect 27910 47470 27922 47504
rect 28098 47470 28110 47504
rect 27910 47458 28110 47470
rect 27910 47282 28110 47294
rect 27910 47248 27922 47282
rect 28098 47248 28110 47282
rect 27910 47236 28110 47248
rect 27910 47194 28110 47206
rect 27910 47160 27922 47194
rect 28098 47160 28110 47194
rect 27910 47148 28110 47160
rect 32900 47592 33100 47604
rect 32900 47558 32912 47592
rect 33088 47558 33100 47592
rect 32900 47546 33100 47558
rect 32900 47504 33100 47516
rect 32900 47470 32912 47504
rect 33088 47470 33100 47504
rect 32900 47458 33100 47470
rect 32900 47282 33100 47294
rect 32900 47248 32912 47282
rect 33088 47248 33100 47282
rect 32900 47236 33100 47248
rect 32900 47194 33100 47206
rect 32900 47160 32912 47194
rect 33088 47160 33100 47194
rect 32900 47148 33100 47160
rect 37890 47592 38090 47604
rect 37890 47558 37902 47592
rect 38078 47558 38090 47592
rect 37890 47546 38090 47558
rect 37890 47504 38090 47516
rect 37890 47470 37902 47504
rect 38078 47470 38090 47504
rect 37890 47458 38090 47470
rect 37890 47282 38090 47294
rect 37890 47248 37902 47282
rect 38078 47248 38090 47282
rect 37890 47236 38090 47248
rect 37890 47194 38090 47206
rect 37890 47160 37902 47194
rect 38078 47160 38090 47194
rect 37890 47148 38090 47160
rect 42880 47592 43080 47604
rect 42880 47558 42892 47592
rect 43068 47558 43080 47592
rect 42880 47546 43080 47558
rect 42880 47504 43080 47516
rect 42880 47470 42892 47504
rect 43068 47470 43080 47504
rect 42880 47458 43080 47470
rect 42880 47282 43080 47294
rect 42880 47248 42892 47282
rect 43068 47248 43080 47282
rect 42880 47236 43080 47248
rect 42880 47194 43080 47206
rect 42880 47160 42892 47194
rect 43068 47160 43080 47194
rect 42880 47148 43080 47160
rect 47870 47592 48070 47604
rect 47870 47558 47882 47592
rect 48058 47558 48070 47592
rect 47870 47546 48070 47558
rect 47870 47504 48070 47516
rect 47870 47470 47882 47504
rect 48058 47470 48070 47504
rect 47870 47458 48070 47470
rect 47870 47282 48070 47294
rect 47870 47248 47882 47282
rect 48058 47248 48070 47282
rect 47870 47236 48070 47248
rect 47870 47194 48070 47206
rect 47870 47160 47882 47194
rect 48058 47160 48070 47194
rect 47870 47148 48070 47160
rect 52860 47592 53060 47604
rect 52860 47558 52872 47592
rect 53048 47558 53060 47592
rect 52860 47546 53060 47558
rect 52860 47504 53060 47516
rect 52860 47470 52872 47504
rect 53048 47470 53060 47504
rect 52860 47458 53060 47470
rect 52860 47282 53060 47294
rect 52860 47248 52872 47282
rect 53048 47248 53060 47282
rect 52860 47236 53060 47248
rect 52860 47194 53060 47206
rect 52860 47160 52872 47194
rect 53048 47160 53060 47194
rect 52860 47148 53060 47160
rect 57850 47592 58050 47604
rect 57850 47558 57862 47592
rect 58038 47558 58050 47592
rect 57850 47546 58050 47558
rect 57850 47504 58050 47516
rect 57850 47470 57862 47504
rect 58038 47470 58050 47504
rect 57850 47458 58050 47470
rect 57850 47282 58050 47294
rect 57850 47248 57862 47282
rect 58038 47248 58050 47282
rect 57850 47236 58050 47248
rect 57850 47194 58050 47206
rect 57850 47160 57862 47194
rect 58038 47160 58050 47194
rect 57850 47148 58050 47160
rect 62840 47592 63040 47604
rect 62840 47558 62852 47592
rect 63028 47558 63040 47592
rect 62840 47546 63040 47558
rect 62840 47504 63040 47516
rect 62840 47470 62852 47504
rect 63028 47470 63040 47504
rect 62840 47458 63040 47470
rect 62840 47282 63040 47294
rect 62840 47248 62852 47282
rect 63028 47248 63040 47282
rect 62840 47236 63040 47248
rect 62840 47194 63040 47206
rect 62840 47160 62852 47194
rect 63028 47160 63040 47194
rect 62840 47148 63040 47160
rect 67830 47592 68030 47604
rect 67830 47558 67842 47592
rect 68018 47558 68030 47592
rect 67830 47546 68030 47558
rect 67830 47504 68030 47516
rect 67830 47470 67842 47504
rect 68018 47470 68030 47504
rect 67830 47458 68030 47470
rect 67830 47282 68030 47294
rect 67830 47248 67842 47282
rect 68018 47248 68030 47282
rect 67830 47236 68030 47248
rect 67830 47194 68030 47206
rect 67830 47160 67842 47194
rect 68018 47160 68030 47194
rect 67830 47148 68030 47160
rect 72820 47592 73020 47604
rect 72820 47558 72832 47592
rect 73008 47558 73020 47592
rect 72820 47546 73020 47558
rect 72820 47504 73020 47516
rect 72820 47470 72832 47504
rect 73008 47470 73020 47504
rect 72820 47458 73020 47470
rect 72820 47282 73020 47294
rect 72820 47248 72832 47282
rect 73008 47248 73020 47282
rect 72820 47236 73020 47248
rect 72820 47194 73020 47206
rect 72820 47160 72832 47194
rect 73008 47160 73020 47194
rect 72820 47148 73020 47160
rect 77810 47592 78010 47604
rect 77810 47558 77822 47592
rect 77998 47558 78010 47592
rect 77810 47546 78010 47558
rect 77810 47504 78010 47516
rect 77810 47470 77822 47504
rect 77998 47470 78010 47504
rect 77810 47458 78010 47470
rect 77810 47282 78010 47294
rect 77810 47248 77822 47282
rect 77998 47248 78010 47282
rect 77810 47236 78010 47248
rect 77810 47194 78010 47206
rect 77810 47160 77822 47194
rect 77998 47160 78010 47194
rect 77810 47148 78010 47160
rect 2960 45882 3160 45894
rect 2960 45848 2972 45882
rect 3148 45848 3160 45882
rect 2960 45836 3160 45848
rect 2960 45794 3160 45806
rect 2960 45760 2972 45794
rect 3148 45760 3160 45794
rect 2960 45748 3160 45760
rect 2960 45572 3160 45584
rect 2960 45538 2972 45572
rect 3148 45538 3160 45572
rect 2960 45526 3160 45538
rect 2960 45484 3160 45496
rect 2960 45450 2972 45484
rect 3148 45450 3160 45484
rect 2960 45438 3160 45450
rect 7950 45882 8150 45894
rect 7950 45848 7962 45882
rect 8138 45848 8150 45882
rect 7950 45836 8150 45848
rect 7950 45794 8150 45806
rect 7950 45760 7962 45794
rect 8138 45760 8150 45794
rect 7950 45748 8150 45760
rect 7950 45572 8150 45584
rect 7950 45538 7962 45572
rect 8138 45538 8150 45572
rect 7950 45526 8150 45538
rect 7950 45484 8150 45496
rect 7950 45450 7962 45484
rect 8138 45450 8150 45484
rect 7950 45438 8150 45450
rect 12940 45882 13140 45894
rect 12940 45848 12952 45882
rect 13128 45848 13140 45882
rect 12940 45836 13140 45848
rect 12940 45794 13140 45806
rect 12940 45760 12952 45794
rect 13128 45760 13140 45794
rect 12940 45748 13140 45760
rect 12940 45572 13140 45584
rect 12940 45538 12952 45572
rect 13128 45538 13140 45572
rect 12940 45526 13140 45538
rect 12940 45484 13140 45496
rect 12940 45450 12952 45484
rect 13128 45450 13140 45484
rect 12940 45438 13140 45450
rect 17930 45882 18130 45894
rect 17930 45848 17942 45882
rect 18118 45848 18130 45882
rect 17930 45836 18130 45848
rect 17930 45794 18130 45806
rect 17930 45760 17942 45794
rect 18118 45760 18130 45794
rect 17930 45748 18130 45760
rect 17930 45572 18130 45584
rect 17930 45538 17942 45572
rect 18118 45538 18130 45572
rect 17930 45526 18130 45538
rect 17930 45484 18130 45496
rect 17930 45450 17942 45484
rect 18118 45450 18130 45484
rect 17930 45438 18130 45450
rect 22920 45882 23120 45894
rect 22920 45848 22932 45882
rect 23108 45848 23120 45882
rect 22920 45836 23120 45848
rect 22920 45794 23120 45806
rect 22920 45760 22932 45794
rect 23108 45760 23120 45794
rect 22920 45748 23120 45760
rect 22920 45572 23120 45584
rect 22920 45538 22932 45572
rect 23108 45538 23120 45572
rect 22920 45526 23120 45538
rect 22920 45484 23120 45496
rect 22920 45450 22932 45484
rect 23108 45450 23120 45484
rect 22920 45438 23120 45450
rect 27910 45882 28110 45894
rect 27910 45848 27922 45882
rect 28098 45848 28110 45882
rect 27910 45836 28110 45848
rect 27910 45794 28110 45806
rect 27910 45760 27922 45794
rect 28098 45760 28110 45794
rect 27910 45748 28110 45760
rect 27910 45572 28110 45584
rect 27910 45538 27922 45572
rect 28098 45538 28110 45572
rect 27910 45526 28110 45538
rect 27910 45484 28110 45496
rect 27910 45450 27922 45484
rect 28098 45450 28110 45484
rect 27910 45438 28110 45450
rect 32900 45882 33100 45894
rect 32900 45848 32912 45882
rect 33088 45848 33100 45882
rect 32900 45836 33100 45848
rect 32900 45794 33100 45806
rect 32900 45760 32912 45794
rect 33088 45760 33100 45794
rect 32900 45748 33100 45760
rect 32900 45572 33100 45584
rect 32900 45538 32912 45572
rect 33088 45538 33100 45572
rect 32900 45526 33100 45538
rect 32900 45484 33100 45496
rect 32900 45450 32912 45484
rect 33088 45450 33100 45484
rect 32900 45438 33100 45450
rect 37890 45882 38090 45894
rect 37890 45848 37902 45882
rect 38078 45848 38090 45882
rect 37890 45836 38090 45848
rect 37890 45794 38090 45806
rect 37890 45760 37902 45794
rect 38078 45760 38090 45794
rect 37890 45748 38090 45760
rect 37890 45572 38090 45584
rect 37890 45538 37902 45572
rect 38078 45538 38090 45572
rect 37890 45526 38090 45538
rect 37890 45484 38090 45496
rect 37890 45450 37902 45484
rect 38078 45450 38090 45484
rect 37890 45438 38090 45450
rect 42880 45882 43080 45894
rect 42880 45848 42892 45882
rect 43068 45848 43080 45882
rect 42880 45836 43080 45848
rect 42880 45794 43080 45806
rect 42880 45760 42892 45794
rect 43068 45760 43080 45794
rect 42880 45748 43080 45760
rect 42880 45572 43080 45584
rect 42880 45538 42892 45572
rect 43068 45538 43080 45572
rect 42880 45526 43080 45538
rect 42880 45484 43080 45496
rect 42880 45450 42892 45484
rect 43068 45450 43080 45484
rect 42880 45438 43080 45450
rect 47870 45882 48070 45894
rect 47870 45848 47882 45882
rect 48058 45848 48070 45882
rect 47870 45836 48070 45848
rect 47870 45794 48070 45806
rect 47870 45760 47882 45794
rect 48058 45760 48070 45794
rect 47870 45748 48070 45760
rect 47870 45572 48070 45584
rect 47870 45538 47882 45572
rect 48058 45538 48070 45572
rect 47870 45526 48070 45538
rect 47870 45484 48070 45496
rect 47870 45450 47882 45484
rect 48058 45450 48070 45484
rect 47870 45438 48070 45450
rect 52860 45882 53060 45894
rect 52860 45848 52872 45882
rect 53048 45848 53060 45882
rect 52860 45836 53060 45848
rect 52860 45794 53060 45806
rect 52860 45760 52872 45794
rect 53048 45760 53060 45794
rect 52860 45748 53060 45760
rect 52860 45572 53060 45584
rect 52860 45538 52872 45572
rect 53048 45538 53060 45572
rect 52860 45526 53060 45538
rect 52860 45484 53060 45496
rect 52860 45450 52872 45484
rect 53048 45450 53060 45484
rect 52860 45438 53060 45450
rect 57850 45882 58050 45894
rect 57850 45848 57862 45882
rect 58038 45848 58050 45882
rect 57850 45836 58050 45848
rect 57850 45794 58050 45806
rect 57850 45760 57862 45794
rect 58038 45760 58050 45794
rect 57850 45748 58050 45760
rect 57850 45572 58050 45584
rect 57850 45538 57862 45572
rect 58038 45538 58050 45572
rect 57850 45526 58050 45538
rect 57850 45484 58050 45496
rect 57850 45450 57862 45484
rect 58038 45450 58050 45484
rect 57850 45438 58050 45450
rect 62840 45882 63040 45894
rect 62840 45848 62852 45882
rect 63028 45848 63040 45882
rect 62840 45836 63040 45848
rect 62840 45794 63040 45806
rect 62840 45760 62852 45794
rect 63028 45760 63040 45794
rect 62840 45748 63040 45760
rect 62840 45572 63040 45584
rect 62840 45538 62852 45572
rect 63028 45538 63040 45572
rect 62840 45526 63040 45538
rect 62840 45484 63040 45496
rect 62840 45450 62852 45484
rect 63028 45450 63040 45484
rect 62840 45438 63040 45450
rect 67830 45882 68030 45894
rect 67830 45848 67842 45882
rect 68018 45848 68030 45882
rect 67830 45836 68030 45848
rect 67830 45794 68030 45806
rect 67830 45760 67842 45794
rect 68018 45760 68030 45794
rect 67830 45748 68030 45760
rect 67830 45572 68030 45584
rect 67830 45538 67842 45572
rect 68018 45538 68030 45572
rect 67830 45526 68030 45538
rect 67830 45484 68030 45496
rect 67830 45450 67842 45484
rect 68018 45450 68030 45484
rect 67830 45438 68030 45450
rect 72820 45882 73020 45894
rect 72820 45848 72832 45882
rect 73008 45848 73020 45882
rect 72820 45836 73020 45848
rect 72820 45794 73020 45806
rect 72820 45760 72832 45794
rect 73008 45760 73020 45794
rect 72820 45748 73020 45760
rect 72820 45572 73020 45584
rect 72820 45538 72832 45572
rect 73008 45538 73020 45572
rect 72820 45526 73020 45538
rect 72820 45484 73020 45496
rect 72820 45450 72832 45484
rect 73008 45450 73020 45484
rect 72820 45438 73020 45450
rect 77810 45882 78010 45894
rect 77810 45848 77822 45882
rect 77998 45848 78010 45882
rect 77810 45836 78010 45848
rect 77810 45794 78010 45806
rect 77810 45760 77822 45794
rect 77998 45760 78010 45794
rect 77810 45748 78010 45760
rect 77810 45572 78010 45584
rect 77810 45538 77822 45572
rect 77998 45538 78010 45572
rect 77810 45526 78010 45538
rect 77810 45484 78010 45496
rect 77810 45450 77822 45484
rect 77998 45450 78010 45484
rect 77810 45438 78010 45450
rect 2960 44172 3160 44184
rect 2960 44138 2972 44172
rect 3148 44138 3160 44172
rect 2960 44126 3160 44138
rect 2960 44084 3160 44096
rect 2960 44050 2972 44084
rect 3148 44050 3160 44084
rect 2960 44038 3160 44050
rect 2960 43862 3160 43874
rect 2960 43828 2972 43862
rect 3148 43828 3160 43862
rect 2960 43816 3160 43828
rect 2960 43774 3160 43786
rect 2960 43740 2972 43774
rect 3148 43740 3160 43774
rect 2960 43728 3160 43740
rect 7950 44172 8150 44184
rect 7950 44138 7962 44172
rect 8138 44138 8150 44172
rect 7950 44126 8150 44138
rect 7950 44084 8150 44096
rect 7950 44050 7962 44084
rect 8138 44050 8150 44084
rect 7950 44038 8150 44050
rect 7950 43862 8150 43874
rect 7950 43828 7962 43862
rect 8138 43828 8150 43862
rect 7950 43816 8150 43828
rect 7950 43774 8150 43786
rect 7950 43740 7962 43774
rect 8138 43740 8150 43774
rect 7950 43728 8150 43740
rect 12940 44172 13140 44184
rect 12940 44138 12952 44172
rect 13128 44138 13140 44172
rect 12940 44126 13140 44138
rect 12940 44084 13140 44096
rect 12940 44050 12952 44084
rect 13128 44050 13140 44084
rect 12940 44038 13140 44050
rect 12940 43862 13140 43874
rect 12940 43828 12952 43862
rect 13128 43828 13140 43862
rect 12940 43816 13140 43828
rect 12940 43774 13140 43786
rect 12940 43740 12952 43774
rect 13128 43740 13140 43774
rect 12940 43728 13140 43740
rect 17930 44172 18130 44184
rect 17930 44138 17942 44172
rect 18118 44138 18130 44172
rect 17930 44126 18130 44138
rect 17930 44084 18130 44096
rect 17930 44050 17942 44084
rect 18118 44050 18130 44084
rect 17930 44038 18130 44050
rect 17930 43862 18130 43874
rect 17930 43828 17942 43862
rect 18118 43828 18130 43862
rect 17930 43816 18130 43828
rect 17930 43774 18130 43786
rect 17930 43740 17942 43774
rect 18118 43740 18130 43774
rect 17930 43728 18130 43740
rect 22920 44172 23120 44184
rect 22920 44138 22932 44172
rect 23108 44138 23120 44172
rect 22920 44126 23120 44138
rect 22920 44084 23120 44096
rect 22920 44050 22932 44084
rect 23108 44050 23120 44084
rect 22920 44038 23120 44050
rect 22920 43862 23120 43874
rect 22920 43828 22932 43862
rect 23108 43828 23120 43862
rect 22920 43816 23120 43828
rect 22920 43774 23120 43786
rect 22920 43740 22932 43774
rect 23108 43740 23120 43774
rect 22920 43728 23120 43740
rect 27910 44172 28110 44184
rect 27910 44138 27922 44172
rect 28098 44138 28110 44172
rect 27910 44126 28110 44138
rect 27910 44084 28110 44096
rect 27910 44050 27922 44084
rect 28098 44050 28110 44084
rect 27910 44038 28110 44050
rect 27910 43862 28110 43874
rect 27910 43828 27922 43862
rect 28098 43828 28110 43862
rect 27910 43816 28110 43828
rect 27910 43774 28110 43786
rect 27910 43740 27922 43774
rect 28098 43740 28110 43774
rect 27910 43728 28110 43740
rect 32900 44172 33100 44184
rect 32900 44138 32912 44172
rect 33088 44138 33100 44172
rect 32900 44126 33100 44138
rect 32900 44084 33100 44096
rect 32900 44050 32912 44084
rect 33088 44050 33100 44084
rect 32900 44038 33100 44050
rect 32900 43862 33100 43874
rect 32900 43828 32912 43862
rect 33088 43828 33100 43862
rect 32900 43816 33100 43828
rect 32900 43774 33100 43786
rect 32900 43740 32912 43774
rect 33088 43740 33100 43774
rect 32900 43728 33100 43740
rect 37890 44172 38090 44184
rect 37890 44138 37902 44172
rect 38078 44138 38090 44172
rect 37890 44126 38090 44138
rect 37890 44084 38090 44096
rect 37890 44050 37902 44084
rect 38078 44050 38090 44084
rect 37890 44038 38090 44050
rect 37890 43862 38090 43874
rect 37890 43828 37902 43862
rect 38078 43828 38090 43862
rect 37890 43816 38090 43828
rect 37890 43774 38090 43786
rect 37890 43740 37902 43774
rect 38078 43740 38090 43774
rect 37890 43728 38090 43740
rect 42880 44172 43080 44184
rect 42880 44138 42892 44172
rect 43068 44138 43080 44172
rect 42880 44126 43080 44138
rect 42880 44084 43080 44096
rect 42880 44050 42892 44084
rect 43068 44050 43080 44084
rect 42880 44038 43080 44050
rect 42880 43862 43080 43874
rect 42880 43828 42892 43862
rect 43068 43828 43080 43862
rect 42880 43816 43080 43828
rect 42880 43774 43080 43786
rect 42880 43740 42892 43774
rect 43068 43740 43080 43774
rect 42880 43728 43080 43740
rect 47870 44172 48070 44184
rect 47870 44138 47882 44172
rect 48058 44138 48070 44172
rect 47870 44126 48070 44138
rect 47870 44084 48070 44096
rect 47870 44050 47882 44084
rect 48058 44050 48070 44084
rect 47870 44038 48070 44050
rect 47870 43862 48070 43874
rect 47870 43828 47882 43862
rect 48058 43828 48070 43862
rect 47870 43816 48070 43828
rect 47870 43774 48070 43786
rect 47870 43740 47882 43774
rect 48058 43740 48070 43774
rect 47870 43728 48070 43740
rect 52860 44172 53060 44184
rect 52860 44138 52872 44172
rect 53048 44138 53060 44172
rect 52860 44126 53060 44138
rect 52860 44084 53060 44096
rect 52860 44050 52872 44084
rect 53048 44050 53060 44084
rect 52860 44038 53060 44050
rect 52860 43862 53060 43874
rect 52860 43828 52872 43862
rect 53048 43828 53060 43862
rect 52860 43816 53060 43828
rect 52860 43774 53060 43786
rect 52860 43740 52872 43774
rect 53048 43740 53060 43774
rect 52860 43728 53060 43740
rect 57850 44172 58050 44184
rect 57850 44138 57862 44172
rect 58038 44138 58050 44172
rect 57850 44126 58050 44138
rect 57850 44084 58050 44096
rect 57850 44050 57862 44084
rect 58038 44050 58050 44084
rect 57850 44038 58050 44050
rect 57850 43862 58050 43874
rect 57850 43828 57862 43862
rect 58038 43828 58050 43862
rect 57850 43816 58050 43828
rect 57850 43774 58050 43786
rect 57850 43740 57862 43774
rect 58038 43740 58050 43774
rect 57850 43728 58050 43740
rect 62840 44172 63040 44184
rect 62840 44138 62852 44172
rect 63028 44138 63040 44172
rect 62840 44126 63040 44138
rect 62840 44084 63040 44096
rect 62840 44050 62852 44084
rect 63028 44050 63040 44084
rect 62840 44038 63040 44050
rect 62840 43862 63040 43874
rect 62840 43828 62852 43862
rect 63028 43828 63040 43862
rect 62840 43816 63040 43828
rect 62840 43774 63040 43786
rect 62840 43740 62852 43774
rect 63028 43740 63040 43774
rect 62840 43728 63040 43740
rect 67830 44172 68030 44184
rect 67830 44138 67842 44172
rect 68018 44138 68030 44172
rect 67830 44126 68030 44138
rect 67830 44084 68030 44096
rect 67830 44050 67842 44084
rect 68018 44050 68030 44084
rect 67830 44038 68030 44050
rect 67830 43862 68030 43874
rect 67830 43828 67842 43862
rect 68018 43828 68030 43862
rect 67830 43816 68030 43828
rect 67830 43774 68030 43786
rect 67830 43740 67842 43774
rect 68018 43740 68030 43774
rect 67830 43728 68030 43740
rect 72820 44172 73020 44184
rect 72820 44138 72832 44172
rect 73008 44138 73020 44172
rect 72820 44126 73020 44138
rect 72820 44084 73020 44096
rect 72820 44050 72832 44084
rect 73008 44050 73020 44084
rect 72820 44038 73020 44050
rect 72820 43862 73020 43874
rect 72820 43828 72832 43862
rect 73008 43828 73020 43862
rect 72820 43816 73020 43828
rect 72820 43774 73020 43786
rect 72820 43740 72832 43774
rect 73008 43740 73020 43774
rect 72820 43728 73020 43740
rect 77810 44172 78010 44184
rect 77810 44138 77822 44172
rect 77998 44138 78010 44172
rect 77810 44126 78010 44138
rect 77810 44084 78010 44096
rect 77810 44050 77822 44084
rect 77998 44050 78010 44084
rect 77810 44038 78010 44050
rect 77810 43862 78010 43874
rect 77810 43828 77822 43862
rect 77998 43828 78010 43862
rect 77810 43816 78010 43828
rect 77810 43774 78010 43786
rect 77810 43740 77822 43774
rect 77998 43740 78010 43774
rect 77810 43728 78010 43740
rect 2960 42462 3160 42474
rect 2960 42428 2972 42462
rect 3148 42428 3160 42462
rect 2960 42416 3160 42428
rect 2960 42374 3160 42386
rect 2960 42340 2972 42374
rect 3148 42340 3160 42374
rect 2960 42328 3160 42340
rect 2960 42152 3160 42164
rect 2960 42118 2972 42152
rect 3148 42118 3160 42152
rect 2960 42106 3160 42118
rect 2960 42064 3160 42076
rect 2960 42030 2972 42064
rect 3148 42030 3160 42064
rect 2960 42018 3160 42030
rect 7950 42462 8150 42474
rect 7950 42428 7962 42462
rect 8138 42428 8150 42462
rect 7950 42416 8150 42428
rect 7950 42374 8150 42386
rect 7950 42340 7962 42374
rect 8138 42340 8150 42374
rect 7950 42328 8150 42340
rect 7950 42152 8150 42164
rect 7950 42118 7962 42152
rect 8138 42118 8150 42152
rect 7950 42106 8150 42118
rect 7950 42064 8150 42076
rect 7950 42030 7962 42064
rect 8138 42030 8150 42064
rect 7950 42018 8150 42030
rect 12940 42462 13140 42474
rect 12940 42428 12952 42462
rect 13128 42428 13140 42462
rect 12940 42416 13140 42428
rect 12940 42374 13140 42386
rect 12940 42340 12952 42374
rect 13128 42340 13140 42374
rect 12940 42328 13140 42340
rect 12940 42152 13140 42164
rect 12940 42118 12952 42152
rect 13128 42118 13140 42152
rect 12940 42106 13140 42118
rect 12940 42064 13140 42076
rect 12940 42030 12952 42064
rect 13128 42030 13140 42064
rect 12940 42018 13140 42030
rect 17930 42462 18130 42474
rect 17930 42428 17942 42462
rect 18118 42428 18130 42462
rect 17930 42416 18130 42428
rect 17930 42374 18130 42386
rect 17930 42340 17942 42374
rect 18118 42340 18130 42374
rect 17930 42328 18130 42340
rect 17930 42152 18130 42164
rect 17930 42118 17942 42152
rect 18118 42118 18130 42152
rect 17930 42106 18130 42118
rect 17930 42064 18130 42076
rect 17930 42030 17942 42064
rect 18118 42030 18130 42064
rect 17930 42018 18130 42030
rect 22920 42462 23120 42474
rect 22920 42428 22932 42462
rect 23108 42428 23120 42462
rect 22920 42416 23120 42428
rect 22920 42374 23120 42386
rect 22920 42340 22932 42374
rect 23108 42340 23120 42374
rect 22920 42328 23120 42340
rect 22920 42152 23120 42164
rect 22920 42118 22932 42152
rect 23108 42118 23120 42152
rect 22920 42106 23120 42118
rect 22920 42064 23120 42076
rect 22920 42030 22932 42064
rect 23108 42030 23120 42064
rect 22920 42018 23120 42030
rect 27910 42462 28110 42474
rect 27910 42428 27922 42462
rect 28098 42428 28110 42462
rect 27910 42416 28110 42428
rect 27910 42374 28110 42386
rect 27910 42340 27922 42374
rect 28098 42340 28110 42374
rect 27910 42328 28110 42340
rect 27910 42152 28110 42164
rect 27910 42118 27922 42152
rect 28098 42118 28110 42152
rect 27910 42106 28110 42118
rect 27910 42064 28110 42076
rect 27910 42030 27922 42064
rect 28098 42030 28110 42064
rect 27910 42018 28110 42030
rect 32900 42462 33100 42474
rect 32900 42428 32912 42462
rect 33088 42428 33100 42462
rect 32900 42416 33100 42428
rect 32900 42374 33100 42386
rect 32900 42340 32912 42374
rect 33088 42340 33100 42374
rect 32900 42328 33100 42340
rect 32900 42152 33100 42164
rect 32900 42118 32912 42152
rect 33088 42118 33100 42152
rect 32900 42106 33100 42118
rect 32900 42064 33100 42076
rect 32900 42030 32912 42064
rect 33088 42030 33100 42064
rect 32900 42018 33100 42030
rect 37890 42462 38090 42474
rect 37890 42428 37902 42462
rect 38078 42428 38090 42462
rect 37890 42416 38090 42428
rect 37890 42374 38090 42386
rect 37890 42340 37902 42374
rect 38078 42340 38090 42374
rect 37890 42328 38090 42340
rect 37890 42152 38090 42164
rect 37890 42118 37902 42152
rect 38078 42118 38090 42152
rect 37890 42106 38090 42118
rect 37890 42064 38090 42076
rect 37890 42030 37902 42064
rect 38078 42030 38090 42064
rect 37890 42018 38090 42030
rect 42880 42462 43080 42474
rect 42880 42428 42892 42462
rect 43068 42428 43080 42462
rect 42880 42416 43080 42428
rect 42880 42374 43080 42386
rect 42880 42340 42892 42374
rect 43068 42340 43080 42374
rect 42880 42328 43080 42340
rect 42880 42152 43080 42164
rect 42880 42118 42892 42152
rect 43068 42118 43080 42152
rect 42880 42106 43080 42118
rect 42880 42064 43080 42076
rect 42880 42030 42892 42064
rect 43068 42030 43080 42064
rect 42880 42018 43080 42030
rect 47870 42462 48070 42474
rect 47870 42428 47882 42462
rect 48058 42428 48070 42462
rect 47870 42416 48070 42428
rect 47870 42374 48070 42386
rect 47870 42340 47882 42374
rect 48058 42340 48070 42374
rect 47870 42328 48070 42340
rect 47870 42152 48070 42164
rect 47870 42118 47882 42152
rect 48058 42118 48070 42152
rect 47870 42106 48070 42118
rect 47870 42064 48070 42076
rect 47870 42030 47882 42064
rect 48058 42030 48070 42064
rect 47870 42018 48070 42030
rect 52860 42462 53060 42474
rect 52860 42428 52872 42462
rect 53048 42428 53060 42462
rect 52860 42416 53060 42428
rect 52860 42374 53060 42386
rect 52860 42340 52872 42374
rect 53048 42340 53060 42374
rect 52860 42328 53060 42340
rect 52860 42152 53060 42164
rect 52860 42118 52872 42152
rect 53048 42118 53060 42152
rect 52860 42106 53060 42118
rect 52860 42064 53060 42076
rect 52860 42030 52872 42064
rect 53048 42030 53060 42064
rect 52860 42018 53060 42030
rect 57850 42462 58050 42474
rect 57850 42428 57862 42462
rect 58038 42428 58050 42462
rect 57850 42416 58050 42428
rect 57850 42374 58050 42386
rect 57850 42340 57862 42374
rect 58038 42340 58050 42374
rect 57850 42328 58050 42340
rect 57850 42152 58050 42164
rect 57850 42118 57862 42152
rect 58038 42118 58050 42152
rect 57850 42106 58050 42118
rect 57850 42064 58050 42076
rect 57850 42030 57862 42064
rect 58038 42030 58050 42064
rect 57850 42018 58050 42030
rect 62840 42462 63040 42474
rect 62840 42428 62852 42462
rect 63028 42428 63040 42462
rect 62840 42416 63040 42428
rect 62840 42374 63040 42386
rect 62840 42340 62852 42374
rect 63028 42340 63040 42374
rect 62840 42328 63040 42340
rect 62840 42152 63040 42164
rect 62840 42118 62852 42152
rect 63028 42118 63040 42152
rect 62840 42106 63040 42118
rect 62840 42064 63040 42076
rect 62840 42030 62852 42064
rect 63028 42030 63040 42064
rect 62840 42018 63040 42030
rect 67830 42462 68030 42474
rect 67830 42428 67842 42462
rect 68018 42428 68030 42462
rect 67830 42416 68030 42428
rect 67830 42374 68030 42386
rect 67830 42340 67842 42374
rect 68018 42340 68030 42374
rect 67830 42328 68030 42340
rect 67830 42152 68030 42164
rect 67830 42118 67842 42152
rect 68018 42118 68030 42152
rect 67830 42106 68030 42118
rect 67830 42064 68030 42076
rect 67830 42030 67842 42064
rect 68018 42030 68030 42064
rect 67830 42018 68030 42030
rect 72820 42462 73020 42474
rect 72820 42428 72832 42462
rect 73008 42428 73020 42462
rect 72820 42416 73020 42428
rect 72820 42374 73020 42386
rect 72820 42340 72832 42374
rect 73008 42340 73020 42374
rect 72820 42328 73020 42340
rect 72820 42152 73020 42164
rect 72820 42118 72832 42152
rect 73008 42118 73020 42152
rect 72820 42106 73020 42118
rect 72820 42064 73020 42076
rect 72820 42030 72832 42064
rect 73008 42030 73020 42064
rect 72820 42018 73020 42030
rect 77810 42462 78010 42474
rect 77810 42428 77822 42462
rect 77998 42428 78010 42462
rect 77810 42416 78010 42428
rect 77810 42374 78010 42386
rect 77810 42340 77822 42374
rect 77998 42340 78010 42374
rect 77810 42328 78010 42340
rect 77810 42152 78010 42164
rect 77810 42118 77822 42152
rect 77998 42118 78010 42152
rect 77810 42106 78010 42118
rect 77810 42064 78010 42076
rect 77810 42030 77822 42064
rect 77998 42030 78010 42064
rect 77810 42018 78010 42030
rect 2960 40752 3160 40764
rect 2960 40718 2972 40752
rect 3148 40718 3160 40752
rect 2960 40706 3160 40718
rect 2960 40664 3160 40676
rect 2960 40630 2972 40664
rect 3148 40630 3160 40664
rect 2960 40618 3160 40630
rect 2960 40442 3160 40454
rect 2960 40408 2972 40442
rect 3148 40408 3160 40442
rect 2960 40396 3160 40408
rect 2960 40354 3160 40366
rect 2960 40320 2972 40354
rect 3148 40320 3160 40354
rect 2960 40308 3160 40320
rect 7950 40752 8150 40764
rect 7950 40718 7962 40752
rect 8138 40718 8150 40752
rect 7950 40706 8150 40718
rect 7950 40664 8150 40676
rect 7950 40630 7962 40664
rect 8138 40630 8150 40664
rect 7950 40618 8150 40630
rect 7950 40442 8150 40454
rect 7950 40408 7962 40442
rect 8138 40408 8150 40442
rect 7950 40396 8150 40408
rect 7950 40354 8150 40366
rect 7950 40320 7962 40354
rect 8138 40320 8150 40354
rect 7950 40308 8150 40320
rect 12940 40752 13140 40764
rect 12940 40718 12952 40752
rect 13128 40718 13140 40752
rect 12940 40706 13140 40718
rect 12940 40664 13140 40676
rect 12940 40630 12952 40664
rect 13128 40630 13140 40664
rect 12940 40618 13140 40630
rect 12940 40442 13140 40454
rect 12940 40408 12952 40442
rect 13128 40408 13140 40442
rect 12940 40396 13140 40408
rect 12940 40354 13140 40366
rect 12940 40320 12952 40354
rect 13128 40320 13140 40354
rect 12940 40308 13140 40320
rect 17930 40752 18130 40764
rect 17930 40718 17942 40752
rect 18118 40718 18130 40752
rect 17930 40706 18130 40718
rect 17930 40664 18130 40676
rect 17930 40630 17942 40664
rect 18118 40630 18130 40664
rect 17930 40618 18130 40630
rect 17930 40442 18130 40454
rect 17930 40408 17942 40442
rect 18118 40408 18130 40442
rect 17930 40396 18130 40408
rect 17930 40354 18130 40366
rect 17930 40320 17942 40354
rect 18118 40320 18130 40354
rect 17930 40308 18130 40320
rect 22920 40752 23120 40764
rect 22920 40718 22932 40752
rect 23108 40718 23120 40752
rect 22920 40706 23120 40718
rect 22920 40664 23120 40676
rect 22920 40630 22932 40664
rect 23108 40630 23120 40664
rect 22920 40618 23120 40630
rect 22920 40442 23120 40454
rect 22920 40408 22932 40442
rect 23108 40408 23120 40442
rect 22920 40396 23120 40408
rect 22920 40354 23120 40366
rect 22920 40320 22932 40354
rect 23108 40320 23120 40354
rect 22920 40308 23120 40320
rect 27910 40752 28110 40764
rect 27910 40718 27922 40752
rect 28098 40718 28110 40752
rect 27910 40706 28110 40718
rect 27910 40664 28110 40676
rect 27910 40630 27922 40664
rect 28098 40630 28110 40664
rect 27910 40618 28110 40630
rect 27910 40442 28110 40454
rect 27910 40408 27922 40442
rect 28098 40408 28110 40442
rect 27910 40396 28110 40408
rect 27910 40354 28110 40366
rect 27910 40320 27922 40354
rect 28098 40320 28110 40354
rect 27910 40308 28110 40320
rect 32900 40752 33100 40764
rect 32900 40718 32912 40752
rect 33088 40718 33100 40752
rect 32900 40706 33100 40718
rect 32900 40664 33100 40676
rect 32900 40630 32912 40664
rect 33088 40630 33100 40664
rect 32900 40618 33100 40630
rect 32900 40442 33100 40454
rect 32900 40408 32912 40442
rect 33088 40408 33100 40442
rect 32900 40396 33100 40408
rect 32900 40354 33100 40366
rect 32900 40320 32912 40354
rect 33088 40320 33100 40354
rect 32900 40308 33100 40320
rect 37890 40752 38090 40764
rect 37890 40718 37902 40752
rect 38078 40718 38090 40752
rect 37890 40706 38090 40718
rect 37890 40664 38090 40676
rect 37890 40630 37902 40664
rect 38078 40630 38090 40664
rect 37890 40618 38090 40630
rect 37890 40442 38090 40454
rect 37890 40408 37902 40442
rect 38078 40408 38090 40442
rect 37890 40396 38090 40408
rect 37890 40354 38090 40366
rect 37890 40320 37902 40354
rect 38078 40320 38090 40354
rect 37890 40308 38090 40320
rect 42880 40752 43080 40764
rect 42880 40718 42892 40752
rect 43068 40718 43080 40752
rect 42880 40706 43080 40718
rect 42880 40664 43080 40676
rect 42880 40630 42892 40664
rect 43068 40630 43080 40664
rect 42880 40618 43080 40630
rect 42880 40442 43080 40454
rect 42880 40408 42892 40442
rect 43068 40408 43080 40442
rect 42880 40396 43080 40408
rect 42880 40354 43080 40366
rect 42880 40320 42892 40354
rect 43068 40320 43080 40354
rect 42880 40308 43080 40320
rect 47870 40752 48070 40764
rect 47870 40718 47882 40752
rect 48058 40718 48070 40752
rect 47870 40706 48070 40718
rect 47870 40664 48070 40676
rect 47870 40630 47882 40664
rect 48058 40630 48070 40664
rect 47870 40618 48070 40630
rect 47870 40442 48070 40454
rect 47870 40408 47882 40442
rect 48058 40408 48070 40442
rect 47870 40396 48070 40408
rect 47870 40354 48070 40366
rect 47870 40320 47882 40354
rect 48058 40320 48070 40354
rect 47870 40308 48070 40320
rect 52860 40752 53060 40764
rect 52860 40718 52872 40752
rect 53048 40718 53060 40752
rect 52860 40706 53060 40718
rect 52860 40664 53060 40676
rect 52860 40630 52872 40664
rect 53048 40630 53060 40664
rect 52860 40618 53060 40630
rect 52860 40442 53060 40454
rect 52860 40408 52872 40442
rect 53048 40408 53060 40442
rect 52860 40396 53060 40408
rect 52860 40354 53060 40366
rect 52860 40320 52872 40354
rect 53048 40320 53060 40354
rect 52860 40308 53060 40320
rect 57850 40752 58050 40764
rect 57850 40718 57862 40752
rect 58038 40718 58050 40752
rect 57850 40706 58050 40718
rect 57850 40664 58050 40676
rect 57850 40630 57862 40664
rect 58038 40630 58050 40664
rect 57850 40618 58050 40630
rect 57850 40442 58050 40454
rect 57850 40408 57862 40442
rect 58038 40408 58050 40442
rect 57850 40396 58050 40408
rect 57850 40354 58050 40366
rect 57850 40320 57862 40354
rect 58038 40320 58050 40354
rect 57850 40308 58050 40320
rect 62840 40752 63040 40764
rect 62840 40718 62852 40752
rect 63028 40718 63040 40752
rect 62840 40706 63040 40718
rect 62840 40664 63040 40676
rect 62840 40630 62852 40664
rect 63028 40630 63040 40664
rect 62840 40618 63040 40630
rect 62840 40442 63040 40454
rect 62840 40408 62852 40442
rect 63028 40408 63040 40442
rect 62840 40396 63040 40408
rect 62840 40354 63040 40366
rect 62840 40320 62852 40354
rect 63028 40320 63040 40354
rect 62840 40308 63040 40320
rect 67830 40752 68030 40764
rect 67830 40718 67842 40752
rect 68018 40718 68030 40752
rect 67830 40706 68030 40718
rect 67830 40664 68030 40676
rect 67830 40630 67842 40664
rect 68018 40630 68030 40664
rect 67830 40618 68030 40630
rect 67830 40442 68030 40454
rect 67830 40408 67842 40442
rect 68018 40408 68030 40442
rect 67830 40396 68030 40408
rect 67830 40354 68030 40366
rect 67830 40320 67842 40354
rect 68018 40320 68030 40354
rect 67830 40308 68030 40320
rect 72820 40752 73020 40764
rect 72820 40718 72832 40752
rect 73008 40718 73020 40752
rect 72820 40706 73020 40718
rect 72820 40664 73020 40676
rect 72820 40630 72832 40664
rect 73008 40630 73020 40664
rect 72820 40618 73020 40630
rect 72820 40442 73020 40454
rect 72820 40408 72832 40442
rect 73008 40408 73020 40442
rect 72820 40396 73020 40408
rect 72820 40354 73020 40366
rect 72820 40320 72832 40354
rect 73008 40320 73020 40354
rect 72820 40308 73020 40320
rect 77810 40752 78010 40764
rect 77810 40718 77822 40752
rect 77998 40718 78010 40752
rect 77810 40706 78010 40718
rect 77810 40664 78010 40676
rect 77810 40630 77822 40664
rect 77998 40630 78010 40664
rect 77810 40618 78010 40630
rect 77810 40442 78010 40454
rect 77810 40408 77822 40442
rect 77998 40408 78010 40442
rect 77810 40396 78010 40408
rect 77810 40354 78010 40366
rect 77810 40320 77822 40354
rect 77998 40320 78010 40354
rect 77810 40308 78010 40320
<< pdiff >>
rect 3458 66402 3658 66414
rect 3458 66368 3470 66402
rect 3646 66368 3658 66402
rect 3458 66356 3658 66368
rect 3458 66314 3658 66326
rect 3458 66280 3470 66314
rect 3646 66280 3658 66314
rect 3458 66268 3658 66280
rect 3458 66092 3658 66104
rect 3458 66058 3470 66092
rect 3646 66058 3658 66092
rect 3458 66046 3658 66058
rect 3458 66004 3658 66016
rect 3458 65970 3470 66004
rect 3646 65970 3658 66004
rect 3458 65958 3658 65970
rect 8448 66402 8648 66414
rect 8448 66368 8460 66402
rect 8636 66368 8648 66402
rect 8448 66356 8648 66368
rect 8448 66314 8648 66326
rect 8448 66280 8460 66314
rect 8636 66280 8648 66314
rect 8448 66268 8648 66280
rect 8448 66092 8648 66104
rect 8448 66058 8460 66092
rect 8636 66058 8648 66092
rect 8448 66046 8648 66058
rect 8448 66004 8648 66016
rect 8448 65970 8460 66004
rect 8636 65970 8648 66004
rect 8448 65958 8648 65970
rect 13438 66402 13638 66414
rect 13438 66368 13450 66402
rect 13626 66368 13638 66402
rect 13438 66356 13638 66368
rect 13438 66314 13638 66326
rect 13438 66280 13450 66314
rect 13626 66280 13638 66314
rect 13438 66268 13638 66280
rect 13438 66092 13638 66104
rect 13438 66058 13450 66092
rect 13626 66058 13638 66092
rect 13438 66046 13638 66058
rect 13438 66004 13638 66016
rect 13438 65970 13450 66004
rect 13626 65970 13638 66004
rect 13438 65958 13638 65970
rect 18428 66402 18628 66414
rect 18428 66368 18440 66402
rect 18616 66368 18628 66402
rect 18428 66356 18628 66368
rect 18428 66314 18628 66326
rect 18428 66280 18440 66314
rect 18616 66280 18628 66314
rect 18428 66268 18628 66280
rect 18428 66092 18628 66104
rect 18428 66058 18440 66092
rect 18616 66058 18628 66092
rect 18428 66046 18628 66058
rect 18428 66004 18628 66016
rect 18428 65970 18440 66004
rect 18616 65970 18628 66004
rect 18428 65958 18628 65970
rect 23418 66402 23618 66414
rect 23418 66368 23430 66402
rect 23606 66368 23618 66402
rect 23418 66356 23618 66368
rect 23418 66314 23618 66326
rect 23418 66280 23430 66314
rect 23606 66280 23618 66314
rect 23418 66268 23618 66280
rect 23418 66092 23618 66104
rect 23418 66058 23430 66092
rect 23606 66058 23618 66092
rect 23418 66046 23618 66058
rect 23418 66004 23618 66016
rect 23418 65970 23430 66004
rect 23606 65970 23618 66004
rect 23418 65958 23618 65970
rect 28408 66402 28608 66414
rect 28408 66368 28420 66402
rect 28596 66368 28608 66402
rect 28408 66356 28608 66368
rect 28408 66314 28608 66326
rect 28408 66280 28420 66314
rect 28596 66280 28608 66314
rect 28408 66268 28608 66280
rect 28408 66092 28608 66104
rect 28408 66058 28420 66092
rect 28596 66058 28608 66092
rect 28408 66046 28608 66058
rect 28408 66004 28608 66016
rect 28408 65970 28420 66004
rect 28596 65970 28608 66004
rect 28408 65958 28608 65970
rect 33398 66402 33598 66414
rect 33398 66368 33410 66402
rect 33586 66368 33598 66402
rect 33398 66356 33598 66368
rect 33398 66314 33598 66326
rect 33398 66280 33410 66314
rect 33586 66280 33598 66314
rect 33398 66268 33598 66280
rect 33398 66092 33598 66104
rect 33398 66058 33410 66092
rect 33586 66058 33598 66092
rect 33398 66046 33598 66058
rect 33398 66004 33598 66016
rect 33398 65970 33410 66004
rect 33586 65970 33598 66004
rect 33398 65958 33598 65970
rect 38388 66402 38588 66414
rect 38388 66368 38400 66402
rect 38576 66368 38588 66402
rect 38388 66356 38588 66368
rect 38388 66314 38588 66326
rect 38388 66280 38400 66314
rect 38576 66280 38588 66314
rect 38388 66268 38588 66280
rect 38388 66092 38588 66104
rect 38388 66058 38400 66092
rect 38576 66058 38588 66092
rect 38388 66046 38588 66058
rect 38388 66004 38588 66016
rect 38388 65970 38400 66004
rect 38576 65970 38588 66004
rect 38388 65958 38588 65970
rect 43378 66402 43578 66414
rect 43378 66368 43390 66402
rect 43566 66368 43578 66402
rect 43378 66356 43578 66368
rect 43378 66314 43578 66326
rect 43378 66280 43390 66314
rect 43566 66280 43578 66314
rect 43378 66268 43578 66280
rect 43378 66092 43578 66104
rect 43378 66058 43390 66092
rect 43566 66058 43578 66092
rect 43378 66046 43578 66058
rect 43378 66004 43578 66016
rect 43378 65970 43390 66004
rect 43566 65970 43578 66004
rect 43378 65958 43578 65970
rect 48368 66402 48568 66414
rect 48368 66368 48380 66402
rect 48556 66368 48568 66402
rect 48368 66356 48568 66368
rect 48368 66314 48568 66326
rect 48368 66280 48380 66314
rect 48556 66280 48568 66314
rect 48368 66268 48568 66280
rect 48368 66092 48568 66104
rect 48368 66058 48380 66092
rect 48556 66058 48568 66092
rect 48368 66046 48568 66058
rect 48368 66004 48568 66016
rect 48368 65970 48380 66004
rect 48556 65970 48568 66004
rect 48368 65958 48568 65970
rect 53358 66402 53558 66414
rect 53358 66368 53370 66402
rect 53546 66368 53558 66402
rect 53358 66356 53558 66368
rect 53358 66314 53558 66326
rect 53358 66280 53370 66314
rect 53546 66280 53558 66314
rect 53358 66268 53558 66280
rect 53358 66092 53558 66104
rect 53358 66058 53370 66092
rect 53546 66058 53558 66092
rect 53358 66046 53558 66058
rect 53358 66004 53558 66016
rect 53358 65970 53370 66004
rect 53546 65970 53558 66004
rect 53358 65958 53558 65970
rect 58348 66402 58548 66414
rect 58348 66368 58360 66402
rect 58536 66368 58548 66402
rect 58348 66356 58548 66368
rect 58348 66314 58548 66326
rect 58348 66280 58360 66314
rect 58536 66280 58548 66314
rect 58348 66268 58548 66280
rect 58348 66092 58548 66104
rect 58348 66058 58360 66092
rect 58536 66058 58548 66092
rect 58348 66046 58548 66058
rect 58348 66004 58548 66016
rect 58348 65970 58360 66004
rect 58536 65970 58548 66004
rect 58348 65958 58548 65970
rect 63338 66402 63538 66414
rect 63338 66368 63350 66402
rect 63526 66368 63538 66402
rect 63338 66356 63538 66368
rect 63338 66314 63538 66326
rect 63338 66280 63350 66314
rect 63526 66280 63538 66314
rect 63338 66268 63538 66280
rect 63338 66092 63538 66104
rect 63338 66058 63350 66092
rect 63526 66058 63538 66092
rect 63338 66046 63538 66058
rect 63338 66004 63538 66016
rect 63338 65970 63350 66004
rect 63526 65970 63538 66004
rect 63338 65958 63538 65970
rect 68328 66402 68528 66414
rect 68328 66368 68340 66402
rect 68516 66368 68528 66402
rect 68328 66356 68528 66368
rect 68328 66314 68528 66326
rect 68328 66280 68340 66314
rect 68516 66280 68528 66314
rect 68328 66268 68528 66280
rect 68328 66092 68528 66104
rect 68328 66058 68340 66092
rect 68516 66058 68528 66092
rect 68328 66046 68528 66058
rect 68328 66004 68528 66016
rect 68328 65970 68340 66004
rect 68516 65970 68528 66004
rect 68328 65958 68528 65970
rect 73318 66402 73518 66414
rect 73318 66368 73330 66402
rect 73506 66368 73518 66402
rect 73318 66356 73518 66368
rect 73318 66314 73518 66326
rect 73318 66280 73330 66314
rect 73506 66280 73518 66314
rect 73318 66268 73518 66280
rect 73318 66092 73518 66104
rect 73318 66058 73330 66092
rect 73506 66058 73518 66092
rect 73318 66046 73518 66058
rect 73318 66004 73518 66016
rect 73318 65970 73330 66004
rect 73506 65970 73518 66004
rect 73318 65958 73518 65970
rect 78308 66402 78508 66414
rect 78308 66368 78320 66402
rect 78496 66368 78508 66402
rect 78308 66356 78508 66368
rect 78308 66314 78508 66326
rect 78308 66280 78320 66314
rect 78496 66280 78508 66314
rect 78308 66268 78508 66280
rect 78308 66092 78508 66104
rect 78308 66058 78320 66092
rect 78496 66058 78508 66092
rect 78308 66046 78508 66058
rect 78308 66004 78508 66016
rect 78308 65970 78320 66004
rect 78496 65970 78508 66004
rect 78308 65958 78508 65970
rect 3458 64692 3658 64704
rect 3458 64658 3470 64692
rect 3646 64658 3658 64692
rect 3458 64646 3658 64658
rect 3458 64604 3658 64616
rect 3458 64570 3470 64604
rect 3646 64570 3658 64604
rect 3458 64558 3658 64570
rect 3458 64382 3658 64394
rect 3458 64348 3470 64382
rect 3646 64348 3658 64382
rect 3458 64336 3658 64348
rect 3458 64294 3658 64306
rect 3458 64260 3470 64294
rect 3646 64260 3658 64294
rect 3458 64248 3658 64260
rect 8448 64692 8648 64704
rect 8448 64658 8460 64692
rect 8636 64658 8648 64692
rect 8448 64646 8648 64658
rect 8448 64604 8648 64616
rect 8448 64570 8460 64604
rect 8636 64570 8648 64604
rect 8448 64558 8648 64570
rect 8448 64382 8648 64394
rect 8448 64348 8460 64382
rect 8636 64348 8648 64382
rect 8448 64336 8648 64348
rect 8448 64294 8648 64306
rect 8448 64260 8460 64294
rect 8636 64260 8648 64294
rect 8448 64248 8648 64260
rect 13438 64692 13638 64704
rect 13438 64658 13450 64692
rect 13626 64658 13638 64692
rect 13438 64646 13638 64658
rect 13438 64604 13638 64616
rect 13438 64570 13450 64604
rect 13626 64570 13638 64604
rect 13438 64558 13638 64570
rect 13438 64382 13638 64394
rect 13438 64348 13450 64382
rect 13626 64348 13638 64382
rect 13438 64336 13638 64348
rect 13438 64294 13638 64306
rect 13438 64260 13450 64294
rect 13626 64260 13638 64294
rect 13438 64248 13638 64260
rect 18428 64692 18628 64704
rect 18428 64658 18440 64692
rect 18616 64658 18628 64692
rect 18428 64646 18628 64658
rect 18428 64604 18628 64616
rect 18428 64570 18440 64604
rect 18616 64570 18628 64604
rect 18428 64558 18628 64570
rect 18428 64382 18628 64394
rect 18428 64348 18440 64382
rect 18616 64348 18628 64382
rect 18428 64336 18628 64348
rect 18428 64294 18628 64306
rect 18428 64260 18440 64294
rect 18616 64260 18628 64294
rect 18428 64248 18628 64260
rect 23418 64692 23618 64704
rect 23418 64658 23430 64692
rect 23606 64658 23618 64692
rect 23418 64646 23618 64658
rect 23418 64604 23618 64616
rect 23418 64570 23430 64604
rect 23606 64570 23618 64604
rect 23418 64558 23618 64570
rect 23418 64382 23618 64394
rect 23418 64348 23430 64382
rect 23606 64348 23618 64382
rect 23418 64336 23618 64348
rect 23418 64294 23618 64306
rect 23418 64260 23430 64294
rect 23606 64260 23618 64294
rect 23418 64248 23618 64260
rect 28408 64692 28608 64704
rect 28408 64658 28420 64692
rect 28596 64658 28608 64692
rect 28408 64646 28608 64658
rect 28408 64604 28608 64616
rect 28408 64570 28420 64604
rect 28596 64570 28608 64604
rect 28408 64558 28608 64570
rect 28408 64382 28608 64394
rect 28408 64348 28420 64382
rect 28596 64348 28608 64382
rect 28408 64336 28608 64348
rect 28408 64294 28608 64306
rect 28408 64260 28420 64294
rect 28596 64260 28608 64294
rect 28408 64248 28608 64260
rect 33398 64692 33598 64704
rect 33398 64658 33410 64692
rect 33586 64658 33598 64692
rect 33398 64646 33598 64658
rect 33398 64604 33598 64616
rect 33398 64570 33410 64604
rect 33586 64570 33598 64604
rect 33398 64558 33598 64570
rect 33398 64382 33598 64394
rect 33398 64348 33410 64382
rect 33586 64348 33598 64382
rect 33398 64336 33598 64348
rect 33398 64294 33598 64306
rect 33398 64260 33410 64294
rect 33586 64260 33598 64294
rect 33398 64248 33598 64260
rect 38388 64692 38588 64704
rect 38388 64658 38400 64692
rect 38576 64658 38588 64692
rect 38388 64646 38588 64658
rect 38388 64604 38588 64616
rect 38388 64570 38400 64604
rect 38576 64570 38588 64604
rect 38388 64558 38588 64570
rect 38388 64382 38588 64394
rect 38388 64348 38400 64382
rect 38576 64348 38588 64382
rect 38388 64336 38588 64348
rect 38388 64294 38588 64306
rect 38388 64260 38400 64294
rect 38576 64260 38588 64294
rect 38388 64248 38588 64260
rect 43378 64692 43578 64704
rect 43378 64658 43390 64692
rect 43566 64658 43578 64692
rect 43378 64646 43578 64658
rect 43378 64604 43578 64616
rect 43378 64570 43390 64604
rect 43566 64570 43578 64604
rect 43378 64558 43578 64570
rect 43378 64382 43578 64394
rect 43378 64348 43390 64382
rect 43566 64348 43578 64382
rect 43378 64336 43578 64348
rect 43378 64294 43578 64306
rect 43378 64260 43390 64294
rect 43566 64260 43578 64294
rect 43378 64248 43578 64260
rect 48368 64692 48568 64704
rect 48368 64658 48380 64692
rect 48556 64658 48568 64692
rect 48368 64646 48568 64658
rect 48368 64604 48568 64616
rect 48368 64570 48380 64604
rect 48556 64570 48568 64604
rect 48368 64558 48568 64570
rect 48368 64382 48568 64394
rect 48368 64348 48380 64382
rect 48556 64348 48568 64382
rect 48368 64336 48568 64348
rect 48368 64294 48568 64306
rect 48368 64260 48380 64294
rect 48556 64260 48568 64294
rect 48368 64248 48568 64260
rect 53358 64692 53558 64704
rect 53358 64658 53370 64692
rect 53546 64658 53558 64692
rect 53358 64646 53558 64658
rect 53358 64604 53558 64616
rect 53358 64570 53370 64604
rect 53546 64570 53558 64604
rect 53358 64558 53558 64570
rect 53358 64382 53558 64394
rect 53358 64348 53370 64382
rect 53546 64348 53558 64382
rect 53358 64336 53558 64348
rect 53358 64294 53558 64306
rect 53358 64260 53370 64294
rect 53546 64260 53558 64294
rect 53358 64248 53558 64260
rect 58348 64692 58548 64704
rect 58348 64658 58360 64692
rect 58536 64658 58548 64692
rect 58348 64646 58548 64658
rect 58348 64604 58548 64616
rect 58348 64570 58360 64604
rect 58536 64570 58548 64604
rect 58348 64558 58548 64570
rect 58348 64382 58548 64394
rect 58348 64348 58360 64382
rect 58536 64348 58548 64382
rect 58348 64336 58548 64348
rect 58348 64294 58548 64306
rect 58348 64260 58360 64294
rect 58536 64260 58548 64294
rect 58348 64248 58548 64260
rect 63338 64692 63538 64704
rect 63338 64658 63350 64692
rect 63526 64658 63538 64692
rect 63338 64646 63538 64658
rect 63338 64604 63538 64616
rect 63338 64570 63350 64604
rect 63526 64570 63538 64604
rect 63338 64558 63538 64570
rect 63338 64382 63538 64394
rect 63338 64348 63350 64382
rect 63526 64348 63538 64382
rect 63338 64336 63538 64348
rect 63338 64294 63538 64306
rect 63338 64260 63350 64294
rect 63526 64260 63538 64294
rect 63338 64248 63538 64260
rect 68328 64692 68528 64704
rect 68328 64658 68340 64692
rect 68516 64658 68528 64692
rect 68328 64646 68528 64658
rect 68328 64604 68528 64616
rect 68328 64570 68340 64604
rect 68516 64570 68528 64604
rect 68328 64558 68528 64570
rect 68328 64382 68528 64394
rect 68328 64348 68340 64382
rect 68516 64348 68528 64382
rect 68328 64336 68528 64348
rect 68328 64294 68528 64306
rect 68328 64260 68340 64294
rect 68516 64260 68528 64294
rect 68328 64248 68528 64260
rect 73318 64692 73518 64704
rect 73318 64658 73330 64692
rect 73506 64658 73518 64692
rect 73318 64646 73518 64658
rect 73318 64604 73518 64616
rect 73318 64570 73330 64604
rect 73506 64570 73518 64604
rect 73318 64558 73518 64570
rect 73318 64382 73518 64394
rect 73318 64348 73330 64382
rect 73506 64348 73518 64382
rect 73318 64336 73518 64348
rect 73318 64294 73518 64306
rect 73318 64260 73330 64294
rect 73506 64260 73518 64294
rect 73318 64248 73518 64260
rect 78308 64692 78508 64704
rect 78308 64658 78320 64692
rect 78496 64658 78508 64692
rect 78308 64646 78508 64658
rect 78308 64604 78508 64616
rect 78308 64570 78320 64604
rect 78496 64570 78508 64604
rect 78308 64558 78508 64570
rect 78308 64382 78508 64394
rect 78308 64348 78320 64382
rect 78496 64348 78508 64382
rect 78308 64336 78508 64348
rect 78308 64294 78508 64306
rect 78308 64260 78320 64294
rect 78496 64260 78508 64294
rect 78308 64248 78508 64260
rect 3458 62982 3658 62994
rect 3458 62948 3470 62982
rect 3646 62948 3658 62982
rect 3458 62936 3658 62948
rect 3458 62894 3658 62906
rect 3458 62860 3470 62894
rect 3646 62860 3658 62894
rect 3458 62848 3658 62860
rect 3458 62672 3658 62684
rect 3458 62638 3470 62672
rect 3646 62638 3658 62672
rect 3458 62626 3658 62638
rect 3458 62584 3658 62596
rect 3458 62550 3470 62584
rect 3646 62550 3658 62584
rect 3458 62538 3658 62550
rect 8448 62982 8648 62994
rect 8448 62948 8460 62982
rect 8636 62948 8648 62982
rect 8448 62936 8648 62948
rect 8448 62894 8648 62906
rect 8448 62860 8460 62894
rect 8636 62860 8648 62894
rect 8448 62848 8648 62860
rect 8448 62672 8648 62684
rect 8448 62638 8460 62672
rect 8636 62638 8648 62672
rect 8448 62626 8648 62638
rect 8448 62584 8648 62596
rect 8448 62550 8460 62584
rect 8636 62550 8648 62584
rect 8448 62538 8648 62550
rect 13438 62982 13638 62994
rect 13438 62948 13450 62982
rect 13626 62948 13638 62982
rect 13438 62936 13638 62948
rect 13438 62894 13638 62906
rect 13438 62860 13450 62894
rect 13626 62860 13638 62894
rect 13438 62848 13638 62860
rect 13438 62672 13638 62684
rect 13438 62638 13450 62672
rect 13626 62638 13638 62672
rect 13438 62626 13638 62638
rect 13438 62584 13638 62596
rect 13438 62550 13450 62584
rect 13626 62550 13638 62584
rect 13438 62538 13638 62550
rect 18428 62982 18628 62994
rect 18428 62948 18440 62982
rect 18616 62948 18628 62982
rect 18428 62936 18628 62948
rect 18428 62894 18628 62906
rect 18428 62860 18440 62894
rect 18616 62860 18628 62894
rect 18428 62848 18628 62860
rect 18428 62672 18628 62684
rect 18428 62638 18440 62672
rect 18616 62638 18628 62672
rect 18428 62626 18628 62638
rect 18428 62584 18628 62596
rect 18428 62550 18440 62584
rect 18616 62550 18628 62584
rect 18428 62538 18628 62550
rect 23418 62982 23618 62994
rect 23418 62948 23430 62982
rect 23606 62948 23618 62982
rect 23418 62936 23618 62948
rect 23418 62894 23618 62906
rect 23418 62860 23430 62894
rect 23606 62860 23618 62894
rect 23418 62848 23618 62860
rect 23418 62672 23618 62684
rect 23418 62638 23430 62672
rect 23606 62638 23618 62672
rect 23418 62626 23618 62638
rect 23418 62584 23618 62596
rect 23418 62550 23430 62584
rect 23606 62550 23618 62584
rect 23418 62538 23618 62550
rect 28408 62982 28608 62994
rect 28408 62948 28420 62982
rect 28596 62948 28608 62982
rect 28408 62936 28608 62948
rect 28408 62894 28608 62906
rect 28408 62860 28420 62894
rect 28596 62860 28608 62894
rect 28408 62848 28608 62860
rect 28408 62672 28608 62684
rect 28408 62638 28420 62672
rect 28596 62638 28608 62672
rect 28408 62626 28608 62638
rect 28408 62584 28608 62596
rect 28408 62550 28420 62584
rect 28596 62550 28608 62584
rect 28408 62538 28608 62550
rect 33398 62982 33598 62994
rect 33398 62948 33410 62982
rect 33586 62948 33598 62982
rect 33398 62936 33598 62948
rect 33398 62894 33598 62906
rect 33398 62860 33410 62894
rect 33586 62860 33598 62894
rect 33398 62848 33598 62860
rect 33398 62672 33598 62684
rect 33398 62638 33410 62672
rect 33586 62638 33598 62672
rect 33398 62626 33598 62638
rect 33398 62584 33598 62596
rect 33398 62550 33410 62584
rect 33586 62550 33598 62584
rect 33398 62538 33598 62550
rect 38388 62982 38588 62994
rect 38388 62948 38400 62982
rect 38576 62948 38588 62982
rect 38388 62936 38588 62948
rect 38388 62894 38588 62906
rect 38388 62860 38400 62894
rect 38576 62860 38588 62894
rect 38388 62848 38588 62860
rect 38388 62672 38588 62684
rect 38388 62638 38400 62672
rect 38576 62638 38588 62672
rect 38388 62626 38588 62638
rect 38388 62584 38588 62596
rect 38388 62550 38400 62584
rect 38576 62550 38588 62584
rect 38388 62538 38588 62550
rect 43378 62982 43578 62994
rect 43378 62948 43390 62982
rect 43566 62948 43578 62982
rect 43378 62936 43578 62948
rect 43378 62894 43578 62906
rect 43378 62860 43390 62894
rect 43566 62860 43578 62894
rect 43378 62848 43578 62860
rect 43378 62672 43578 62684
rect 43378 62638 43390 62672
rect 43566 62638 43578 62672
rect 43378 62626 43578 62638
rect 43378 62584 43578 62596
rect 43378 62550 43390 62584
rect 43566 62550 43578 62584
rect 43378 62538 43578 62550
rect 48368 62982 48568 62994
rect 48368 62948 48380 62982
rect 48556 62948 48568 62982
rect 48368 62936 48568 62948
rect 48368 62894 48568 62906
rect 48368 62860 48380 62894
rect 48556 62860 48568 62894
rect 48368 62848 48568 62860
rect 48368 62672 48568 62684
rect 48368 62638 48380 62672
rect 48556 62638 48568 62672
rect 48368 62626 48568 62638
rect 48368 62584 48568 62596
rect 48368 62550 48380 62584
rect 48556 62550 48568 62584
rect 48368 62538 48568 62550
rect 53358 62982 53558 62994
rect 53358 62948 53370 62982
rect 53546 62948 53558 62982
rect 53358 62936 53558 62948
rect 53358 62894 53558 62906
rect 53358 62860 53370 62894
rect 53546 62860 53558 62894
rect 53358 62848 53558 62860
rect 53358 62672 53558 62684
rect 53358 62638 53370 62672
rect 53546 62638 53558 62672
rect 53358 62626 53558 62638
rect 53358 62584 53558 62596
rect 53358 62550 53370 62584
rect 53546 62550 53558 62584
rect 53358 62538 53558 62550
rect 58348 62982 58548 62994
rect 58348 62948 58360 62982
rect 58536 62948 58548 62982
rect 58348 62936 58548 62948
rect 58348 62894 58548 62906
rect 58348 62860 58360 62894
rect 58536 62860 58548 62894
rect 58348 62848 58548 62860
rect 58348 62672 58548 62684
rect 58348 62638 58360 62672
rect 58536 62638 58548 62672
rect 58348 62626 58548 62638
rect 58348 62584 58548 62596
rect 58348 62550 58360 62584
rect 58536 62550 58548 62584
rect 58348 62538 58548 62550
rect 63338 62982 63538 62994
rect 63338 62948 63350 62982
rect 63526 62948 63538 62982
rect 63338 62936 63538 62948
rect 63338 62894 63538 62906
rect 63338 62860 63350 62894
rect 63526 62860 63538 62894
rect 63338 62848 63538 62860
rect 63338 62672 63538 62684
rect 63338 62638 63350 62672
rect 63526 62638 63538 62672
rect 63338 62626 63538 62638
rect 63338 62584 63538 62596
rect 63338 62550 63350 62584
rect 63526 62550 63538 62584
rect 63338 62538 63538 62550
rect 68328 62982 68528 62994
rect 68328 62948 68340 62982
rect 68516 62948 68528 62982
rect 68328 62936 68528 62948
rect 68328 62894 68528 62906
rect 68328 62860 68340 62894
rect 68516 62860 68528 62894
rect 68328 62848 68528 62860
rect 68328 62672 68528 62684
rect 68328 62638 68340 62672
rect 68516 62638 68528 62672
rect 68328 62626 68528 62638
rect 68328 62584 68528 62596
rect 68328 62550 68340 62584
rect 68516 62550 68528 62584
rect 68328 62538 68528 62550
rect 73318 62982 73518 62994
rect 73318 62948 73330 62982
rect 73506 62948 73518 62982
rect 73318 62936 73518 62948
rect 73318 62894 73518 62906
rect 73318 62860 73330 62894
rect 73506 62860 73518 62894
rect 73318 62848 73518 62860
rect 73318 62672 73518 62684
rect 73318 62638 73330 62672
rect 73506 62638 73518 62672
rect 73318 62626 73518 62638
rect 73318 62584 73518 62596
rect 73318 62550 73330 62584
rect 73506 62550 73518 62584
rect 73318 62538 73518 62550
rect 78308 62982 78508 62994
rect 78308 62948 78320 62982
rect 78496 62948 78508 62982
rect 78308 62936 78508 62948
rect 78308 62894 78508 62906
rect 78308 62860 78320 62894
rect 78496 62860 78508 62894
rect 78308 62848 78508 62860
rect 78308 62672 78508 62684
rect 78308 62638 78320 62672
rect 78496 62638 78508 62672
rect 78308 62626 78508 62638
rect 78308 62584 78508 62596
rect 78308 62550 78320 62584
rect 78496 62550 78508 62584
rect 78308 62538 78508 62550
rect 3458 61272 3658 61284
rect 3458 61238 3470 61272
rect 3646 61238 3658 61272
rect 3458 61226 3658 61238
rect 3458 61184 3658 61196
rect 3458 61150 3470 61184
rect 3646 61150 3658 61184
rect 3458 61138 3658 61150
rect 3458 60962 3658 60974
rect 3458 60928 3470 60962
rect 3646 60928 3658 60962
rect 3458 60916 3658 60928
rect 3458 60874 3658 60886
rect 3458 60840 3470 60874
rect 3646 60840 3658 60874
rect 3458 60828 3658 60840
rect 8448 61272 8648 61284
rect 8448 61238 8460 61272
rect 8636 61238 8648 61272
rect 8448 61226 8648 61238
rect 8448 61184 8648 61196
rect 8448 61150 8460 61184
rect 8636 61150 8648 61184
rect 8448 61138 8648 61150
rect 8448 60962 8648 60974
rect 8448 60928 8460 60962
rect 8636 60928 8648 60962
rect 8448 60916 8648 60928
rect 8448 60874 8648 60886
rect 8448 60840 8460 60874
rect 8636 60840 8648 60874
rect 8448 60828 8648 60840
rect 13438 61272 13638 61284
rect 13438 61238 13450 61272
rect 13626 61238 13638 61272
rect 13438 61226 13638 61238
rect 13438 61184 13638 61196
rect 13438 61150 13450 61184
rect 13626 61150 13638 61184
rect 13438 61138 13638 61150
rect 13438 60962 13638 60974
rect 13438 60928 13450 60962
rect 13626 60928 13638 60962
rect 13438 60916 13638 60928
rect 13438 60874 13638 60886
rect 13438 60840 13450 60874
rect 13626 60840 13638 60874
rect 13438 60828 13638 60840
rect 18428 61272 18628 61284
rect 18428 61238 18440 61272
rect 18616 61238 18628 61272
rect 18428 61226 18628 61238
rect 18428 61184 18628 61196
rect 18428 61150 18440 61184
rect 18616 61150 18628 61184
rect 18428 61138 18628 61150
rect 18428 60962 18628 60974
rect 18428 60928 18440 60962
rect 18616 60928 18628 60962
rect 18428 60916 18628 60928
rect 18428 60874 18628 60886
rect 18428 60840 18440 60874
rect 18616 60840 18628 60874
rect 18428 60828 18628 60840
rect 23418 61272 23618 61284
rect 23418 61238 23430 61272
rect 23606 61238 23618 61272
rect 23418 61226 23618 61238
rect 23418 61184 23618 61196
rect 23418 61150 23430 61184
rect 23606 61150 23618 61184
rect 23418 61138 23618 61150
rect 23418 60962 23618 60974
rect 23418 60928 23430 60962
rect 23606 60928 23618 60962
rect 23418 60916 23618 60928
rect 23418 60874 23618 60886
rect 23418 60840 23430 60874
rect 23606 60840 23618 60874
rect 23418 60828 23618 60840
rect 28408 61272 28608 61284
rect 28408 61238 28420 61272
rect 28596 61238 28608 61272
rect 28408 61226 28608 61238
rect 28408 61184 28608 61196
rect 28408 61150 28420 61184
rect 28596 61150 28608 61184
rect 28408 61138 28608 61150
rect 28408 60962 28608 60974
rect 28408 60928 28420 60962
rect 28596 60928 28608 60962
rect 28408 60916 28608 60928
rect 28408 60874 28608 60886
rect 28408 60840 28420 60874
rect 28596 60840 28608 60874
rect 28408 60828 28608 60840
rect 33398 61272 33598 61284
rect 33398 61238 33410 61272
rect 33586 61238 33598 61272
rect 33398 61226 33598 61238
rect 33398 61184 33598 61196
rect 33398 61150 33410 61184
rect 33586 61150 33598 61184
rect 33398 61138 33598 61150
rect 33398 60962 33598 60974
rect 33398 60928 33410 60962
rect 33586 60928 33598 60962
rect 33398 60916 33598 60928
rect 33398 60874 33598 60886
rect 33398 60840 33410 60874
rect 33586 60840 33598 60874
rect 33398 60828 33598 60840
rect 38388 61272 38588 61284
rect 38388 61238 38400 61272
rect 38576 61238 38588 61272
rect 38388 61226 38588 61238
rect 38388 61184 38588 61196
rect 38388 61150 38400 61184
rect 38576 61150 38588 61184
rect 38388 61138 38588 61150
rect 38388 60962 38588 60974
rect 38388 60928 38400 60962
rect 38576 60928 38588 60962
rect 38388 60916 38588 60928
rect 38388 60874 38588 60886
rect 38388 60840 38400 60874
rect 38576 60840 38588 60874
rect 38388 60828 38588 60840
rect 43378 61272 43578 61284
rect 43378 61238 43390 61272
rect 43566 61238 43578 61272
rect 43378 61226 43578 61238
rect 43378 61184 43578 61196
rect 43378 61150 43390 61184
rect 43566 61150 43578 61184
rect 43378 61138 43578 61150
rect 43378 60962 43578 60974
rect 43378 60928 43390 60962
rect 43566 60928 43578 60962
rect 43378 60916 43578 60928
rect 43378 60874 43578 60886
rect 43378 60840 43390 60874
rect 43566 60840 43578 60874
rect 43378 60828 43578 60840
rect 48368 61272 48568 61284
rect 48368 61238 48380 61272
rect 48556 61238 48568 61272
rect 48368 61226 48568 61238
rect 48368 61184 48568 61196
rect 48368 61150 48380 61184
rect 48556 61150 48568 61184
rect 48368 61138 48568 61150
rect 48368 60962 48568 60974
rect 48368 60928 48380 60962
rect 48556 60928 48568 60962
rect 48368 60916 48568 60928
rect 48368 60874 48568 60886
rect 48368 60840 48380 60874
rect 48556 60840 48568 60874
rect 48368 60828 48568 60840
rect 53358 61272 53558 61284
rect 53358 61238 53370 61272
rect 53546 61238 53558 61272
rect 53358 61226 53558 61238
rect 53358 61184 53558 61196
rect 53358 61150 53370 61184
rect 53546 61150 53558 61184
rect 53358 61138 53558 61150
rect 53358 60962 53558 60974
rect 53358 60928 53370 60962
rect 53546 60928 53558 60962
rect 53358 60916 53558 60928
rect 53358 60874 53558 60886
rect 53358 60840 53370 60874
rect 53546 60840 53558 60874
rect 53358 60828 53558 60840
rect 58348 61272 58548 61284
rect 58348 61238 58360 61272
rect 58536 61238 58548 61272
rect 58348 61226 58548 61238
rect 58348 61184 58548 61196
rect 58348 61150 58360 61184
rect 58536 61150 58548 61184
rect 58348 61138 58548 61150
rect 58348 60962 58548 60974
rect 58348 60928 58360 60962
rect 58536 60928 58548 60962
rect 58348 60916 58548 60928
rect 58348 60874 58548 60886
rect 58348 60840 58360 60874
rect 58536 60840 58548 60874
rect 58348 60828 58548 60840
rect 63338 61272 63538 61284
rect 63338 61238 63350 61272
rect 63526 61238 63538 61272
rect 63338 61226 63538 61238
rect 63338 61184 63538 61196
rect 63338 61150 63350 61184
rect 63526 61150 63538 61184
rect 63338 61138 63538 61150
rect 63338 60962 63538 60974
rect 63338 60928 63350 60962
rect 63526 60928 63538 60962
rect 63338 60916 63538 60928
rect 63338 60874 63538 60886
rect 63338 60840 63350 60874
rect 63526 60840 63538 60874
rect 63338 60828 63538 60840
rect 68328 61272 68528 61284
rect 68328 61238 68340 61272
rect 68516 61238 68528 61272
rect 68328 61226 68528 61238
rect 68328 61184 68528 61196
rect 68328 61150 68340 61184
rect 68516 61150 68528 61184
rect 68328 61138 68528 61150
rect 68328 60962 68528 60974
rect 68328 60928 68340 60962
rect 68516 60928 68528 60962
rect 68328 60916 68528 60928
rect 68328 60874 68528 60886
rect 68328 60840 68340 60874
rect 68516 60840 68528 60874
rect 68328 60828 68528 60840
rect 73318 61272 73518 61284
rect 73318 61238 73330 61272
rect 73506 61238 73518 61272
rect 73318 61226 73518 61238
rect 73318 61184 73518 61196
rect 73318 61150 73330 61184
rect 73506 61150 73518 61184
rect 73318 61138 73518 61150
rect 73318 60962 73518 60974
rect 73318 60928 73330 60962
rect 73506 60928 73518 60962
rect 73318 60916 73518 60928
rect 73318 60874 73518 60886
rect 73318 60840 73330 60874
rect 73506 60840 73518 60874
rect 73318 60828 73518 60840
rect 78308 61272 78508 61284
rect 78308 61238 78320 61272
rect 78496 61238 78508 61272
rect 78308 61226 78508 61238
rect 78308 61184 78508 61196
rect 78308 61150 78320 61184
rect 78496 61150 78508 61184
rect 78308 61138 78508 61150
rect 78308 60962 78508 60974
rect 78308 60928 78320 60962
rect 78496 60928 78508 60962
rect 78308 60916 78508 60928
rect 78308 60874 78508 60886
rect 78308 60840 78320 60874
rect 78496 60840 78508 60874
rect 78308 60828 78508 60840
rect 3458 59562 3658 59574
rect 3458 59528 3470 59562
rect 3646 59528 3658 59562
rect 3458 59516 3658 59528
rect 3458 59474 3658 59486
rect 3458 59440 3470 59474
rect 3646 59440 3658 59474
rect 3458 59428 3658 59440
rect 3458 59252 3658 59264
rect 3458 59218 3470 59252
rect 3646 59218 3658 59252
rect 3458 59206 3658 59218
rect 3458 59164 3658 59176
rect 3458 59130 3470 59164
rect 3646 59130 3658 59164
rect 3458 59118 3658 59130
rect 8448 59562 8648 59574
rect 8448 59528 8460 59562
rect 8636 59528 8648 59562
rect 8448 59516 8648 59528
rect 8448 59474 8648 59486
rect 8448 59440 8460 59474
rect 8636 59440 8648 59474
rect 8448 59428 8648 59440
rect 8448 59252 8648 59264
rect 8448 59218 8460 59252
rect 8636 59218 8648 59252
rect 8448 59206 8648 59218
rect 8448 59164 8648 59176
rect 8448 59130 8460 59164
rect 8636 59130 8648 59164
rect 8448 59118 8648 59130
rect 13438 59562 13638 59574
rect 13438 59528 13450 59562
rect 13626 59528 13638 59562
rect 13438 59516 13638 59528
rect 13438 59474 13638 59486
rect 13438 59440 13450 59474
rect 13626 59440 13638 59474
rect 13438 59428 13638 59440
rect 13438 59252 13638 59264
rect 13438 59218 13450 59252
rect 13626 59218 13638 59252
rect 13438 59206 13638 59218
rect 13438 59164 13638 59176
rect 13438 59130 13450 59164
rect 13626 59130 13638 59164
rect 13438 59118 13638 59130
rect 18428 59562 18628 59574
rect 18428 59528 18440 59562
rect 18616 59528 18628 59562
rect 18428 59516 18628 59528
rect 18428 59474 18628 59486
rect 18428 59440 18440 59474
rect 18616 59440 18628 59474
rect 18428 59428 18628 59440
rect 18428 59252 18628 59264
rect 18428 59218 18440 59252
rect 18616 59218 18628 59252
rect 18428 59206 18628 59218
rect 18428 59164 18628 59176
rect 18428 59130 18440 59164
rect 18616 59130 18628 59164
rect 18428 59118 18628 59130
rect 23418 59562 23618 59574
rect 23418 59528 23430 59562
rect 23606 59528 23618 59562
rect 23418 59516 23618 59528
rect 23418 59474 23618 59486
rect 23418 59440 23430 59474
rect 23606 59440 23618 59474
rect 23418 59428 23618 59440
rect 23418 59252 23618 59264
rect 23418 59218 23430 59252
rect 23606 59218 23618 59252
rect 23418 59206 23618 59218
rect 23418 59164 23618 59176
rect 23418 59130 23430 59164
rect 23606 59130 23618 59164
rect 23418 59118 23618 59130
rect 28408 59562 28608 59574
rect 28408 59528 28420 59562
rect 28596 59528 28608 59562
rect 28408 59516 28608 59528
rect 28408 59474 28608 59486
rect 28408 59440 28420 59474
rect 28596 59440 28608 59474
rect 28408 59428 28608 59440
rect 28408 59252 28608 59264
rect 28408 59218 28420 59252
rect 28596 59218 28608 59252
rect 28408 59206 28608 59218
rect 28408 59164 28608 59176
rect 28408 59130 28420 59164
rect 28596 59130 28608 59164
rect 28408 59118 28608 59130
rect 33398 59562 33598 59574
rect 33398 59528 33410 59562
rect 33586 59528 33598 59562
rect 33398 59516 33598 59528
rect 33398 59474 33598 59486
rect 33398 59440 33410 59474
rect 33586 59440 33598 59474
rect 33398 59428 33598 59440
rect 33398 59252 33598 59264
rect 33398 59218 33410 59252
rect 33586 59218 33598 59252
rect 33398 59206 33598 59218
rect 33398 59164 33598 59176
rect 33398 59130 33410 59164
rect 33586 59130 33598 59164
rect 33398 59118 33598 59130
rect 38388 59562 38588 59574
rect 38388 59528 38400 59562
rect 38576 59528 38588 59562
rect 38388 59516 38588 59528
rect 38388 59474 38588 59486
rect 38388 59440 38400 59474
rect 38576 59440 38588 59474
rect 38388 59428 38588 59440
rect 38388 59252 38588 59264
rect 38388 59218 38400 59252
rect 38576 59218 38588 59252
rect 38388 59206 38588 59218
rect 38388 59164 38588 59176
rect 38388 59130 38400 59164
rect 38576 59130 38588 59164
rect 38388 59118 38588 59130
rect 43378 59562 43578 59574
rect 43378 59528 43390 59562
rect 43566 59528 43578 59562
rect 43378 59516 43578 59528
rect 43378 59474 43578 59486
rect 43378 59440 43390 59474
rect 43566 59440 43578 59474
rect 43378 59428 43578 59440
rect 43378 59252 43578 59264
rect 43378 59218 43390 59252
rect 43566 59218 43578 59252
rect 43378 59206 43578 59218
rect 43378 59164 43578 59176
rect 43378 59130 43390 59164
rect 43566 59130 43578 59164
rect 43378 59118 43578 59130
rect 48368 59562 48568 59574
rect 48368 59528 48380 59562
rect 48556 59528 48568 59562
rect 48368 59516 48568 59528
rect 48368 59474 48568 59486
rect 48368 59440 48380 59474
rect 48556 59440 48568 59474
rect 48368 59428 48568 59440
rect 48368 59252 48568 59264
rect 48368 59218 48380 59252
rect 48556 59218 48568 59252
rect 48368 59206 48568 59218
rect 48368 59164 48568 59176
rect 48368 59130 48380 59164
rect 48556 59130 48568 59164
rect 48368 59118 48568 59130
rect 53358 59562 53558 59574
rect 53358 59528 53370 59562
rect 53546 59528 53558 59562
rect 53358 59516 53558 59528
rect 53358 59474 53558 59486
rect 53358 59440 53370 59474
rect 53546 59440 53558 59474
rect 53358 59428 53558 59440
rect 53358 59252 53558 59264
rect 53358 59218 53370 59252
rect 53546 59218 53558 59252
rect 53358 59206 53558 59218
rect 53358 59164 53558 59176
rect 53358 59130 53370 59164
rect 53546 59130 53558 59164
rect 53358 59118 53558 59130
rect 58348 59562 58548 59574
rect 58348 59528 58360 59562
rect 58536 59528 58548 59562
rect 58348 59516 58548 59528
rect 58348 59474 58548 59486
rect 58348 59440 58360 59474
rect 58536 59440 58548 59474
rect 58348 59428 58548 59440
rect 58348 59252 58548 59264
rect 58348 59218 58360 59252
rect 58536 59218 58548 59252
rect 58348 59206 58548 59218
rect 58348 59164 58548 59176
rect 58348 59130 58360 59164
rect 58536 59130 58548 59164
rect 58348 59118 58548 59130
rect 63338 59562 63538 59574
rect 63338 59528 63350 59562
rect 63526 59528 63538 59562
rect 63338 59516 63538 59528
rect 63338 59474 63538 59486
rect 63338 59440 63350 59474
rect 63526 59440 63538 59474
rect 63338 59428 63538 59440
rect 63338 59252 63538 59264
rect 63338 59218 63350 59252
rect 63526 59218 63538 59252
rect 63338 59206 63538 59218
rect 63338 59164 63538 59176
rect 63338 59130 63350 59164
rect 63526 59130 63538 59164
rect 63338 59118 63538 59130
rect 68328 59562 68528 59574
rect 68328 59528 68340 59562
rect 68516 59528 68528 59562
rect 68328 59516 68528 59528
rect 68328 59474 68528 59486
rect 68328 59440 68340 59474
rect 68516 59440 68528 59474
rect 68328 59428 68528 59440
rect 68328 59252 68528 59264
rect 68328 59218 68340 59252
rect 68516 59218 68528 59252
rect 68328 59206 68528 59218
rect 68328 59164 68528 59176
rect 68328 59130 68340 59164
rect 68516 59130 68528 59164
rect 68328 59118 68528 59130
rect 73318 59562 73518 59574
rect 73318 59528 73330 59562
rect 73506 59528 73518 59562
rect 73318 59516 73518 59528
rect 73318 59474 73518 59486
rect 73318 59440 73330 59474
rect 73506 59440 73518 59474
rect 73318 59428 73518 59440
rect 73318 59252 73518 59264
rect 73318 59218 73330 59252
rect 73506 59218 73518 59252
rect 73318 59206 73518 59218
rect 73318 59164 73518 59176
rect 73318 59130 73330 59164
rect 73506 59130 73518 59164
rect 73318 59118 73518 59130
rect 78308 59562 78508 59574
rect 78308 59528 78320 59562
rect 78496 59528 78508 59562
rect 78308 59516 78508 59528
rect 78308 59474 78508 59486
rect 78308 59440 78320 59474
rect 78496 59440 78508 59474
rect 78308 59428 78508 59440
rect 78308 59252 78508 59264
rect 78308 59218 78320 59252
rect 78496 59218 78508 59252
rect 78308 59206 78508 59218
rect 78308 59164 78508 59176
rect 78308 59130 78320 59164
rect 78496 59130 78508 59164
rect 78308 59118 78508 59130
rect 3458 57852 3658 57864
rect 3458 57818 3470 57852
rect 3646 57818 3658 57852
rect 3458 57806 3658 57818
rect 3458 57764 3658 57776
rect 3458 57730 3470 57764
rect 3646 57730 3658 57764
rect 3458 57718 3658 57730
rect 3458 57542 3658 57554
rect 3458 57508 3470 57542
rect 3646 57508 3658 57542
rect 3458 57496 3658 57508
rect 3458 57454 3658 57466
rect 3458 57420 3470 57454
rect 3646 57420 3658 57454
rect 3458 57408 3658 57420
rect 8448 57852 8648 57864
rect 8448 57818 8460 57852
rect 8636 57818 8648 57852
rect 8448 57806 8648 57818
rect 8448 57764 8648 57776
rect 8448 57730 8460 57764
rect 8636 57730 8648 57764
rect 8448 57718 8648 57730
rect 8448 57542 8648 57554
rect 8448 57508 8460 57542
rect 8636 57508 8648 57542
rect 8448 57496 8648 57508
rect 8448 57454 8648 57466
rect 8448 57420 8460 57454
rect 8636 57420 8648 57454
rect 8448 57408 8648 57420
rect 13438 57852 13638 57864
rect 13438 57818 13450 57852
rect 13626 57818 13638 57852
rect 13438 57806 13638 57818
rect 13438 57764 13638 57776
rect 13438 57730 13450 57764
rect 13626 57730 13638 57764
rect 13438 57718 13638 57730
rect 13438 57542 13638 57554
rect 13438 57508 13450 57542
rect 13626 57508 13638 57542
rect 13438 57496 13638 57508
rect 13438 57454 13638 57466
rect 13438 57420 13450 57454
rect 13626 57420 13638 57454
rect 13438 57408 13638 57420
rect 18428 57852 18628 57864
rect 18428 57818 18440 57852
rect 18616 57818 18628 57852
rect 18428 57806 18628 57818
rect 18428 57764 18628 57776
rect 18428 57730 18440 57764
rect 18616 57730 18628 57764
rect 18428 57718 18628 57730
rect 18428 57542 18628 57554
rect 18428 57508 18440 57542
rect 18616 57508 18628 57542
rect 18428 57496 18628 57508
rect 18428 57454 18628 57466
rect 18428 57420 18440 57454
rect 18616 57420 18628 57454
rect 18428 57408 18628 57420
rect 23418 57852 23618 57864
rect 23418 57818 23430 57852
rect 23606 57818 23618 57852
rect 23418 57806 23618 57818
rect 23418 57764 23618 57776
rect 23418 57730 23430 57764
rect 23606 57730 23618 57764
rect 23418 57718 23618 57730
rect 23418 57542 23618 57554
rect 23418 57508 23430 57542
rect 23606 57508 23618 57542
rect 23418 57496 23618 57508
rect 23418 57454 23618 57466
rect 23418 57420 23430 57454
rect 23606 57420 23618 57454
rect 23418 57408 23618 57420
rect 28408 57852 28608 57864
rect 28408 57818 28420 57852
rect 28596 57818 28608 57852
rect 28408 57806 28608 57818
rect 28408 57764 28608 57776
rect 28408 57730 28420 57764
rect 28596 57730 28608 57764
rect 28408 57718 28608 57730
rect 28408 57542 28608 57554
rect 28408 57508 28420 57542
rect 28596 57508 28608 57542
rect 28408 57496 28608 57508
rect 28408 57454 28608 57466
rect 28408 57420 28420 57454
rect 28596 57420 28608 57454
rect 28408 57408 28608 57420
rect 33398 57852 33598 57864
rect 33398 57818 33410 57852
rect 33586 57818 33598 57852
rect 33398 57806 33598 57818
rect 33398 57764 33598 57776
rect 33398 57730 33410 57764
rect 33586 57730 33598 57764
rect 33398 57718 33598 57730
rect 33398 57542 33598 57554
rect 33398 57508 33410 57542
rect 33586 57508 33598 57542
rect 33398 57496 33598 57508
rect 33398 57454 33598 57466
rect 33398 57420 33410 57454
rect 33586 57420 33598 57454
rect 33398 57408 33598 57420
rect 38388 57852 38588 57864
rect 38388 57818 38400 57852
rect 38576 57818 38588 57852
rect 38388 57806 38588 57818
rect 38388 57764 38588 57776
rect 38388 57730 38400 57764
rect 38576 57730 38588 57764
rect 38388 57718 38588 57730
rect 38388 57542 38588 57554
rect 38388 57508 38400 57542
rect 38576 57508 38588 57542
rect 38388 57496 38588 57508
rect 38388 57454 38588 57466
rect 38388 57420 38400 57454
rect 38576 57420 38588 57454
rect 38388 57408 38588 57420
rect 43378 57852 43578 57864
rect 43378 57818 43390 57852
rect 43566 57818 43578 57852
rect 43378 57806 43578 57818
rect 43378 57764 43578 57776
rect 43378 57730 43390 57764
rect 43566 57730 43578 57764
rect 43378 57718 43578 57730
rect 43378 57542 43578 57554
rect 43378 57508 43390 57542
rect 43566 57508 43578 57542
rect 43378 57496 43578 57508
rect 43378 57454 43578 57466
rect 43378 57420 43390 57454
rect 43566 57420 43578 57454
rect 43378 57408 43578 57420
rect 48368 57852 48568 57864
rect 48368 57818 48380 57852
rect 48556 57818 48568 57852
rect 48368 57806 48568 57818
rect 48368 57764 48568 57776
rect 48368 57730 48380 57764
rect 48556 57730 48568 57764
rect 48368 57718 48568 57730
rect 48368 57542 48568 57554
rect 48368 57508 48380 57542
rect 48556 57508 48568 57542
rect 48368 57496 48568 57508
rect 48368 57454 48568 57466
rect 48368 57420 48380 57454
rect 48556 57420 48568 57454
rect 48368 57408 48568 57420
rect 53358 57852 53558 57864
rect 53358 57818 53370 57852
rect 53546 57818 53558 57852
rect 53358 57806 53558 57818
rect 53358 57764 53558 57776
rect 53358 57730 53370 57764
rect 53546 57730 53558 57764
rect 53358 57718 53558 57730
rect 53358 57542 53558 57554
rect 53358 57508 53370 57542
rect 53546 57508 53558 57542
rect 53358 57496 53558 57508
rect 53358 57454 53558 57466
rect 53358 57420 53370 57454
rect 53546 57420 53558 57454
rect 53358 57408 53558 57420
rect 58348 57852 58548 57864
rect 58348 57818 58360 57852
rect 58536 57818 58548 57852
rect 58348 57806 58548 57818
rect 58348 57764 58548 57776
rect 58348 57730 58360 57764
rect 58536 57730 58548 57764
rect 58348 57718 58548 57730
rect 58348 57542 58548 57554
rect 58348 57508 58360 57542
rect 58536 57508 58548 57542
rect 58348 57496 58548 57508
rect 58348 57454 58548 57466
rect 58348 57420 58360 57454
rect 58536 57420 58548 57454
rect 58348 57408 58548 57420
rect 63338 57852 63538 57864
rect 63338 57818 63350 57852
rect 63526 57818 63538 57852
rect 63338 57806 63538 57818
rect 63338 57764 63538 57776
rect 63338 57730 63350 57764
rect 63526 57730 63538 57764
rect 63338 57718 63538 57730
rect 63338 57542 63538 57554
rect 63338 57508 63350 57542
rect 63526 57508 63538 57542
rect 63338 57496 63538 57508
rect 63338 57454 63538 57466
rect 63338 57420 63350 57454
rect 63526 57420 63538 57454
rect 63338 57408 63538 57420
rect 68328 57852 68528 57864
rect 68328 57818 68340 57852
rect 68516 57818 68528 57852
rect 68328 57806 68528 57818
rect 68328 57764 68528 57776
rect 68328 57730 68340 57764
rect 68516 57730 68528 57764
rect 68328 57718 68528 57730
rect 68328 57542 68528 57554
rect 68328 57508 68340 57542
rect 68516 57508 68528 57542
rect 68328 57496 68528 57508
rect 68328 57454 68528 57466
rect 68328 57420 68340 57454
rect 68516 57420 68528 57454
rect 68328 57408 68528 57420
rect 73318 57852 73518 57864
rect 73318 57818 73330 57852
rect 73506 57818 73518 57852
rect 73318 57806 73518 57818
rect 73318 57764 73518 57776
rect 73318 57730 73330 57764
rect 73506 57730 73518 57764
rect 73318 57718 73518 57730
rect 73318 57542 73518 57554
rect 73318 57508 73330 57542
rect 73506 57508 73518 57542
rect 73318 57496 73518 57508
rect 73318 57454 73518 57466
rect 73318 57420 73330 57454
rect 73506 57420 73518 57454
rect 73318 57408 73518 57420
rect 78308 57852 78508 57864
rect 78308 57818 78320 57852
rect 78496 57818 78508 57852
rect 78308 57806 78508 57818
rect 78308 57764 78508 57776
rect 78308 57730 78320 57764
rect 78496 57730 78508 57764
rect 78308 57718 78508 57730
rect 78308 57542 78508 57554
rect 78308 57508 78320 57542
rect 78496 57508 78508 57542
rect 78308 57496 78508 57508
rect 78308 57454 78508 57466
rect 78308 57420 78320 57454
rect 78496 57420 78508 57454
rect 78308 57408 78508 57420
rect 3458 56142 3658 56154
rect 3458 56108 3470 56142
rect 3646 56108 3658 56142
rect 3458 56096 3658 56108
rect 3458 56054 3658 56066
rect 3458 56020 3470 56054
rect 3646 56020 3658 56054
rect 3458 56008 3658 56020
rect 3458 55832 3658 55844
rect 3458 55798 3470 55832
rect 3646 55798 3658 55832
rect 3458 55786 3658 55798
rect 3458 55744 3658 55756
rect 3458 55710 3470 55744
rect 3646 55710 3658 55744
rect 3458 55698 3658 55710
rect 8448 56142 8648 56154
rect 8448 56108 8460 56142
rect 8636 56108 8648 56142
rect 8448 56096 8648 56108
rect 8448 56054 8648 56066
rect 8448 56020 8460 56054
rect 8636 56020 8648 56054
rect 8448 56008 8648 56020
rect 8448 55832 8648 55844
rect 8448 55798 8460 55832
rect 8636 55798 8648 55832
rect 8448 55786 8648 55798
rect 8448 55744 8648 55756
rect 8448 55710 8460 55744
rect 8636 55710 8648 55744
rect 8448 55698 8648 55710
rect 13438 56142 13638 56154
rect 13438 56108 13450 56142
rect 13626 56108 13638 56142
rect 13438 56096 13638 56108
rect 13438 56054 13638 56066
rect 13438 56020 13450 56054
rect 13626 56020 13638 56054
rect 13438 56008 13638 56020
rect 13438 55832 13638 55844
rect 13438 55798 13450 55832
rect 13626 55798 13638 55832
rect 13438 55786 13638 55798
rect 13438 55744 13638 55756
rect 13438 55710 13450 55744
rect 13626 55710 13638 55744
rect 13438 55698 13638 55710
rect 18428 56142 18628 56154
rect 18428 56108 18440 56142
rect 18616 56108 18628 56142
rect 18428 56096 18628 56108
rect 18428 56054 18628 56066
rect 18428 56020 18440 56054
rect 18616 56020 18628 56054
rect 18428 56008 18628 56020
rect 18428 55832 18628 55844
rect 18428 55798 18440 55832
rect 18616 55798 18628 55832
rect 18428 55786 18628 55798
rect 18428 55744 18628 55756
rect 18428 55710 18440 55744
rect 18616 55710 18628 55744
rect 18428 55698 18628 55710
rect 23418 56142 23618 56154
rect 23418 56108 23430 56142
rect 23606 56108 23618 56142
rect 23418 56096 23618 56108
rect 23418 56054 23618 56066
rect 23418 56020 23430 56054
rect 23606 56020 23618 56054
rect 23418 56008 23618 56020
rect 23418 55832 23618 55844
rect 23418 55798 23430 55832
rect 23606 55798 23618 55832
rect 23418 55786 23618 55798
rect 23418 55744 23618 55756
rect 23418 55710 23430 55744
rect 23606 55710 23618 55744
rect 23418 55698 23618 55710
rect 28408 56142 28608 56154
rect 28408 56108 28420 56142
rect 28596 56108 28608 56142
rect 28408 56096 28608 56108
rect 28408 56054 28608 56066
rect 28408 56020 28420 56054
rect 28596 56020 28608 56054
rect 28408 56008 28608 56020
rect 28408 55832 28608 55844
rect 28408 55798 28420 55832
rect 28596 55798 28608 55832
rect 28408 55786 28608 55798
rect 28408 55744 28608 55756
rect 28408 55710 28420 55744
rect 28596 55710 28608 55744
rect 28408 55698 28608 55710
rect 33398 56142 33598 56154
rect 33398 56108 33410 56142
rect 33586 56108 33598 56142
rect 33398 56096 33598 56108
rect 33398 56054 33598 56066
rect 33398 56020 33410 56054
rect 33586 56020 33598 56054
rect 33398 56008 33598 56020
rect 33398 55832 33598 55844
rect 33398 55798 33410 55832
rect 33586 55798 33598 55832
rect 33398 55786 33598 55798
rect 33398 55744 33598 55756
rect 33398 55710 33410 55744
rect 33586 55710 33598 55744
rect 33398 55698 33598 55710
rect 38388 56142 38588 56154
rect 38388 56108 38400 56142
rect 38576 56108 38588 56142
rect 38388 56096 38588 56108
rect 38388 56054 38588 56066
rect 38388 56020 38400 56054
rect 38576 56020 38588 56054
rect 38388 56008 38588 56020
rect 38388 55832 38588 55844
rect 38388 55798 38400 55832
rect 38576 55798 38588 55832
rect 38388 55786 38588 55798
rect 38388 55744 38588 55756
rect 38388 55710 38400 55744
rect 38576 55710 38588 55744
rect 38388 55698 38588 55710
rect 43378 56142 43578 56154
rect 43378 56108 43390 56142
rect 43566 56108 43578 56142
rect 43378 56096 43578 56108
rect 43378 56054 43578 56066
rect 43378 56020 43390 56054
rect 43566 56020 43578 56054
rect 43378 56008 43578 56020
rect 43378 55832 43578 55844
rect 43378 55798 43390 55832
rect 43566 55798 43578 55832
rect 43378 55786 43578 55798
rect 43378 55744 43578 55756
rect 43378 55710 43390 55744
rect 43566 55710 43578 55744
rect 43378 55698 43578 55710
rect 48368 56142 48568 56154
rect 48368 56108 48380 56142
rect 48556 56108 48568 56142
rect 48368 56096 48568 56108
rect 48368 56054 48568 56066
rect 48368 56020 48380 56054
rect 48556 56020 48568 56054
rect 48368 56008 48568 56020
rect 48368 55832 48568 55844
rect 48368 55798 48380 55832
rect 48556 55798 48568 55832
rect 48368 55786 48568 55798
rect 48368 55744 48568 55756
rect 48368 55710 48380 55744
rect 48556 55710 48568 55744
rect 48368 55698 48568 55710
rect 53358 56142 53558 56154
rect 53358 56108 53370 56142
rect 53546 56108 53558 56142
rect 53358 56096 53558 56108
rect 53358 56054 53558 56066
rect 53358 56020 53370 56054
rect 53546 56020 53558 56054
rect 53358 56008 53558 56020
rect 53358 55832 53558 55844
rect 53358 55798 53370 55832
rect 53546 55798 53558 55832
rect 53358 55786 53558 55798
rect 53358 55744 53558 55756
rect 53358 55710 53370 55744
rect 53546 55710 53558 55744
rect 53358 55698 53558 55710
rect 58348 56142 58548 56154
rect 58348 56108 58360 56142
rect 58536 56108 58548 56142
rect 58348 56096 58548 56108
rect 58348 56054 58548 56066
rect 58348 56020 58360 56054
rect 58536 56020 58548 56054
rect 58348 56008 58548 56020
rect 58348 55832 58548 55844
rect 58348 55798 58360 55832
rect 58536 55798 58548 55832
rect 58348 55786 58548 55798
rect 58348 55744 58548 55756
rect 58348 55710 58360 55744
rect 58536 55710 58548 55744
rect 58348 55698 58548 55710
rect 63338 56142 63538 56154
rect 63338 56108 63350 56142
rect 63526 56108 63538 56142
rect 63338 56096 63538 56108
rect 63338 56054 63538 56066
rect 63338 56020 63350 56054
rect 63526 56020 63538 56054
rect 63338 56008 63538 56020
rect 63338 55832 63538 55844
rect 63338 55798 63350 55832
rect 63526 55798 63538 55832
rect 63338 55786 63538 55798
rect 63338 55744 63538 55756
rect 63338 55710 63350 55744
rect 63526 55710 63538 55744
rect 63338 55698 63538 55710
rect 68328 56142 68528 56154
rect 68328 56108 68340 56142
rect 68516 56108 68528 56142
rect 68328 56096 68528 56108
rect 68328 56054 68528 56066
rect 68328 56020 68340 56054
rect 68516 56020 68528 56054
rect 68328 56008 68528 56020
rect 68328 55832 68528 55844
rect 68328 55798 68340 55832
rect 68516 55798 68528 55832
rect 68328 55786 68528 55798
rect 68328 55744 68528 55756
rect 68328 55710 68340 55744
rect 68516 55710 68528 55744
rect 68328 55698 68528 55710
rect 73318 56142 73518 56154
rect 73318 56108 73330 56142
rect 73506 56108 73518 56142
rect 73318 56096 73518 56108
rect 73318 56054 73518 56066
rect 73318 56020 73330 56054
rect 73506 56020 73518 56054
rect 73318 56008 73518 56020
rect 73318 55832 73518 55844
rect 73318 55798 73330 55832
rect 73506 55798 73518 55832
rect 73318 55786 73518 55798
rect 73318 55744 73518 55756
rect 73318 55710 73330 55744
rect 73506 55710 73518 55744
rect 73318 55698 73518 55710
rect 78308 56142 78508 56154
rect 78308 56108 78320 56142
rect 78496 56108 78508 56142
rect 78308 56096 78508 56108
rect 78308 56054 78508 56066
rect 78308 56020 78320 56054
rect 78496 56020 78508 56054
rect 78308 56008 78508 56020
rect 78308 55832 78508 55844
rect 78308 55798 78320 55832
rect 78496 55798 78508 55832
rect 78308 55786 78508 55798
rect 78308 55744 78508 55756
rect 78308 55710 78320 55744
rect 78496 55710 78508 55744
rect 78308 55698 78508 55710
rect 3458 54432 3658 54444
rect 3458 54398 3470 54432
rect 3646 54398 3658 54432
rect 3458 54386 3658 54398
rect 3458 54344 3658 54356
rect 3458 54310 3470 54344
rect 3646 54310 3658 54344
rect 3458 54298 3658 54310
rect 3458 54122 3658 54134
rect 3458 54088 3470 54122
rect 3646 54088 3658 54122
rect 3458 54076 3658 54088
rect 3458 54034 3658 54046
rect 3458 54000 3470 54034
rect 3646 54000 3658 54034
rect 3458 53988 3658 54000
rect 8448 54432 8648 54444
rect 8448 54398 8460 54432
rect 8636 54398 8648 54432
rect 8448 54386 8648 54398
rect 8448 54344 8648 54356
rect 8448 54310 8460 54344
rect 8636 54310 8648 54344
rect 8448 54298 8648 54310
rect 8448 54122 8648 54134
rect 8448 54088 8460 54122
rect 8636 54088 8648 54122
rect 8448 54076 8648 54088
rect 8448 54034 8648 54046
rect 8448 54000 8460 54034
rect 8636 54000 8648 54034
rect 8448 53988 8648 54000
rect 13438 54432 13638 54444
rect 13438 54398 13450 54432
rect 13626 54398 13638 54432
rect 13438 54386 13638 54398
rect 13438 54344 13638 54356
rect 13438 54310 13450 54344
rect 13626 54310 13638 54344
rect 13438 54298 13638 54310
rect 13438 54122 13638 54134
rect 13438 54088 13450 54122
rect 13626 54088 13638 54122
rect 13438 54076 13638 54088
rect 13438 54034 13638 54046
rect 13438 54000 13450 54034
rect 13626 54000 13638 54034
rect 13438 53988 13638 54000
rect 18428 54432 18628 54444
rect 18428 54398 18440 54432
rect 18616 54398 18628 54432
rect 18428 54386 18628 54398
rect 18428 54344 18628 54356
rect 18428 54310 18440 54344
rect 18616 54310 18628 54344
rect 18428 54298 18628 54310
rect 18428 54122 18628 54134
rect 18428 54088 18440 54122
rect 18616 54088 18628 54122
rect 18428 54076 18628 54088
rect 18428 54034 18628 54046
rect 18428 54000 18440 54034
rect 18616 54000 18628 54034
rect 18428 53988 18628 54000
rect 23418 54432 23618 54444
rect 23418 54398 23430 54432
rect 23606 54398 23618 54432
rect 23418 54386 23618 54398
rect 23418 54344 23618 54356
rect 23418 54310 23430 54344
rect 23606 54310 23618 54344
rect 23418 54298 23618 54310
rect 23418 54122 23618 54134
rect 23418 54088 23430 54122
rect 23606 54088 23618 54122
rect 23418 54076 23618 54088
rect 23418 54034 23618 54046
rect 23418 54000 23430 54034
rect 23606 54000 23618 54034
rect 23418 53988 23618 54000
rect 28408 54432 28608 54444
rect 28408 54398 28420 54432
rect 28596 54398 28608 54432
rect 28408 54386 28608 54398
rect 28408 54344 28608 54356
rect 28408 54310 28420 54344
rect 28596 54310 28608 54344
rect 28408 54298 28608 54310
rect 28408 54122 28608 54134
rect 28408 54088 28420 54122
rect 28596 54088 28608 54122
rect 28408 54076 28608 54088
rect 28408 54034 28608 54046
rect 28408 54000 28420 54034
rect 28596 54000 28608 54034
rect 28408 53988 28608 54000
rect 33398 54432 33598 54444
rect 33398 54398 33410 54432
rect 33586 54398 33598 54432
rect 33398 54386 33598 54398
rect 33398 54344 33598 54356
rect 33398 54310 33410 54344
rect 33586 54310 33598 54344
rect 33398 54298 33598 54310
rect 33398 54122 33598 54134
rect 33398 54088 33410 54122
rect 33586 54088 33598 54122
rect 33398 54076 33598 54088
rect 33398 54034 33598 54046
rect 33398 54000 33410 54034
rect 33586 54000 33598 54034
rect 33398 53988 33598 54000
rect 38388 54432 38588 54444
rect 38388 54398 38400 54432
rect 38576 54398 38588 54432
rect 38388 54386 38588 54398
rect 38388 54344 38588 54356
rect 38388 54310 38400 54344
rect 38576 54310 38588 54344
rect 38388 54298 38588 54310
rect 38388 54122 38588 54134
rect 38388 54088 38400 54122
rect 38576 54088 38588 54122
rect 38388 54076 38588 54088
rect 38388 54034 38588 54046
rect 38388 54000 38400 54034
rect 38576 54000 38588 54034
rect 38388 53988 38588 54000
rect 43378 54432 43578 54444
rect 43378 54398 43390 54432
rect 43566 54398 43578 54432
rect 43378 54386 43578 54398
rect 43378 54344 43578 54356
rect 43378 54310 43390 54344
rect 43566 54310 43578 54344
rect 43378 54298 43578 54310
rect 43378 54122 43578 54134
rect 43378 54088 43390 54122
rect 43566 54088 43578 54122
rect 43378 54076 43578 54088
rect 43378 54034 43578 54046
rect 43378 54000 43390 54034
rect 43566 54000 43578 54034
rect 43378 53988 43578 54000
rect 48368 54432 48568 54444
rect 48368 54398 48380 54432
rect 48556 54398 48568 54432
rect 48368 54386 48568 54398
rect 48368 54344 48568 54356
rect 48368 54310 48380 54344
rect 48556 54310 48568 54344
rect 48368 54298 48568 54310
rect 48368 54122 48568 54134
rect 48368 54088 48380 54122
rect 48556 54088 48568 54122
rect 48368 54076 48568 54088
rect 48368 54034 48568 54046
rect 48368 54000 48380 54034
rect 48556 54000 48568 54034
rect 48368 53988 48568 54000
rect 53358 54432 53558 54444
rect 53358 54398 53370 54432
rect 53546 54398 53558 54432
rect 53358 54386 53558 54398
rect 53358 54344 53558 54356
rect 53358 54310 53370 54344
rect 53546 54310 53558 54344
rect 53358 54298 53558 54310
rect 53358 54122 53558 54134
rect 53358 54088 53370 54122
rect 53546 54088 53558 54122
rect 53358 54076 53558 54088
rect 53358 54034 53558 54046
rect 53358 54000 53370 54034
rect 53546 54000 53558 54034
rect 53358 53988 53558 54000
rect 58348 54432 58548 54444
rect 58348 54398 58360 54432
rect 58536 54398 58548 54432
rect 58348 54386 58548 54398
rect 58348 54344 58548 54356
rect 58348 54310 58360 54344
rect 58536 54310 58548 54344
rect 58348 54298 58548 54310
rect 58348 54122 58548 54134
rect 58348 54088 58360 54122
rect 58536 54088 58548 54122
rect 58348 54076 58548 54088
rect 58348 54034 58548 54046
rect 58348 54000 58360 54034
rect 58536 54000 58548 54034
rect 58348 53988 58548 54000
rect 63338 54432 63538 54444
rect 63338 54398 63350 54432
rect 63526 54398 63538 54432
rect 63338 54386 63538 54398
rect 63338 54344 63538 54356
rect 63338 54310 63350 54344
rect 63526 54310 63538 54344
rect 63338 54298 63538 54310
rect 63338 54122 63538 54134
rect 63338 54088 63350 54122
rect 63526 54088 63538 54122
rect 63338 54076 63538 54088
rect 63338 54034 63538 54046
rect 63338 54000 63350 54034
rect 63526 54000 63538 54034
rect 63338 53988 63538 54000
rect 68328 54432 68528 54444
rect 68328 54398 68340 54432
rect 68516 54398 68528 54432
rect 68328 54386 68528 54398
rect 68328 54344 68528 54356
rect 68328 54310 68340 54344
rect 68516 54310 68528 54344
rect 68328 54298 68528 54310
rect 68328 54122 68528 54134
rect 68328 54088 68340 54122
rect 68516 54088 68528 54122
rect 68328 54076 68528 54088
rect 68328 54034 68528 54046
rect 68328 54000 68340 54034
rect 68516 54000 68528 54034
rect 68328 53988 68528 54000
rect 73318 54432 73518 54444
rect 73318 54398 73330 54432
rect 73506 54398 73518 54432
rect 73318 54386 73518 54398
rect 73318 54344 73518 54356
rect 73318 54310 73330 54344
rect 73506 54310 73518 54344
rect 73318 54298 73518 54310
rect 73318 54122 73518 54134
rect 73318 54088 73330 54122
rect 73506 54088 73518 54122
rect 73318 54076 73518 54088
rect 73318 54034 73518 54046
rect 73318 54000 73330 54034
rect 73506 54000 73518 54034
rect 73318 53988 73518 54000
rect 78308 54432 78508 54444
rect 78308 54398 78320 54432
rect 78496 54398 78508 54432
rect 78308 54386 78508 54398
rect 78308 54344 78508 54356
rect 78308 54310 78320 54344
rect 78496 54310 78508 54344
rect 78308 54298 78508 54310
rect 78308 54122 78508 54134
rect 78308 54088 78320 54122
rect 78496 54088 78508 54122
rect 78308 54076 78508 54088
rect 78308 54034 78508 54046
rect 78308 54000 78320 54034
rect 78496 54000 78508 54034
rect 78308 53988 78508 54000
rect 3458 52722 3658 52734
rect 3458 52688 3470 52722
rect 3646 52688 3658 52722
rect 3458 52676 3658 52688
rect 3458 52634 3658 52646
rect 3458 52600 3470 52634
rect 3646 52600 3658 52634
rect 3458 52588 3658 52600
rect 3458 52412 3658 52424
rect 3458 52378 3470 52412
rect 3646 52378 3658 52412
rect 3458 52366 3658 52378
rect 3458 52324 3658 52336
rect 3458 52290 3470 52324
rect 3646 52290 3658 52324
rect 3458 52278 3658 52290
rect 8448 52722 8648 52734
rect 8448 52688 8460 52722
rect 8636 52688 8648 52722
rect 8448 52676 8648 52688
rect 8448 52634 8648 52646
rect 8448 52600 8460 52634
rect 8636 52600 8648 52634
rect 8448 52588 8648 52600
rect 8448 52412 8648 52424
rect 8448 52378 8460 52412
rect 8636 52378 8648 52412
rect 8448 52366 8648 52378
rect 8448 52324 8648 52336
rect 8448 52290 8460 52324
rect 8636 52290 8648 52324
rect 8448 52278 8648 52290
rect 13438 52722 13638 52734
rect 13438 52688 13450 52722
rect 13626 52688 13638 52722
rect 13438 52676 13638 52688
rect 13438 52634 13638 52646
rect 13438 52600 13450 52634
rect 13626 52600 13638 52634
rect 13438 52588 13638 52600
rect 13438 52412 13638 52424
rect 13438 52378 13450 52412
rect 13626 52378 13638 52412
rect 13438 52366 13638 52378
rect 13438 52324 13638 52336
rect 13438 52290 13450 52324
rect 13626 52290 13638 52324
rect 13438 52278 13638 52290
rect 18428 52722 18628 52734
rect 18428 52688 18440 52722
rect 18616 52688 18628 52722
rect 18428 52676 18628 52688
rect 18428 52634 18628 52646
rect 18428 52600 18440 52634
rect 18616 52600 18628 52634
rect 18428 52588 18628 52600
rect 18428 52412 18628 52424
rect 18428 52378 18440 52412
rect 18616 52378 18628 52412
rect 18428 52366 18628 52378
rect 18428 52324 18628 52336
rect 18428 52290 18440 52324
rect 18616 52290 18628 52324
rect 18428 52278 18628 52290
rect 23418 52722 23618 52734
rect 23418 52688 23430 52722
rect 23606 52688 23618 52722
rect 23418 52676 23618 52688
rect 23418 52634 23618 52646
rect 23418 52600 23430 52634
rect 23606 52600 23618 52634
rect 23418 52588 23618 52600
rect 23418 52412 23618 52424
rect 23418 52378 23430 52412
rect 23606 52378 23618 52412
rect 23418 52366 23618 52378
rect 23418 52324 23618 52336
rect 23418 52290 23430 52324
rect 23606 52290 23618 52324
rect 23418 52278 23618 52290
rect 28408 52722 28608 52734
rect 28408 52688 28420 52722
rect 28596 52688 28608 52722
rect 28408 52676 28608 52688
rect 28408 52634 28608 52646
rect 28408 52600 28420 52634
rect 28596 52600 28608 52634
rect 28408 52588 28608 52600
rect 28408 52412 28608 52424
rect 28408 52378 28420 52412
rect 28596 52378 28608 52412
rect 28408 52366 28608 52378
rect 28408 52324 28608 52336
rect 28408 52290 28420 52324
rect 28596 52290 28608 52324
rect 28408 52278 28608 52290
rect 33398 52722 33598 52734
rect 33398 52688 33410 52722
rect 33586 52688 33598 52722
rect 33398 52676 33598 52688
rect 33398 52634 33598 52646
rect 33398 52600 33410 52634
rect 33586 52600 33598 52634
rect 33398 52588 33598 52600
rect 33398 52412 33598 52424
rect 33398 52378 33410 52412
rect 33586 52378 33598 52412
rect 33398 52366 33598 52378
rect 33398 52324 33598 52336
rect 33398 52290 33410 52324
rect 33586 52290 33598 52324
rect 33398 52278 33598 52290
rect 38388 52722 38588 52734
rect 38388 52688 38400 52722
rect 38576 52688 38588 52722
rect 38388 52676 38588 52688
rect 38388 52634 38588 52646
rect 38388 52600 38400 52634
rect 38576 52600 38588 52634
rect 38388 52588 38588 52600
rect 38388 52412 38588 52424
rect 38388 52378 38400 52412
rect 38576 52378 38588 52412
rect 38388 52366 38588 52378
rect 38388 52324 38588 52336
rect 38388 52290 38400 52324
rect 38576 52290 38588 52324
rect 38388 52278 38588 52290
rect 43378 52722 43578 52734
rect 43378 52688 43390 52722
rect 43566 52688 43578 52722
rect 43378 52676 43578 52688
rect 43378 52634 43578 52646
rect 43378 52600 43390 52634
rect 43566 52600 43578 52634
rect 43378 52588 43578 52600
rect 43378 52412 43578 52424
rect 43378 52378 43390 52412
rect 43566 52378 43578 52412
rect 43378 52366 43578 52378
rect 43378 52324 43578 52336
rect 43378 52290 43390 52324
rect 43566 52290 43578 52324
rect 43378 52278 43578 52290
rect 48368 52722 48568 52734
rect 48368 52688 48380 52722
rect 48556 52688 48568 52722
rect 48368 52676 48568 52688
rect 48368 52634 48568 52646
rect 48368 52600 48380 52634
rect 48556 52600 48568 52634
rect 48368 52588 48568 52600
rect 48368 52412 48568 52424
rect 48368 52378 48380 52412
rect 48556 52378 48568 52412
rect 48368 52366 48568 52378
rect 48368 52324 48568 52336
rect 48368 52290 48380 52324
rect 48556 52290 48568 52324
rect 48368 52278 48568 52290
rect 53358 52722 53558 52734
rect 53358 52688 53370 52722
rect 53546 52688 53558 52722
rect 53358 52676 53558 52688
rect 53358 52634 53558 52646
rect 53358 52600 53370 52634
rect 53546 52600 53558 52634
rect 53358 52588 53558 52600
rect 53358 52412 53558 52424
rect 53358 52378 53370 52412
rect 53546 52378 53558 52412
rect 53358 52366 53558 52378
rect 53358 52324 53558 52336
rect 53358 52290 53370 52324
rect 53546 52290 53558 52324
rect 53358 52278 53558 52290
rect 58348 52722 58548 52734
rect 58348 52688 58360 52722
rect 58536 52688 58548 52722
rect 58348 52676 58548 52688
rect 58348 52634 58548 52646
rect 58348 52600 58360 52634
rect 58536 52600 58548 52634
rect 58348 52588 58548 52600
rect 58348 52412 58548 52424
rect 58348 52378 58360 52412
rect 58536 52378 58548 52412
rect 58348 52366 58548 52378
rect 58348 52324 58548 52336
rect 58348 52290 58360 52324
rect 58536 52290 58548 52324
rect 58348 52278 58548 52290
rect 63338 52722 63538 52734
rect 63338 52688 63350 52722
rect 63526 52688 63538 52722
rect 63338 52676 63538 52688
rect 63338 52634 63538 52646
rect 63338 52600 63350 52634
rect 63526 52600 63538 52634
rect 63338 52588 63538 52600
rect 63338 52412 63538 52424
rect 63338 52378 63350 52412
rect 63526 52378 63538 52412
rect 63338 52366 63538 52378
rect 63338 52324 63538 52336
rect 63338 52290 63350 52324
rect 63526 52290 63538 52324
rect 63338 52278 63538 52290
rect 68328 52722 68528 52734
rect 68328 52688 68340 52722
rect 68516 52688 68528 52722
rect 68328 52676 68528 52688
rect 68328 52634 68528 52646
rect 68328 52600 68340 52634
rect 68516 52600 68528 52634
rect 68328 52588 68528 52600
rect 68328 52412 68528 52424
rect 68328 52378 68340 52412
rect 68516 52378 68528 52412
rect 68328 52366 68528 52378
rect 68328 52324 68528 52336
rect 68328 52290 68340 52324
rect 68516 52290 68528 52324
rect 68328 52278 68528 52290
rect 73318 52722 73518 52734
rect 73318 52688 73330 52722
rect 73506 52688 73518 52722
rect 73318 52676 73518 52688
rect 73318 52634 73518 52646
rect 73318 52600 73330 52634
rect 73506 52600 73518 52634
rect 73318 52588 73518 52600
rect 73318 52412 73518 52424
rect 73318 52378 73330 52412
rect 73506 52378 73518 52412
rect 73318 52366 73518 52378
rect 73318 52324 73518 52336
rect 73318 52290 73330 52324
rect 73506 52290 73518 52324
rect 73318 52278 73518 52290
rect 78308 52722 78508 52734
rect 78308 52688 78320 52722
rect 78496 52688 78508 52722
rect 78308 52676 78508 52688
rect 78308 52634 78508 52646
rect 78308 52600 78320 52634
rect 78496 52600 78508 52634
rect 78308 52588 78508 52600
rect 78308 52412 78508 52424
rect 78308 52378 78320 52412
rect 78496 52378 78508 52412
rect 78308 52366 78508 52378
rect 78308 52324 78508 52336
rect 78308 52290 78320 52324
rect 78496 52290 78508 52324
rect 78308 52278 78508 52290
rect 3458 51012 3658 51024
rect 3458 50978 3470 51012
rect 3646 50978 3658 51012
rect 3458 50966 3658 50978
rect 3458 50924 3658 50936
rect 3458 50890 3470 50924
rect 3646 50890 3658 50924
rect 3458 50878 3658 50890
rect 3458 50702 3658 50714
rect 3458 50668 3470 50702
rect 3646 50668 3658 50702
rect 3458 50656 3658 50668
rect 3458 50614 3658 50626
rect 3458 50580 3470 50614
rect 3646 50580 3658 50614
rect 3458 50568 3658 50580
rect 8448 51012 8648 51024
rect 8448 50978 8460 51012
rect 8636 50978 8648 51012
rect 8448 50966 8648 50978
rect 8448 50924 8648 50936
rect 8448 50890 8460 50924
rect 8636 50890 8648 50924
rect 8448 50878 8648 50890
rect 8448 50702 8648 50714
rect 8448 50668 8460 50702
rect 8636 50668 8648 50702
rect 8448 50656 8648 50668
rect 8448 50614 8648 50626
rect 8448 50580 8460 50614
rect 8636 50580 8648 50614
rect 8448 50568 8648 50580
rect 13438 51012 13638 51024
rect 13438 50978 13450 51012
rect 13626 50978 13638 51012
rect 13438 50966 13638 50978
rect 13438 50924 13638 50936
rect 13438 50890 13450 50924
rect 13626 50890 13638 50924
rect 13438 50878 13638 50890
rect 13438 50702 13638 50714
rect 13438 50668 13450 50702
rect 13626 50668 13638 50702
rect 13438 50656 13638 50668
rect 13438 50614 13638 50626
rect 13438 50580 13450 50614
rect 13626 50580 13638 50614
rect 13438 50568 13638 50580
rect 18428 51012 18628 51024
rect 18428 50978 18440 51012
rect 18616 50978 18628 51012
rect 18428 50966 18628 50978
rect 18428 50924 18628 50936
rect 18428 50890 18440 50924
rect 18616 50890 18628 50924
rect 18428 50878 18628 50890
rect 18428 50702 18628 50714
rect 18428 50668 18440 50702
rect 18616 50668 18628 50702
rect 18428 50656 18628 50668
rect 18428 50614 18628 50626
rect 18428 50580 18440 50614
rect 18616 50580 18628 50614
rect 18428 50568 18628 50580
rect 23418 51012 23618 51024
rect 23418 50978 23430 51012
rect 23606 50978 23618 51012
rect 23418 50966 23618 50978
rect 23418 50924 23618 50936
rect 23418 50890 23430 50924
rect 23606 50890 23618 50924
rect 23418 50878 23618 50890
rect 23418 50702 23618 50714
rect 23418 50668 23430 50702
rect 23606 50668 23618 50702
rect 23418 50656 23618 50668
rect 23418 50614 23618 50626
rect 23418 50580 23430 50614
rect 23606 50580 23618 50614
rect 23418 50568 23618 50580
rect 28408 51012 28608 51024
rect 28408 50978 28420 51012
rect 28596 50978 28608 51012
rect 28408 50966 28608 50978
rect 28408 50924 28608 50936
rect 28408 50890 28420 50924
rect 28596 50890 28608 50924
rect 28408 50878 28608 50890
rect 28408 50702 28608 50714
rect 28408 50668 28420 50702
rect 28596 50668 28608 50702
rect 28408 50656 28608 50668
rect 28408 50614 28608 50626
rect 28408 50580 28420 50614
rect 28596 50580 28608 50614
rect 28408 50568 28608 50580
rect 33398 51012 33598 51024
rect 33398 50978 33410 51012
rect 33586 50978 33598 51012
rect 33398 50966 33598 50978
rect 33398 50924 33598 50936
rect 33398 50890 33410 50924
rect 33586 50890 33598 50924
rect 33398 50878 33598 50890
rect 33398 50702 33598 50714
rect 33398 50668 33410 50702
rect 33586 50668 33598 50702
rect 33398 50656 33598 50668
rect 33398 50614 33598 50626
rect 33398 50580 33410 50614
rect 33586 50580 33598 50614
rect 33398 50568 33598 50580
rect 38388 51012 38588 51024
rect 38388 50978 38400 51012
rect 38576 50978 38588 51012
rect 38388 50966 38588 50978
rect 38388 50924 38588 50936
rect 38388 50890 38400 50924
rect 38576 50890 38588 50924
rect 38388 50878 38588 50890
rect 38388 50702 38588 50714
rect 38388 50668 38400 50702
rect 38576 50668 38588 50702
rect 38388 50656 38588 50668
rect 38388 50614 38588 50626
rect 38388 50580 38400 50614
rect 38576 50580 38588 50614
rect 38388 50568 38588 50580
rect 43378 51012 43578 51024
rect 43378 50978 43390 51012
rect 43566 50978 43578 51012
rect 43378 50966 43578 50978
rect 43378 50924 43578 50936
rect 43378 50890 43390 50924
rect 43566 50890 43578 50924
rect 43378 50878 43578 50890
rect 43378 50702 43578 50714
rect 43378 50668 43390 50702
rect 43566 50668 43578 50702
rect 43378 50656 43578 50668
rect 43378 50614 43578 50626
rect 43378 50580 43390 50614
rect 43566 50580 43578 50614
rect 43378 50568 43578 50580
rect 48368 51012 48568 51024
rect 48368 50978 48380 51012
rect 48556 50978 48568 51012
rect 48368 50966 48568 50978
rect 48368 50924 48568 50936
rect 48368 50890 48380 50924
rect 48556 50890 48568 50924
rect 48368 50878 48568 50890
rect 48368 50702 48568 50714
rect 48368 50668 48380 50702
rect 48556 50668 48568 50702
rect 48368 50656 48568 50668
rect 48368 50614 48568 50626
rect 48368 50580 48380 50614
rect 48556 50580 48568 50614
rect 48368 50568 48568 50580
rect 53358 51012 53558 51024
rect 53358 50978 53370 51012
rect 53546 50978 53558 51012
rect 53358 50966 53558 50978
rect 53358 50924 53558 50936
rect 53358 50890 53370 50924
rect 53546 50890 53558 50924
rect 53358 50878 53558 50890
rect 53358 50702 53558 50714
rect 53358 50668 53370 50702
rect 53546 50668 53558 50702
rect 53358 50656 53558 50668
rect 53358 50614 53558 50626
rect 53358 50580 53370 50614
rect 53546 50580 53558 50614
rect 53358 50568 53558 50580
rect 58348 51012 58548 51024
rect 58348 50978 58360 51012
rect 58536 50978 58548 51012
rect 58348 50966 58548 50978
rect 58348 50924 58548 50936
rect 58348 50890 58360 50924
rect 58536 50890 58548 50924
rect 58348 50878 58548 50890
rect 58348 50702 58548 50714
rect 58348 50668 58360 50702
rect 58536 50668 58548 50702
rect 58348 50656 58548 50668
rect 58348 50614 58548 50626
rect 58348 50580 58360 50614
rect 58536 50580 58548 50614
rect 58348 50568 58548 50580
rect 63338 51012 63538 51024
rect 63338 50978 63350 51012
rect 63526 50978 63538 51012
rect 63338 50966 63538 50978
rect 63338 50924 63538 50936
rect 63338 50890 63350 50924
rect 63526 50890 63538 50924
rect 63338 50878 63538 50890
rect 63338 50702 63538 50714
rect 63338 50668 63350 50702
rect 63526 50668 63538 50702
rect 63338 50656 63538 50668
rect 63338 50614 63538 50626
rect 63338 50580 63350 50614
rect 63526 50580 63538 50614
rect 63338 50568 63538 50580
rect 68328 51012 68528 51024
rect 68328 50978 68340 51012
rect 68516 50978 68528 51012
rect 68328 50966 68528 50978
rect 68328 50924 68528 50936
rect 68328 50890 68340 50924
rect 68516 50890 68528 50924
rect 68328 50878 68528 50890
rect 68328 50702 68528 50714
rect 68328 50668 68340 50702
rect 68516 50668 68528 50702
rect 68328 50656 68528 50668
rect 68328 50614 68528 50626
rect 68328 50580 68340 50614
rect 68516 50580 68528 50614
rect 68328 50568 68528 50580
rect 73318 51012 73518 51024
rect 73318 50978 73330 51012
rect 73506 50978 73518 51012
rect 73318 50966 73518 50978
rect 73318 50924 73518 50936
rect 73318 50890 73330 50924
rect 73506 50890 73518 50924
rect 73318 50878 73518 50890
rect 73318 50702 73518 50714
rect 73318 50668 73330 50702
rect 73506 50668 73518 50702
rect 73318 50656 73518 50668
rect 73318 50614 73518 50626
rect 73318 50580 73330 50614
rect 73506 50580 73518 50614
rect 73318 50568 73518 50580
rect 78308 51012 78508 51024
rect 78308 50978 78320 51012
rect 78496 50978 78508 51012
rect 78308 50966 78508 50978
rect 78308 50924 78508 50936
rect 78308 50890 78320 50924
rect 78496 50890 78508 50924
rect 78308 50878 78508 50890
rect 78308 50702 78508 50714
rect 78308 50668 78320 50702
rect 78496 50668 78508 50702
rect 78308 50656 78508 50668
rect 78308 50614 78508 50626
rect 78308 50580 78320 50614
rect 78496 50580 78508 50614
rect 78308 50568 78508 50580
rect 3458 49302 3658 49314
rect 3458 49268 3470 49302
rect 3646 49268 3658 49302
rect 3458 49256 3658 49268
rect 3458 49214 3658 49226
rect 3458 49180 3470 49214
rect 3646 49180 3658 49214
rect 3458 49168 3658 49180
rect 3458 48992 3658 49004
rect 3458 48958 3470 48992
rect 3646 48958 3658 48992
rect 3458 48946 3658 48958
rect 3458 48904 3658 48916
rect 3458 48870 3470 48904
rect 3646 48870 3658 48904
rect 3458 48858 3658 48870
rect 8448 49302 8648 49314
rect 8448 49268 8460 49302
rect 8636 49268 8648 49302
rect 8448 49256 8648 49268
rect 8448 49214 8648 49226
rect 8448 49180 8460 49214
rect 8636 49180 8648 49214
rect 8448 49168 8648 49180
rect 8448 48992 8648 49004
rect 8448 48958 8460 48992
rect 8636 48958 8648 48992
rect 8448 48946 8648 48958
rect 8448 48904 8648 48916
rect 8448 48870 8460 48904
rect 8636 48870 8648 48904
rect 8448 48858 8648 48870
rect 13438 49302 13638 49314
rect 13438 49268 13450 49302
rect 13626 49268 13638 49302
rect 13438 49256 13638 49268
rect 13438 49214 13638 49226
rect 13438 49180 13450 49214
rect 13626 49180 13638 49214
rect 13438 49168 13638 49180
rect 13438 48992 13638 49004
rect 13438 48958 13450 48992
rect 13626 48958 13638 48992
rect 13438 48946 13638 48958
rect 13438 48904 13638 48916
rect 13438 48870 13450 48904
rect 13626 48870 13638 48904
rect 13438 48858 13638 48870
rect 18428 49302 18628 49314
rect 18428 49268 18440 49302
rect 18616 49268 18628 49302
rect 18428 49256 18628 49268
rect 18428 49214 18628 49226
rect 18428 49180 18440 49214
rect 18616 49180 18628 49214
rect 18428 49168 18628 49180
rect 18428 48992 18628 49004
rect 18428 48958 18440 48992
rect 18616 48958 18628 48992
rect 18428 48946 18628 48958
rect 18428 48904 18628 48916
rect 18428 48870 18440 48904
rect 18616 48870 18628 48904
rect 18428 48858 18628 48870
rect 23418 49302 23618 49314
rect 23418 49268 23430 49302
rect 23606 49268 23618 49302
rect 23418 49256 23618 49268
rect 23418 49214 23618 49226
rect 23418 49180 23430 49214
rect 23606 49180 23618 49214
rect 23418 49168 23618 49180
rect 23418 48992 23618 49004
rect 23418 48958 23430 48992
rect 23606 48958 23618 48992
rect 23418 48946 23618 48958
rect 23418 48904 23618 48916
rect 23418 48870 23430 48904
rect 23606 48870 23618 48904
rect 23418 48858 23618 48870
rect 28408 49302 28608 49314
rect 28408 49268 28420 49302
rect 28596 49268 28608 49302
rect 28408 49256 28608 49268
rect 28408 49214 28608 49226
rect 28408 49180 28420 49214
rect 28596 49180 28608 49214
rect 28408 49168 28608 49180
rect 28408 48992 28608 49004
rect 28408 48958 28420 48992
rect 28596 48958 28608 48992
rect 28408 48946 28608 48958
rect 28408 48904 28608 48916
rect 28408 48870 28420 48904
rect 28596 48870 28608 48904
rect 28408 48858 28608 48870
rect 33398 49302 33598 49314
rect 33398 49268 33410 49302
rect 33586 49268 33598 49302
rect 33398 49256 33598 49268
rect 33398 49214 33598 49226
rect 33398 49180 33410 49214
rect 33586 49180 33598 49214
rect 33398 49168 33598 49180
rect 33398 48992 33598 49004
rect 33398 48958 33410 48992
rect 33586 48958 33598 48992
rect 33398 48946 33598 48958
rect 33398 48904 33598 48916
rect 33398 48870 33410 48904
rect 33586 48870 33598 48904
rect 33398 48858 33598 48870
rect 38388 49302 38588 49314
rect 38388 49268 38400 49302
rect 38576 49268 38588 49302
rect 38388 49256 38588 49268
rect 38388 49214 38588 49226
rect 38388 49180 38400 49214
rect 38576 49180 38588 49214
rect 38388 49168 38588 49180
rect 38388 48992 38588 49004
rect 38388 48958 38400 48992
rect 38576 48958 38588 48992
rect 38388 48946 38588 48958
rect 38388 48904 38588 48916
rect 38388 48870 38400 48904
rect 38576 48870 38588 48904
rect 38388 48858 38588 48870
rect 43378 49302 43578 49314
rect 43378 49268 43390 49302
rect 43566 49268 43578 49302
rect 43378 49256 43578 49268
rect 43378 49214 43578 49226
rect 43378 49180 43390 49214
rect 43566 49180 43578 49214
rect 43378 49168 43578 49180
rect 43378 48992 43578 49004
rect 43378 48958 43390 48992
rect 43566 48958 43578 48992
rect 43378 48946 43578 48958
rect 43378 48904 43578 48916
rect 43378 48870 43390 48904
rect 43566 48870 43578 48904
rect 43378 48858 43578 48870
rect 48368 49302 48568 49314
rect 48368 49268 48380 49302
rect 48556 49268 48568 49302
rect 48368 49256 48568 49268
rect 48368 49214 48568 49226
rect 48368 49180 48380 49214
rect 48556 49180 48568 49214
rect 48368 49168 48568 49180
rect 48368 48992 48568 49004
rect 48368 48958 48380 48992
rect 48556 48958 48568 48992
rect 48368 48946 48568 48958
rect 48368 48904 48568 48916
rect 48368 48870 48380 48904
rect 48556 48870 48568 48904
rect 48368 48858 48568 48870
rect 53358 49302 53558 49314
rect 53358 49268 53370 49302
rect 53546 49268 53558 49302
rect 53358 49256 53558 49268
rect 53358 49214 53558 49226
rect 53358 49180 53370 49214
rect 53546 49180 53558 49214
rect 53358 49168 53558 49180
rect 53358 48992 53558 49004
rect 53358 48958 53370 48992
rect 53546 48958 53558 48992
rect 53358 48946 53558 48958
rect 53358 48904 53558 48916
rect 53358 48870 53370 48904
rect 53546 48870 53558 48904
rect 53358 48858 53558 48870
rect 58348 49302 58548 49314
rect 58348 49268 58360 49302
rect 58536 49268 58548 49302
rect 58348 49256 58548 49268
rect 58348 49214 58548 49226
rect 58348 49180 58360 49214
rect 58536 49180 58548 49214
rect 58348 49168 58548 49180
rect 58348 48992 58548 49004
rect 58348 48958 58360 48992
rect 58536 48958 58548 48992
rect 58348 48946 58548 48958
rect 58348 48904 58548 48916
rect 58348 48870 58360 48904
rect 58536 48870 58548 48904
rect 58348 48858 58548 48870
rect 63338 49302 63538 49314
rect 63338 49268 63350 49302
rect 63526 49268 63538 49302
rect 63338 49256 63538 49268
rect 63338 49214 63538 49226
rect 63338 49180 63350 49214
rect 63526 49180 63538 49214
rect 63338 49168 63538 49180
rect 63338 48992 63538 49004
rect 63338 48958 63350 48992
rect 63526 48958 63538 48992
rect 63338 48946 63538 48958
rect 63338 48904 63538 48916
rect 63338 48870 63350 48904
rect 63526 48870 63538 48904
rect 63338 48858 63538 48870
rect 68328 49302 68528 49314
rect 68328 49268 68340 49302
rect 68516 49268 68528 49302
rect 68328 49256 68528 49268
rect 68328 49214 68528 49226
rect 68328 49180 68340 49214
rect 68516 49180 68528 49214
rect 68328 49168 68528 49180
rect 68328 48992 68528 49004
rect 68328 48958 68340 48992
rect 68516 48958 68528 48992
rect 68328 48946 68528 48958
rect 68328 48904 68528 48916
rect 68328 48870 68340 48904
rect 68516 48870 68528 48904
rect 68328 48858 68528 48870
rect 73318 49302 73518 49314
rect 73318 49268 73330 49302
rect 73506 49268 73518 49302
rect 73318 49256 73518 49268
rect 73318 49214 73518 49226
rect 73318 49180 73330 49214
rect 73506 49180 73518 49214
rect 73318 49168 73518 49180
rect 73318 48992 73518 49004
rect 73318 48958 73330 48992
rect 73506 48958 73518 48992
rect 73318 48946 73518 48958
rect 73318 48904 73518 48916
rect 73318 48870 73330 48904
rect 73506 48870 73518 48904
rect 73318 48858 73518 48870
rect 78308 49302 78508 49314
rect 78308 49268 78320 49302
rect 78496 49268 78508 49302
rect 78308 49256 78508 49268
rect 78308 49214 78508 49226
rect 78308 49180 78320 49214
rect 78496 49180 78508 49214
rect 78308 49168 78508 49180
rect 78308 48992 78508 49004
rect 78308 48958 78320 48992
rect 78496 48958 78508 48992
rect 78308 48946 78508 48958
rect 78308 48904 78508 48916
rect 78308 48870 78320 48904
rect 78496 48870 78508 48904
rect 78308 48858 78508 48870
rect 3458 47592 3658 47604
rect 3458 47558 3470 47592
rect 3646 47558 3658 47592
rect 3458 47546 3658 47558
rect 3458 47504 3658 47516
rect 3458 47470 3470 47504
rect 3646 47470 3658 47504
rect 3458 47458 3658 47470
rect 3458 47282 3658 47294
rect 3458 47248 3470 47282
rect 3646 47248 3658 47282
rect 3458 47236 3658 47248
rect 3458 47194 3658 47206
rect 3458 47160 3470 47194
rect 3646 47160 3658 47194
rect 3458 47148 3658 47160
rect 8448 47592 8648 47604
rect 8448 47558 8460 47592
rect 8636 47558 8648 47592
rect 8448 47546 8648 47558
rect 8448 47504 8648 47516
rect 8448 47470 8460 47504
rect 8636 47470 8648 47504
rect 8448 47458 8648 47470
rect 8448 47282 8648 47294
rect 8448 47248 8460 47282
rect 8636 47248 8648 47282
rect 8448 47236 8648 47248
rect 8448 47194 8648 47206
rect 8448 47160 8460 47194
rect 8636 47160 8648 47194
rect 8448 47148 8648 47160
rect 13438 47592 13638 47604
rect 13438 47558 13450 47592
rect 13626 47558 13638 47592
rect 13438 47546 13638 47558
rect 13438 47504 13638 47516
rect 13438 47470 13450 47504
rect 13626 47470 13638 47504
rect 13438 47458 13638 47470
rect 13438 47282 13638 47294
rect 13438 47248 13450 47282
rect 13626 47248 13638 47282
rect 13438 47236 13638 47248
rect 13438 47194 13638 47206
rect 13438 47160 13450 47194
rect 13626 47160 13638 47194
rect 13438 47148 13638 47160
rect 18428 47592 18628 47604
rect 18428 47558 18440 47592
rect 18616 47558 18628 47592
rect 18428 47546 18628 47558
rect 18428 47504 18628 47516
rect 18428 47470 18440 47504
rect 18616 47470 18628 47504
rect 18428 47458 18628 47470
rect 18428 47282 18628 47294
rect 18428 47248 18440 47282
rect 18616 47248 18628 47282
rect 18428 47236 18628 47248
rect 18428 47194 18628 47206
rect 18428 47160 18440 47194
rect 18616 47160 18628 47194
rect 18428 47148 18628 47160
rect 23418 47592 23618 47604
rect 23418 47558 23430 47592
rect 23606 47558 23618 47592
rect 23418 47546 23618 47558
rect 23418 47504 23618 47516
rect 23418 47470 23430 47504
rect 23606 47470 23618 47504
rect 23418 47458 23618 47470
rect 23418 47282 23618 47294
rect 23418 47248 23430 47282
rect 23606 47248 23618 47282
rect 23418 47236 23618 47248
rect 23418 47194 23618 47206
rect 23418 47160 23430 47194
rect 23606 47160 23618 47194
rect 23418 47148 23618 47160
rect 28408 47592 28608 47604
rect 28408 47558 28420 47592
rect 28596 47558 28608 47592
rect 28408 47546 28608 47558
rect 28408 47504 28608 47516
rect 28408 47470 28420 47504
rect 28596 47470 28608 47504
rect 28408 47458 28608 47470
rect 28408 47282 28608 47294
rect 28408 47248 28420 47282
rect 28596 47248 28608 47282
rect 28408 47236 28608 47248
rect 28408 47194 28608 47206
rect 28408 47160 28420 47194
rect 28596 47160 28608 47194
rect 28408 47148 28608 47160
rect 33398 47592 33598 47604
rect 33398 47558 33410 47592
rect 33586 47558 33598 47592
rect 33398 47546 33598 47558
rect 33398 47504 33598 47516
rect 33398 47470 33410 47504
rect 33586 47470 33598 47504
rect 33398 47458 33598 47470
rect 33398 47282 33598 47294
rect 33398 47248 33410 47282
rect 33586 47248 33598 47282
rect 33398 47236 33598 47248
rect 33398 47194 33598 47206
rect 33398 47160 33410 47194
rect 33586 47160 33598 47194
rect 33398 47148 33598 47160
rect 38388 47592 38588 47604
rect 38388 47558 38400 47592
rect 38576 47558 38588 47592
rect 38388 47546 38588 47558
rect 38388 47504 38588 47516
rect 38388 47470 38400 47504
rect 38576 47470 38588 47504
rect 38388 47458 38588 47470
rect 38388 47282 38588 47294
rect 38388 47248 38400 47282
rect 38576 47248 38588 47282
rect 38388 47236 38588 47248
rect 38388 47194 38588 47206
rect 38388 47160 38400 47194
rect 38576 47160 38588 47194
rect 38388 47148 38588 47160
rect 43378 47592 43578 47604
rect 43378 47558 43390 47592
rect 43566 47558 43578 47592
rect 43378 47546 43578 47558
rect 43378 47504 43578 47516
rect 43378 47470 43390 47504
rect 43566 47470 43578 47504
rect 43378 47458 43578 47470
rect 43378 47282 43578 47294
rect 43378 47248 43390 47282
rect 43566 47248 43578 47282
rect 43378 47236 43578 47248
rect 43378 47194 43578 47206
rect 43378 47160 43390 47194
rect 43566 47160 43578 47194
rect 43378 47148 43578 47160
rect 48368 47592 48568 47604
rect 48368 47558 48380 47592
rect 48556 47558 48568 47592
rect 48368 47546 48568 47558
rect 48368 47504 48568 47516
rect 48368 47470 48380 47504
rect 48556 47470 48568 47504
rect 48368 47458 48568 47470
rect 48368 47282 48568 47294
rect 48368 47248 48380 47282
rect 48556 47248 48568 47282
rect 48368 47236 48568 47248
rect 48368 47194 48568 47206
rect 48368 47160 48380 47194
rect 48556 47160 48568 47194
rect 48368 47148 48568 47160
rect 53358 47592 53558 47604
rect 53358 47558 53370 47592
rect 53546 47558 53558 47592
rect 53358 47546 53558 47558
rect 53358 47504 53558 47516
rect 53358 47470 53370 47504
rect 53546 47470 53558 47504
rect 53358 47458 53558 47470
rect 53358 47282 53558 47294
rect 53358 47248 53370 47282
rect 53546 47248 53558 47282
rect 53358 47236 53558 47248
rect 53358 47194 53558 47206
rect 53358 47160 53370 47194
rect 53546 47160 53558 47194
rect 53358 47148 53558 47160
rect 58348 47592 58548 47604
rect 58348 47558 58360 47592
rect 58536 47558 58548 47592
rect 58348 47546 58548 47558
rect 58348 47504 58548 47516
rect 58348 47470 58360 47504
rect 58536 47470 58548 47504
rect 58348 47458 58548 47470
rect 58348 47282 58548 47294
rect 58348 47248 58360 47282
rect 58536 47248 58548 47282
rect 58348 47236 58548 47248
rect 58348 47194 58548 47206
rect 58348 47160 58360 47194
rect 58536 47160 58548 47194
rect 58348 47148 58548 47160
rect 63338 47592 63538 47604
rect 63338 47558 63350 47592
rect 63526 47558 63538 47592
rect 63338 47546 63538 47558
rect 63338 47504 63538 47516
rect 63338 47470 63350 47504
rect 63526 47470 63538 47504
rect 63338 47458 63538 47470
rect 63338 47282 63538 47294
rect 63338 47248 63350 47282
rect 63526 47248 63538 47282
rect 63338 47236 63538 47248
rect 63338 47194 63538 47206
rect 63338 47160 63350 47194
rect 63526 47160 63538 47194
rect 63338 47148 63538 47160
rect 68328 47592 68528 47604
rect 68328 47558 68340 47592
rect 68516 47558 68528 47592
rect 68328 47546 68528 47558
rect 68328 47504 68528 47516
rect 68328 47470 68340 47504
rect 68516 47470 68528 47504
rect 68328 47458 68528 47470
rect 68328 47282 68528 47294
rect 68328 47248 68340 47282
rect 68516 47248 68528 47282
rect 68328 47236 68528 47248
rect 68328 47194 68528 47206
rect 68328 47160 68340 47194
rect 68516 47160 68528 47194
rect 68328 47148 68528 47160
rect 73318 47592 73518 47604
rect 73318 47558 73330 47592
rect 73506 47558 73518 47592
rect 73318 47546 73518 47558
rect 73318 47504 73518 47516
rect 73318 47470 73330 47504
rect 73506 47470 73518 47504
rect 73318 47458 73518 47470
rect 73318 47282 73518 47294
rect 73318 47248 73330 47282
rect 73506 47248 73518 47282
rect 73318 47236 73518 47248
rect 73318 47194 73518 47206
rect 73318 47160 73330 47194
rect 73506 47160 73518 47194
rect 73318 47148 73518 47160
rect 78308 47592 78508 47604
rect 78308 47558 78320 47592
rect 78496 47558 78508 47592
rect 78308 47546 78508 47558
rect 78308 47504 78508 47516
rect 78308 47470 78320 47504
rect 78496 47470 78508 47504
rect 78308 47458 78508 47470
rect 78308 47282 78508 47294
rect 78308 47248 78320 47282
rect 78496 47248 78508 47282
rect 78308 47236 78508 47248
rect 78308 47194 78508 47206
rect 78308 47160 78320 47194
rect 78496 47160 78508 47194
rect 78308 47148 78508 47160
rect 3458 45882 3658 45894
rect 3458 45848 3470 45882
rect 3646 45848 3658 45882
rect 3458 45836 3658 45848
rect 3458 45794 3658 45806
rect 3458 45760 3470 45794
rect 3646 45760 3658 45794
rect 3458 45748 3658 45760
rect 3458 45572 3658 45584
rect 3458 45538 3470 45572
rect 3646 45538 3658 45572
rect 3458 45526 3658 45538
rect 3458 45484 3658 45496
rect 3458 45450 3470 45484
rect 3646 45450 3658 45484
rect 3458 45438 3658 45450
rect 8448 45882 8648 45894
rect 8448 45848 8460 45882
rect 8636 45848 8648 45882
rect 8448 45836 8648 45848
rect 8448 45794 8648 45806
rect 8448 45760 8460 45794
rect 8636 45760 8648 45794
rect 8448 45748 8648 45760
rect 8448 45572 8648 45584
rect 8448 45538 8460 45572
rect 8636 45538 8648 45572
rect 8448 45526 8648 45538
rect 8448 45484 8648 45496
rect 8448 45450 8460 45484
rect 8636 45450 8648 45484
rect 8448 45438 8648 45450
rect 13438 45882 13638 45894
rect 13438 45848 13450 45882
rect 13626 45848 13638 45882
rect 13438 45836 13638 45848
rect 13438 45794 13638 45806
rect 13438 45760 13450 45794
rect 13626 45760 13638 45794
rect 13438 45748 13638 45760
rect 13438 45572 13638 45584
rect 13438 45538 13450 45572
rect 13626 45538 13638 45572
rect 13438 45526 13638 45538
rect 13438 45484 13638 45496
rect 13438 45450 13450 45484
rect 13626 45450 13638 45484
rect 13438 45438 13638 45450
rect 18428 45882 18628 45894
rect 18428 45848 18440 45882
rect 18616 45848 18628 45882
rect 18428 45836 18628 45848
rect 18428 45794 18628 45806
rect 18428 45760 18440 45794
rect 18616 45760 18628 45794
rect 18428 45748 18628 45760
rect 18428 45572 18628 45584
rect 18428 45538 18440 45572
rect 18616 45538 18628 45572
rect 18428 45526 18628 45538
rect 18428 45484 18628 45496
rect 18428 45450 18440 45484
rect 18616 45450 18628 45484
rect 18428 45438 18628 45450
rect 23418 45882 23618 45894
rect 23418 45848 23430 45882
rect 23606 45848 23618 45882
rect 23418 45836 23618 45848
rect 23418 45794 23618 45806
rect 23418 45760 23430 45794
rect 23606 45760 23618 45794
rect 23418 45748 23618 45760
rect 23418 45572 23618 45584
rect 23418 45538 23430 45572
rect 23606 45538 23618 45572
rect 23418 45526 23618 45538
rect 23418 45484 23618 45496
rect 23418 45450 23430 45484
rect 23606 45450 23618 45484
rect 23418 45438 23618 45450
rect 28408 45882 28608 45894
rect 28408 45848 28420 45882
rect 28596 45848 28608 45882
rect 28408 45836 28608 45848
rect 28408 45794 28608 45806
rect 28408 45760 28420 45794
rect 28596 45760 28608 45794
rect 28408 45748 28608 45760
rect 28408 45572 28608 45584
rect 28408 45538 28420 45572
rect 28596 45538 28608 45572
rect 28408 45526 28608 45538
rect 28408 45484 28608 45496
rect 28408 45450 28420 45484
rect 28596 45450 28608 45484
rect 28408 45438 28608 45450
rect 33398 45882 33598 45894
rect 33398 45848 33410 45882
rect 33586 45848 33598 45882
rect 33398 45836 33598 45848
rect 33398 45794 33598 45806
rect 33398 45760 33410 45794
rect 33586 45760 33598 45794
rect 33398 45748 33598 45760
rect 33398 45572 33598 45584
rect 33398 45538 33410 45572
rect 33586 45538 33598 45572
rect 33398 45526 33598 45538
rect 33398 45484 33598 45496
rect 33398 45450 33410 45484
rect 33586 45450 33598 45484
rect 33398 45438 33598 45450
rect 38388 45882 38588 45894
rect 38388 45848 38400 45882
rect 38576 45848 38588 45882
rect 38388 45836 38588 45848
rect 38388 45794 38588 45806
rect 38388 45760 38400 45794
rect 38576 45760 38588 45794
rect 38388 45748 38588 45760
rect 38388 45572 38588 45584
rect 38388 45538 38400 45572
rect 38576 45538 38588 45572
rect 38388 45526 38588 45538
rect 38388 45484 38588 45496
rect 38388 45450 38400 45484
rect 38576 45450 38588 45484
rect 38388 45438 38588 45450
rect 43378 45882 43578 45894
rect 43378 45848 43390 45882
rect 43566 45848 43578 45882
rect 43378 45836 43578 45848
rect 43378 45794 43578 45806
rect 43378 45760 43390 45794
rect 43566 45760 43578 45794
rect 43378 45748 43578 45760
rect 43378 45572 43578 45584
rect 43378 45538 43390 45572
rect 43566 45538 43578 45572
rect 43378 45526 43578 45538
rect 43378 45484 43578 45496
rect 43378 45450 43390 45484
rect 43566 45450 43578 45484
rect 43378 45438 43578 45450
rect 48368 45882 48568 45894
rect 48368 45848 48380 45882
rect 48556 45848 48568 45882
rect 48368 45836 48568 45848
rect 48368 45794 48568 45806
rect 48368 45760 48380 45794
rect 48556 45760 48568 45794
rect 48368 45748 48568 45760
rect 48368 45572 48568 45584
rect 48368 45538 48380 45572
rect 48556 45538 48568 45572
rect 48368 45526 48568 45538
rect 48368 45484 48568 45496
rect 48368 45450 48380 45484
rect 48556 45450 48568 45484
rect 48368 45438 48568 45450
rect 53358 45882 53558 45894
rect 53358 45848 53370 45882
rect 53546 45848 53558 45882
rect 53358 45836 53558 45848
rect 53358 45794 53558 45806
rect 53358 45760 53370 45794
rect 53546 45760 53558 45794
rect 53358 45748 53558 45760
rect 53358 45572 53558 45584
rect 53358 45538 53370 45572
rect 53546 45538 53558 45572
rect 53358 45526 53558 45538
rect 53358 45484 53558 45496
rect 53358 45450 53370 45484
rect 53546 45450 53558 45484
rect 53358 45438 53558 45450
rect 58348 45882 58548 45894
rect 58348 45848 58360 45882
rect 58536 45848 58548 45882
rect 58348 45836 58548 45848
rect 58348 45794 58548 45806
rect 58348 45760 58360 45794
rect 58536 45760 58548 45794
rect 58348 45748 58548 45760
rect 58348 45572 58548 45584
rect 58348 45538 58360 45572
rect 58536 45538 58548 45572
rect 58348 45526 58548 45538
rect 58348 45484 58548 45496
rect 58348 45450 58360 45484
rect 58536 45450 58548 45484
rect 58348 45438 58548 45450
rect 63338 45882 63538 45894
rect 63338 45848 63350 45882
rect 63526 45848 63538 45882
rect 63338 45836 63538 45848
rect 63338 45794 63538 45806
rect 63338 45760 63350 45794
rect 63526 45760 63538 45794
rect 63338 45748 63538 45760
rect 63338 45572 63538 45584
rect 63338 45538 63350 45572
rect 63526 45538 63538 45572
rect 63338 45526 63538 45538
rect 63338 45484 63538 45496
rect 63338 45450 63350 45484
rect 63526 45450 63538 45484
rect 63338 45438 63538 45450
rect 68328 45882 68528 45894
rect 68328 45848 68340 45882
rect 68516 45848 68528 45882
rect 68328 45836 68528 45848
rect 68328 45794 68528 45806
rect 68328 45760 68340 45794
rect 68516 45760 68528 45794
rect 68328 45748 68528 45760
rect 68328 45572 68528 45584
rect 68328 45538 68340 45572
rect 68516 45538 68528 45572
rect 68328 45526 68528 45538
rect 68328 45484 68528 45496
rect 68328 45450 68340 45484
rect 68516 45450 68528 45484
rect 68328 45438 68528 45450
rect 73318 45882 73518 45894
rect 73318 45848 73330 45882
rect 73506 45848 73518 45882
rect 73318 45836 73518 45848
rect 73318 45794 73518 45806
rect 73318 45760 73330 45794
rect 73506 45760 73518 45794
rect 73318 45748 73518 45760
rect 73318 45572 73518 45584
rect 73318 45538 73330 45572
rect 73506 45538 73518 45572
rect 73318 45526 73518 45538
rect 73318 45484 73518 45496
rect 73318 45450 73330 45484
rect 73506 45450 73518 45484
rect 73318 45438 73518 45450
rect 78308 45882 78508 45894
rect 78308 45848 78320 45882
rect 78496 45848 78508 45882
rect 78308 45836 78508 45848
rect 78308 45794 78508 45806
rect 78308 45760 78320 45794
rect 78496 45760 78508 45794
rect 78308 45748 78508 45760
rect 78308 45572 78508 45584
rect 78308 45538 78320 45572
rect 78496 45538 78508 45572
rect 78308 45526 78508 45538
rect 78308 45484 78508 45496
rect 78308 45450 78320 45484
rect 78496 45450 78508 45484
rect 78308 45438 78508 45450
rect 3458 44172 3658 44184
rect 3458 44138 3470 44172
rect 3646 44138 3658 44172
rect 3458 44126 3658 44138
rect 3458 44084 3658 44096
rect 3458 44050 3470 44084
rect 3646 44050 3658 44084
rect 3458 44038 3658 44050
rect 3458 43862 3658 43874
rect 3458 43828 3470 43862
rect 3646 43828 3658 43862
rect 3458 43816 3658 43828
rect 3458 43774 3658 43786
rect 3458 43740 3470 43774
rect 3646 43740 3658 43774
rect 3458 43728 3658 43740
rect 8448 44172 8648 44184
rect 8448 44138 8460 44172
rect 8636 44138 8648 44172
rect 8448 44126 8648 44138
rect 8448 44084 8648 44096
rect 8448 44050 8460 44084
rect 8636 44050 8648 44084
rect 8448 44038 8648 44050
rect 8448 43862 8648 43874
rect 8448 43828 8460 43862
rect 8636 43828 8648 43862
rect 8448 43816 8648 43828
rect 8448 43774 8648 43786
rect 8448 43740 8460 43774
rect 8636 43740 8648 43774
rect 8448 43728 8648 43740
rect 13438 44172 13638 44184
rect 13438 44138 13450 44172
rect 13626 44138 13638 44172
rect 13438 44126 13638 44138
rect 13438 44084 13638 44096
rect 13438 44050 13450 44084
rect 13626 44050 13638 44084
rect 13438 44038 13638 44050
rect 13438 43862 13638 43874
rect 13438 43828 13450 43862
rect 13626 43828 13638 43862
rect 13438 43816 13638 43828
rect 13438 43774 13638 43786
rect 13438 43740 13450 43774
rect 13626 43740 13638 43774
rect 13438 43728 13638 43740
rect 18428 44172 18628 44184
rect 18428 44138 18440 44172
rect 18616 44138 18628 44172
rect 18428 44126 18628 44138
rect 18428 44084 18628 44096
rect 18428 44050 18440 44084
rect 18616 44050 18628 44084
rect 18428 44038 18628 44050
rect 18428 43862 18628 43874
rect 18428 43828 18440 43862
rect 18616 43828 18628 43862
rect 18428 43816 18628 43828
rect 18428 43774 18628 43786
rect 18428 43740 18440 43774
rect 18616 43740 18628 43774
rect 18428 43728 18628 43740
rect 23418 44172 23618 44184
rect 23418 44138 23430 44172
rect 23606 44138 23618 44172
rect 23418 44126 23618 44138
rect 23418 44084 23618 44096
rect 23418 44050 23430 44084
rect 23606 44050 23618 44084
rect 23418 44038 23618 44050
rect 23418 43862 23618 43874
rect 23418 43828 23430 43862
rect 23606 43828 23618 43862
rect 23418 43816 23618 43828
rect 23418 43774 23618 43786
rect 23418 43740 23430 43774
rect 23606 43740 23618 43774
rect 23418 43728 23618 43740
rect 28408 44172 28608 44184
rect 28408 44138 28420 44172
rect 28596 44138 28608 44172
rect 28408 44126 28608 44138
rect 28408 44084 28608 44096
rect 28408 44050 28420 44084
rect 28596 44050 28608 44084
rect 28408 44038 28608 44050
rect 28408 43862 28608 43874
rect 28408 43828 28420 43862
rect 28596 43828 28608 43862
rect 28408 43816 28608 43828
rect 28408 43774 28608 43786
rect 28408 43740 28420 43774
rect 28596 43740 28608 43774
rect 28408 43728 28608 43740
rect 33398 44172 33598 44184
rect 33398 44138 33410 44172
rect 33586 44138 33598 44172
rect 33398 44126 33598 44138
rect 33398 44084 33598 44096
rect 33398 44050 33410 44084
rect 33586 44050 33598 44084
rect 33398 44038 33598 44050
rect 33398 43862 33598 43874
rect 33398 43828 33410 43862
rect 33586 43828 33598 43862
rect 33398 43816 33598 43828
rect 33398 43774 33598 43786
rect 33398 43740 33410 43774
rect 33586 43740 33598 43774
rect 33398 43728 33598 43740
rect 38388 44172 38588 44184
rect 38388 44138 38400 44172
rect 38576 44138 38588 44172
rect 38388 44126 38588 44138
rect 38388 44084 38588 44096
rect 38388 44050 38400 44084
rect 38576 44050 38588 44084
rect 38388 44038 38588 44050
rect 38388 43862 38588 43874
rect 38388 43828 38400 43862
rect 38576 43828 38588 43862
rect 38388 43816 38588 43828
rect 38388 43774 38588 43786
rect 38388 43740 38400 43774
rect 38576 43740 38588 43774
rect 38388 43728 38588 43740
rect 43378 44172 43578 44184
rect 43378 44138 43390 44172
rect 43566 44138 43578 44172
rect 43378 44126 43578 44138
rect 43378 44084 43578 44096
rect 43378 44050 43390 44084
rect 43566 44050 43578 44084
rect 43378 44038 43578 44050
rect 43378 43862 43578 43874
rect 43378 43828 43390 43862
rect 43566 43828 43578 43862
rect 43378 43816 43578 43828
rect 43378 43774 43578 43786
rect 43378 43740 43390 43774
rect 43566 43740 43578 43774
rect 43378 43728 43578 43740
rect 48368 44172 48568 44184
rect 48368 44138 48380 44172
rect 48556 44138 48568 44172
rect 48368 44126 48568 44138
rect 48368 44084 48568 44096
rect 48368 44050 48380 44084
rect 48556 44050 48568 44084
rect 48368 44038 48568 44050
rect 48368 43862 48568 43874
rect 48368 43828 48380 43862
rect 48556 43828 48568 43862
rect 48368 43816 48568 43828
rect 48368 43774 48568 43786
rect 48368 43740 48380 43774
rect 48556 43740 48568 43774
rect 48368 43728 48568 43740
rect 53358 44172 53558 44184
rect 53358 44138 53370 44172
rect 53546 44138 53558 44172
rect 53358 44126 53558 44138
rect 53358 44084 53558 44096
rect 53358 44050 53370 44084
rect 53546 44050 53558 44084
rect 53358 44038 53558 44050
rect 53358 43862 53558 43874
rect 53358 43828 53370 43862
rect 53546 43828 53558 43862
rect 53358 43816 53558 43828
rect 53358 43774 53558 43786
rect 53358 43740 53370 43774
rect 53546 43740 53558 43774
rect 53358 43728 53558 43740
rect 58348 44172 58548 44184
rect 58348 44138 58360 44172
rect 58536 44138 58548 44172
rect 58348 44126 58548 44138
rect 58348 44084 58548 44096
rect 58348 44050 58360 44084
rect 58536 44050 58548 44084
rect 58348 44038 58548 44050
rect 58348 43862 58548 43874
rect 58348 43828 58360 43862
rect 58536 43828 58548 43862
rect 58348 43816 58548 43828
rect 58348 43774 58548 43786
rect 58348 43740 58360 43774
rect 58536 43740 58548 43774
rect 58348 43728 58548 43740
rect 63338 44172 63538 44184
rect 63338 44138 63350 44172
rect 63526 44138 63538 44172
rect 63338 44126 63538 44138
rect 63338 44084 63538 44096
rect 63338 44050 63350 44084
rect 63526 44050 63538 44084
rect 63338 44038 63538 44050
rect 63338 43862 63538 43874
rect 63338 43828 63350 43862
rect 63526 43828 63538 43862
rect 63338 43816 63538 43828
rect 63338 43774 63538 43786
rect 63338 43740 63350 43774
rect 63526 43740 63538 43774
rect 63338 43728 63538 43740
rect 68328 44172 68528 44184
rect 68328 44138 68340 44172
rect 68516 44138 68528 44172
rect 68328 44126 68528 44138
rect 68328 44084 68528 44096
rect 68328 44050 68340 44084
rect 68516 44050 68528 44084
rect 68328 44038 68528 44050
rect 68328 43862 68528 43874
rect 68328 43828 68340 43862
rect 68516 43828 68528 43862
rect 68328 43816 68528 43828
rect 68328 43774 68528 43786
rect 68328 43740 68340 43774
rect 68516 43740 68528 43774
rect 68328 43728 68528 43740
rect 73318 44172 73518 44184
rect 73318 44138 73330 44172
rect 73506 44138 73518 44172
rect 73318 44126 73518 44138
rect 73318 44084 73518 44096
rect 73318 44050 73330 44084
rect 73506 44050 73518 44084
rect 73318 44038 73518 44050
rect 73318 43862 73518 43874
rect 73318 43828 73330 43862
rect 73506 43828 73518 43862
rect 73318 43816 73518 43828
rect 73318 43774 73518 43786
rect 73318 43740 73330 43774
rect 73506 43740 73518 43774
rect 73318 43728 73518 43740
rect 78308 44172 78508 44184
rect 78308 44138 78320 44172
rect 78496 44138 78508 44172
rect 78308 44126 78508 44138
rect 78308 44084 78508 44096
rect 78308 44050 78320 44084
rect 78496 44050 78508 44084
rect 78308 44038 78508 44050
rect 78308 43862 78508 43874
rect 78308 43828 78320 43862
rect 78496 43828 78508 43862
rect 78308 43816 78508 43828
rect 78308 43774 78508 43786
rect 78308 43740 78320 43774
rect 78496 43740 78508 43774
rect 78308 43728 78508 43740
rect 3458 42462 3658 42474
rect 3458 42428 3470 42462
rect 3646 42428 3658 42462
rect 3458 42416 3658 42428
rect 3458 42374 3658 42386
rect 3458 42340 3470 42374
rect 3646 42340 3658 42374
rect 3458 42328 3658 42340
rect 3458 42152 3658 42164
rect 3458 42118 3470 42152
rect 3646 42118 3658 42152
rect 3458 42106 3658 42118
rect 3458 42064 3658 42076
rect 3458 42030 3470 42064
rect 3646 42030 3658 42064
rect 3458 42018 3658 42030
rect 8448 42462 8648 42474
rect 8448 42428 8460 42462
rect 8636 42428 8648 42462
rect 8448 42416 8648 42428
rect 8448 42374 8648 42386
rect 8448 42340 8460 42374
rect 8636 42340 8648 42374
rect 8448 42328 8648 42340
rect 8448 42152 8648 42164
rect 8448 42118 8460 42152
rect 8636 42118 8648 42152
rect 8448 42106 8648 42118
rect 8448 42064 8648 42076
rect 8448 42030 8460 42064
rect 8636 42030 8648 42064
rect 8448 42018 8648 42030
rect 13438 42462 13638 42474
rect 13438 42428 13450 42462
rect 13626 42428 13638 42462
rect 13438 42416 13638 42428
rect 13438 42374 13638 42386
rect 13438 42340 13450 42374
rect 13626 42340 13638 42374
rect 13438 42328 13638 42340
rect 13438 42152 13638 42164
rect 13438 42118 13450 42152
rect 13626 42118 13638 42152
rect 13438 42106 13638 42118
rect 13438 42064 13638 42076
rect 13438 42030 13450 42064
rect 13626 42030 13638 42064
rect 13438 42018 13638 42030
rect 18428 42462 18628 42474
rect 18428 42428 18440 42462
rect 18616 42428 18628 42462
rect 18428 42416 18628 42428
rect 18428 42374 18628 42386
rect 18428 42340 18440 42374
rect 18616 42340 18628 42374
rect 18428 42328 18628 42340
rect 18428 42152 18628 42164
rect 18428 42118 18440 42152
rect 18616 42118 18628 42152
rect 18428 42106 18628 42118
rect 18428 42064 18628 42076
rect 18428 42030 18440 42064
rect 18616 42030 18628 42064
rect 18428 42018 18628 42030
rect 23418 42462 23618 42474
rect 23418 42428 23430 42462
rect 23606 42428 23618 42462
rect 23418 42416 23618 42428
rect 23418 42374 23618 42386
rect 23418 42340 23430 42374
rect 23606 42340 23618 42374
rect 23418 42328 23618 42340
rect 23418 42152 23618 42164
rect 23418 42118 23430 42152
rect 23606 42118 23618 42152
rect 23418 42106 23618 42118
rect 23418 42064 23618 42076
rect 23418 42030 23430 42064
rect 23606 42030 23618 42064
rect 23418 42018 23618 42030
rect 28408 42462 28608 42474
rect 28408 42428 28420 42462
rect 28596 42428 28608 42462
rect 28408 42416 28608 42428
rect 28408 42374 28608 42386
rect 28408 42340 28420 42374
rect 28596 42340 28608 42374
rect 28408 42328 28608 42340
rect 28408 42152 28608 42164
rect 28408 42118 28420 42152
rect 28596 42118 28608 42152
rect 28408 42106 28608 42118
rect 28408 42064 28608 42076
rect 28408 42030 28420 42064
rect 28596 42030 28608 42064
rect 28408 42018 28608 42030
rect 33398 42462 33598 42474
rect 33398 42428 33410 42462
rect 33586 42428 33598 42462
rect 33398 42416 33598 42428
rect 33398 42374 33598 42386
rect 33398 42340 33410 42374
rect 33586 42340 33598 42374
rect 33398 42328 33598 42340
rect 33398 42152 33598 42164
rect 33398 42118 33410 42152
rect 33586 42118 33598 42152
rect 33398 42106 33598 42118
rect 33398 42064 33598 42076
rect 33398 42030 33410 42064
rect 33586 42030 33598 42064
rect 33398 42018 33598 42030
rect 38388 42462 38588 42474
rect 38388 42428 38400 42462
rect 38576 42428 38588 42462
rect 38388 42416 38588 42428
rect 38388 42374 38588 42386
rect 38388 42340 38400 42374
rect 38576 42340 38588 42374
rect 38388 42328 38588 42340
rect 38388 42152 38588 42164
rect 38388 42118 38400 42152
rect 38576 42118 38588 42152
rect 38388 42106 38588 42118
rect 38388 42064 38588 42076
rect 38388 42030 38400 42064
rect 38576 42030 38588 42064
rect 38388 42018 38588 42030
rect 43378 42462 43578 42474
rect 43378 42428 43390 42462
rect 43566 42428 43578 42462
rect 43378 42416 43578 42428
rect 43378 42374 43578 42386
rect 43378 42340 43390 42374
rect 43566 42340 43578 42374
rect 43378 42328 43578 42340
rect 43378 42152 43578 42164
rect 43378 42118 43390 42152
rect 43566 42118 43578 42152
rect 43378 42106 43578 42118
rect 43378 42064 43578 42076
rect 43378 42030 43390 42064
rect 43566 42030 43578 42064
rect 43378 42018 43578 42030
rect 48368 42462 48568 42474
rect 48368 42428 48380 42462
rect 48556 42428 48568 42462
rect 48368 42416 48568 42428
rect 48368 42374 48568 42386
rect 48368 42340 48380 42374
rect 48556 42340 48568 42374
rect 48368 42328 48568 42340
rect 48368 42152 48568 42164
rect 48368 42118 48380 42152
rect 48556 42118 48568 42152
rect 48368 42106 48568 42118
rect 48368 42064 48568 42076
rect 48368 42030 48380 42064
rect 48556 42030 48568 42064
rect 48368 42018 48568 42030
rect 53358 42462 53558 42474
rect 53358 42428 53370 42462
rect 53546 42428 53558 42462
rect 53358 42416 53558 42428
rect 53358 42374 53558 42386
rect 53358 42340 53370 42374
rect 53546 42340 53558 42374
rect 53358 42328 53558 42340
rect 53358 42152 53558 42164
rect 53358 42118 53370 42152
rect 53546 42118 53558 42152
rect 53358 42106 53558 42118
rect 53358 42064 53558 42076
rect 53358 42030 53370 42064
rect 53546 42030 53558 42064
rect 53358 42018 53558 42030
rect 58348 42462 58548 42474
rect 58348 42428 58360 42462
rect 58536 42428 58548 42462
rect 58348 42416 58548 42428
rect 58348 42374 58548 42386
rect 58348 42340 58360 42374
rect 58536 42340 58548 42374
rect 58348 42328 58548 42340
rect 58348 42152 58548 42164
rect 58348 42118 58360 42152
rect 58536 42118 58548 42152
rect 58348 42106 58548 42118
rect 58348 42064 58548 42076
rect 58348 42030 58360 42064
rect 58536 42030 58548 42064
rect 58348 42018 58548 42030
rect 63338 42462 63538 42474
rect 63338 42428 63350 42462
rect 63526 42428 63538 42462
rect 63338 42416 63538 42428
rect 63338 42374 63538 42386
rect 63338 42340 63350 42374
rect 63526 42340 63538 42374
rect 63338 42328 63538 42340
rect 63338 42152 63538 42164
rect 63338 42118 63350 42152
rect 63526 42118 63538 42152
rect 63338 42106 63538 42118
rect 63338 42064 63538 42076
rect 63338 42030 63350 42064
rect 63526 42030 63538 42064
rect 63338 42018 63538 42030
rect 68328 42462 68528 42474
rect 68328 42428 68340 42462
rect 68516 42428 68528 42462
rect 68328 42416 68528 42428
rect 68328 42374 68528 42386
rect 68328 42340 68340 42374
rect 68516 42340 68528 42374
rect 68328 42328 68528 42340
rect 68328 42152 68528 42164
rect 68328 42118 68340 42152
rect 68516 42118 68528 42152
rect 68328 42106 68528 42118
rect 68328 42064 68528 42076
rect 68328 42030 68340 42064
rect 68516 42030 68528 42064
rect 68328 42018 68528 42030
rect 73318 42462 73518 42474
rect 73318 42428 73330 42462
rect 73506 42428 73518 42462
rect 73318 42416 73518 42428
rect 73318 42374 73518 42386
rect 73318 42340 73330 42374
rect 73506 42340 73518 42374
rect 73318 42328 73518 42340
rect 73318 42152 73518 42164
rect 73318 42118 73330 42152
rect 73506 42118 73518 42152
rect 73318 42106 73518 42118
rect 73318 42064 73518 42076
rect 73318 42030 73330 42064
rect 73506 42030 73518 42064
rect 73318 42018 73518 42030
rect 78308 42462 78508 42474
rect 78308 42428 78320 42462
rect 78496 42428 78508 42462
rect 78308 42416 78508 42428
rect 78308 42374 78508 42386
rect 78308 42340 78320 42374
rect 78496 42340 78508 42374
rect 78308 42328 78508 42340
rect 78308 42152 78508 42164
rect 78308 42118 78320 42152
rect 78496 42118 78508 42152
rect 78308 42106 78508 42118
rect 78308 42064 78508 42076
rect 78308 42030 78320 42064
rect 78496 42030 78508 42064
rect 78308 42018 78508 42030
rect 3458 40752 3658 40764
rect 3458 40718 3470 40752
rect 3646 40718 3658 40752
rect 3458 40706 3658 40718
rect 3458 40664 3658 40676
rect 3458 40630 3470 40664
rect 3646 40630 3658 40664
rect 3458 40618 3658 40630
rect 3458 40442 3658 40454
rect 3458 40408 3470 40442
rect 3646 40408 3658 40442
rect 3458 40396 3658 40408
rect 3458 40354 3658 40366
rect 3458 40320 3470 40354
rect 3646 40320 3658 40354
rect 3458 40308 3658 40320
rect 8448 40752 8648 40764
rect 8448 40718 8460 40752
rect 8636 40718 8648 40752
rect 8448 40706 8648 40718
rect 8448 40664 8648 40676
rect 8448 40630 8460 40664
rect 8636 40630 8648 40664
rect 8448 40618 8648 40630
rect 8448 40442 8648 40454
rect 8448 40408 8460 40442
rect 8636 40408 8648 40442
rect 8448 40396 8648 40408
rect 8448 40354 8648 40366
rect 8448 40320 8460 40354
rect 8636 40320 8648 40354
rect 8448 40308 8648 40320
rect 13438 40752 13638 40764
rect 13438 40718 13450 40752
rect 13626 40718 13638 40752
rect 13438 40706 13638 40718
rect 13438 40664 13638 40676
rect 13438 40630 13450 40664
rect 13626 40630 13638 40664
rect 13438 40618 13638 40630
rect 13438 40442 13638 40454
rect 13438 40408 13450 40442
rect 13626 40408 13638 40442
rect 13438 40396 13638 40408
rect 13438 40354 13638 40366
rect 13438 40320 13450 40354
rect 13626 40320 13638 40354
rect 13438 40308 13638 40320
rect 18428 40752 18628 40764
rect 18428 40718 18440 40752
rect 18616 40718 18628 40752
rect 18428 40706 18628 40718
rect 18428 40664 18628 40676
rect 18428 40630 18440 40664
rect 18616 40630 18628 40664
rect 18428 40618 18628 40630
rect 18428 40442 18628 40454
rect 18428 40408 18440 40442
rect 18616 40408 18628 40442
rect 18428 40396 18628 40408
rect 18428 40354 18628 40366
rect 18428 40320 18440 40354
rect 18616 40320 18628 40354
rect 18428 40308 18628 40320
rect 23418 40752 23618 40764
rect 23418 40718 23430 40752
rect 23606 40718 23618 40752
rect 23418 40706 23618 40718
rect 23418 40664 23618 40676
rect 23418 40630 23430 40664
rect 23606 40630 23618 40664
rect 23418 40618 23618 40630
rect 23418 40442 23618 40454
rect 23418 40408 23430 40442
rect 23606 40408 23618 40442
rect 23418 40396 23618 40408
rect 23418 40354 23618 40366
rect 23418 40320 23430 40354
rect 23606 40320 23618 40354
rect 23418 40308 23618 40320
rect 28408 40752 28608 40764
rect 28408 40718 28420 40752
rect 28596 40718 28608 40752
rect 28408 40706 28608 40718
rect 28408 40664 28608 40676
rect 28408 40630 28420 40664
rect 28596 40630 28608 40664
rect 28408 40618 28608 40630
rect 28408 40442 28608 40454
rect 28408 40408 28420 40442
rect 28596 40408 28608 40442
rect 28408 40396 28608 40408
rect 28408 40354 28608 40366
rect 28408 40320 28420 40354
rect 28596 40320 28608 40354
rect 28408 40308 28608 40320
rect 33398 40752 33598 40764
rect 33398 40718 33410 40752
rect 33586 40718 33598 40752
rect 33398 40706 33598 40718
rect 33398 40664 33598 40676
rect 33398 40630 33410 40664
rect 33586 40630 33598 40664
rect 33398 40618 33598 40630
rect 33398 40442 33598 40454
rect 33398 40408 33410 40442
rect 33586 40408 33598 40442
rect 33398 40396 33598 40408
rect 33398 40354 33598 40366
rect 33398 40320 33410 40354
rect 33586 40320 33598 40354
rect 33398 40308 33598 40320
rect 38388 40752 38588 40764
rect 38388 40718 38400 40752
rect 38576 40718 38588 40752
rect 38388 40706 38588 40718
rect 38388 40664 38588 40676
rect 38388 40630 38400 40664
rect 38576 40630 38588 40664
rect 38388 40618 38588 40630
rect 38388 40442 38588 40454
rect 38388 40408 38400 40442
rect 38576 40408 38588 40442
rect 38388 40396 38588 40408
rect 38388 40354 38588 40366
rect 38388 40320 38400 40354
rect 38576 40320 38588 40354
rect 38388 40308 38588 40320
rect 43378 40752 43578 40764
rect 43378 40718 43390 40752
rect 43566 40718 43578 40752
rect 43378 40706 43578 40718
rect 43378 40664 43578 40676
rect 43378 40630 43390 40664
rect 43566 40630 43578 40664
rect 43378 40618 43578 40630
rect 43378 40442 43578 40454
rect 43378 40408 43390 40442
rect 43566 40408 43578 40442
rect 43378 40396 43578 40408
rect 43378 40354 43578 40366
rect 43378 40320 43390 40354
rect 43566 40320 43578 40354
rect 43378 40308 43578 40320
rect 48368 40752 48568 40764
rect 48368 40718 48380 40752
rect 48556 40718 48568 40752
rect 48368 40706 48568 40718
rect 48368 40664 48568 40676
rect 48368 40630 48380 40664
rect 48556 40630 48568 40664
rect 48368 40618 48568 40630
rect 48368 40442 48568 40454
rect 48368 40408 48380 40442
rect 48556 40408 48568 40442
rect 48368 40396 48568 40408
rect 48368 40354 48568 40366
rect 48368 40320 48380 40354
rect 48556 40320 48568 40354
rect 48368 40308 48568 40320
rect 53358 40752 53558 40764
rect 53358 40718 53370 40752
rect 53546 40718 53558 40752
rect 53358 40706 53558 40718
rect 53358 40664 53558 40676
rect 53358 40630 53370 40664
rect 53546 40630 53558 40664
rect 53358 40618 53558 40630
rect 53358 40442 53558 40454
rect 53358 40408 53370 40442
rect 53546 40408 53558 40442
rect 53358 40396 53558 40408
rect 53358 40354 53558 40366
rect 53358 40320 53370 40354
rect 53546 40320 53558 40354
rect 53358 40308 53558 40320
rect 58348 40752 58548 40764
rect 58348 40718 58360 40752
rect 58536 40718 58548 40752
rect 58348 40706 58548 40718
rect 58348 40664 58548 40676
rect 58348 40630 58360 40664
rect 58536 40630 58548 40664
rect 58348 40618 58548 40630
rect 58348 40442 58548 40454
rect 58348 40408 58360 40442
rect 58536 40408 58548 40442
rect 58348 40396 58548 40408
rect 58348 40354 58548 40366
rect 58348 40320 58360 40354
rect 58536 40320 58548 40354
rect 58348 40308 58548 40320
rect 63338 40752 63538 40764
rect 63338 40718 63350 40752
rect 63526 40718 63538 40752
rect 63338 40706 63538 40718
rect 63338 40664 63538 40676
rect 63338 40630 63350 40664
rect 63526 40630 63538 40664
rect 63338 40618 63538 40630
rect 63338 40442 63538 40454
rect 63338 40408 63350 40442
rect 63526 40408 63538 40442
rect 63338 40396 63538 40408
rect 63338 40354 63538 40366
rect 63338 40320 63350 40354
rect 63526 40320 63538 40354
rect 63338 40308 63538 40320
rect 68328 40752 68528 40764
rect 68328 40718 68340 40752
rect 68516 40718 68528 40752
rect 68328 40706 68528 40718
rect 68328 40664 68528 40676
rect 68328 40630 68340 40664
rect 68516 40630 68528 40664
rect 68328 40618 68528 40630
rect 68328 40442 68528 40454
rect 68328 40408 68340 40442
rect 68516 40408 68528 40442
rect 68328 40396 68528 40408
rect 68328 40354 68528 40366
rect 68328 40320 68340 40354
rect 68516 40320 68528 40354
rect 68328 40308 68528 40320
rect 73318 40752 73518 40764
rect 73318 40718 73330 40752
rect 73506 40718 73518 40752
rect 73318 40706 73518 40718
rect 73318 40664 73518 40676
rect 73318 40630 73330 40664
rect 73506 40630 73518 40664
rect 73318 40618 73518 40630
rect 73318 40442 73518 40454
rect 73318 40408 73330 40442
rect 73506 40408 73518 40442
rect 73318 40396 73518 40408
rect 73318 40354 73518 40366
rect 73318 40320 73330 40354
rect 73506 40320 73518 40354
rect 73318 40308 73518 40320
rect 78308 40752 78508 40764
rect 78308 40718 78320 40752
rect 78496 40718 78508 40752
rect 78308 40706 78508 40718
rect 78308 40664 78508 40676
rect 78308 40630 78320 40664
rect 78496 40630 78508 40664
rect 78308 40618 78508 40630
rect 78308 40442 78508 40454
rect 78308 40408 78320 40442
rect 78496 40408 78508 40442
rect 78308 40396 78508 40408
rect 78308 40354 78508 40366
rect 78308 40320 78320 40354
rect 78496 40320 78508 40354
rect 78308 40308 78508 40320
<< ndiffc >>
rect 2972 66368 3148 66402
rect 2972 66280 3148 66314
rect 2972 66058 3148 66092
rect 2972 65970 3148 66004
rect 7962 66368 8138 66402
rect 7962 66280 8138 66314
rect 7962 66058 8138 66092
rect 7962 65970 8138 66004
rect 12952 66368 13128 66402
rect 12952 66280 13128 66314
rect 12952 66058 13128 66092
rect 12952 65970 13128 66004
rect 17942 66368 18118 66402
rect 17942 66280 18118 66314
rect 17942 66058 18118 66092
rect 17942 65970 18118 66004
rect 22932 66368 23108 66402
rect 22932 66280 23108 66314
rect 22932 66058 23108 66092
rect 22932 65970 23108 66004
rect 27922 66368 28098 66402
rect 27922 66280 28098 66314
rect 27922 66058 28098 66092
rect 27922 65970 28098 66004
rect 32912 66368 33088 66402
rect 32912 66280 33088 66314
rect 32912 66058 33088 66092
rect 32912 65970 33088 66004
rect 37902 66368 38078 66402
rect 37902 66280 38078 66314
rect 37902 66058 38078 66092
rect 37902 65970 38078 66004
rect 42892 66368 43068 66402
rect 42892 66280 43068 66314
rect 42892 66058 43068 66092
rect 42892 65970 43068 66004
rect 47882 66368 48058 66402
rect 47882 66280 48058 66314
rect 47882 66058 48058 66092
rect 47882 65970 48058 66004
rect 52872 66368 53048 66402
rect 52872 66280 53048 66314
rect 52872 66058 53048 66092
rect 52872 65970 53048 66004
rect 57862 66368 58038 66402
rect 57862 66280 58038 66314
rect 57862 66058 58038 66092
rect 57862 65970 58038 66004
rect 62852 66368 63028 66402
rect 62852 66280 63028 66314
rect 62852 66058 63028 66092
rect 62852 65970 63028 66004
rect 67842 66368 68018 66402
rect 67842 66280 68018 66314
rect 67842 66058 68018 66092
rect 67842 65970 68018 66004
rect 72832 66368 73008 66402
rect 72832 66280 73008 66314
rect 72832 66058 73008 66092
rect 72832 65970 73008 66004
rect 77822 66368 77998 66402
rect 77822 66280 77998 66314
rect 77822 66058 77998 66092
rect 77822 65970 77998 66004
rect 2972 64658 3148 64692
rect 2972 64570 3148 64604
rect 2972 64348 3148 64382
rect 2972 64260 3148 64294
rect 7962 64658 8138 64692
rect 7962 64570 8138 64604
rect 7962 64348 8138 64382
rect 7962 64260 8138 64294
rect 12952 64658 13128 64692
rect 12952 64570 13128 64604
rect 12952 64348 13128 64382
rect 12952 64260 13128 64294
rect 17942 64658 18118 64692
rect 17942 64570 18118 64604
rect 17942 64348 18118 64382
rect 17942 64260 18118 64294
rect 22932 64658 23108 64692
rect 22932 64570 23108 64604
rect 22932 64348 23108 64382
rect 22932 64260 23108 64294
rect 27922 64658 28098 64692
rect 27922 64570 28098 64604
rect 27922 64348 28098 64382
rect 27922 64260 28098 64294
rect 32912 64658 33088 64692
rect 32912 64570 33088 64604
rect 32912 64348 33088 64382
rect 32912 64260 33088 64294
rect 37902 64658 38078 64692
rect 37902 64570 38078 64604
rect 37902 64348 38078 64382
rect 37902 64260 38078 64294
rect 42892 64658 43068 64692
rect 42892 64570 43068 64604
rect 42892 64348 43068 64382
rect 42892 64260 43068 64294
rect 47882 64658 48058 64692
rect 47882 64570 48058 64604
rect 47882 64348 48058 64382
rect 47882 64260 48058 64294
rect 52872 64658 53048 64692
rect 52872 64570 53048 64604
rect 52872 64348 53048 64382
rect 52872 64260 53048 64294
rect 57862 64658 58038 64692
rect 57862 64570 58038 64604
rect 57862 64348 58038 64382
rect 57862 64260 58038 64294
rect 62852 64658 63028 64692
rect 62852 64570 63028 64604
rect 62852 64348 63028 64382
rect 62852 64260 63028 64294
rect 67842 64658 68018 64692
rect 67842 64570 68018 64604
rect 67842 64348 68018 64382
rect 67842 64260 68018 64294
rect 72832 64658 73008 64692
rect 72832 64570 73008 64604
rect 72832 64348 73008 64382
rect 72832 64260 73008 64294
rect 77822 64658 77998 64692
rect 77822 64570 77998 64604
rect 77822 64348 77998 64382
rect 77822 64260 77998 64294
rect 2972 62948 3148 62982
rect 2972 62860 3148 62894
rect 2972 62638 3148 62672
rect 2972 62550 3148 62584
rect 7962 62948 8138 62982
rect 7962 62860 8138 62894
rect 7962 62638 8138 62672
rect 7962 62550 8138 62584
rect 12952 62948 13128 62982
rect 12952 62860 13128 62894
rect 12952 62638 13128 62672
rect 12952 62550 13128 62584
rect 17942 62948 18118 62982
rect 17942 62860 18118 62894
rect 17942 62638 18118 62672
rect 17942 62550 18118 62584
rect 22932 62948 23108 62982
rect 22932 62860 23108 62894
rect 22932 62638 23108 62672
rect 22932 62550 23108 62584
rect 27922 62948 28098 62982
rect 27922 62860 28098 62894
rect 27922 62638 28098 62672
rect 27922 62550 28098 62584
rect 32912 62948 33088 62982
rect 32912 62860 33088 62894
rect 32912 62638 33088 62672
rect 32912 62550 33088 62584
rect 37902 62948 38078 62982
rect 37902 62860 38078 62894
rect 37902 62638 38078 62672
rect 37902 62550 38078 62584
rect 42892 62948 43068 62982
rect 42892 62860 43068 62894
rect 42892 62638 43068 62672
rect 42892 62550 43068 62584
rect 47882 62948 48058 62982
rect 47882 62860 48058 62894
rect 47882 62638 48058 62672
rect 47882 62550 48058 62584
rect 52872 62948 53048 62982
rect 52872 62860 53048 62894
rect 52872 62638 53048 62672
rect 52872 62550 53048 62584
rect 57862 62948 58038 62982
rect 57862 62860 58038 62894
rect 57862 62638 58038 62672
rect 57862 62550 58038 62584
rect 62852 62948 63028 62982
rect 62852 62860 63028 62894
rect 62852 62638 63028 62672
rect 62852 62550 63028 62584
rect 67842 62948 68018 62982
rect 67842 62860 68018 62894
rect 67842 62638 68018 62672
rect 67842 62550 68018 62584
rect 72832 62948 73008 62982
rect 72832 62860 73008 62894
rect 72832 62638 73008 62672
rect 72832 62550 73008 62584
rect 77822 62948 77998 62982
rect 77822 62860 77998 62894
rect 77822 62638 77998 62672
rect 77822 62550 77998 62584
rect 2972 61238 3148 61272
rect 2972 61150 3148 61184
rect 2972 60928 3148 60962
rect 2972 60840 3148 60874
rect 7962 61238 8138 61272
rect 7962 61150 8138 61184
rect 7962 60928 8138 60962
rect 7962 60840 8138 60874
rect 12952 61238 13128 61272
rect 12952 61150 13128 61184
rect 12952 60928 13128 60962
rect 12952 60840 13128 60874
rect 17942 61238 18118 61272
rect 17942 61150 18118 61184
rect 17942 60928 18118 60962
rect 17942 60840 18118 60874
rect 22932 61238 23108 61272
rect 22932 61150 23108 61184
rect 22932 60928 23108 60962
rect 22932 60840 23108 60874
rect 27922 61238 28098 61272
rect 27922 61150 28098 61184
rect 27922 60928 28098 60962
rect 27922 60840 28098 60874
rect 32912 61238 33088 61272
rect 32912 61150 33088 61184
rect 32912 60928 33088 60962
rect 32912 60840 33088 60874
rect 37902 61238 38078 61272
rect 37902 61150 38078 61184
rect 37902 60928 38078 60962
rect 37902 60840 38078 60874
rect 42892 61238 43068 61272
rect 42892 61150 43068 61184
rect 42892 60928 43068 60962
rect 42892 60840 43068 60874
rect 47882 61238 48058 61272
rect 47882 61150 48058 61184
rect 47882 60928 48058 60962
rect 47882 60840 48058 60874
rect 52872 61238 53048 61272
rect 52872 61150 53048 61184
rect 52872 60928 53048 60962
rect 52872 60840 53048 60874
rect 57862 61238 58038 61272
rect 57862 61150 58038 61184
rect 57862 60928 58038 60962
rect 57862 60840 58038 60874
rect 62852 61238 63028 61272
rect 62852 61150 63028 61184
rect 62852 60928 63028 60962
rect 62852 60840 63028 60874
rect 67842 61238 68018 61272
rect 67842 61150 68018 61184
rect 67842 60928 68018 60962
rect 67842 60840 68018 60874
rect 72832 61238 73008 61272
rect 72832 61150 73008 61184
rect 72832 60928 73008 60962
rect 72832 60840 73008 60874
rect 77822 61238 77998 61272
rect 77822 61150 77998 61184
rect 77822 60928 77998 60962
rect 77822 60840 77998 60874
rect 2972 59528 3148 59562
rect 2972 59440 3148 59474
rect 2972 59218 3148 59252
rect 2972 59130 3148 59164
rect 7962 59528 8138 59562
rect 7962 59440 8138 59474
rect 7962 59218 8138 59252
rect 7962 59130 8138 59164
rect 12952 59528 13128 59562
rect 12952 59440 13128 59474
rect 12952 59218 13128 59252
rect 12952 59130 13128 59164
rect 17942 59528 18118 59562
rect 17942 59440 18118 59474
rect 17942 59218 18118 59252
rect 17942 59130 18118 59164
rect 22932 59528 23108 59562
rect 22932 59440 23108 59474
rect 22932 59218 23108 59252
rect 22932 59130 23108 59164
rect 27922 59528 28098 59562
rect 27922 59440 28098 59474
rect 27922 59218 28098 59252
rect 27922 59130 28098 59164
rect 32912 59528 33088 59562
rect 32912 59440 33088 59474
rect 32912 59218 33088 59252
rect 32912 59130 33088 59164
rect 37902 59528 38078 59562
rect 37902 59440 38078 59474
rect 37902 59218 38078 59252
rect 37902 59130 38078 59164
rect 42892 59528 43068 59562
rect 42892 59440 43068 59474
rect 42892 59218 43068 59252
rect 42892 59130 43068 59164
rect 47882 59528 48058 59562
rect 47882 59440 48058 59474
rect 47882 59218 48058 59252
rect 47882 59130 48058 59164
rect 52872 59528 53048 59562
rect 52872 59440 53048 59474
rect 52872 59218 53048 59252
rect 52872 59130 53048 59164
rect 57862 59528 58038 59562
rect 57862 59440 58038 59474
rect 57862 59218 58038 59252
rect 57862 59130 58038 59164
rect 62852 59528 63028 59562
rect 62852 59440 63028 59474
rect 62852 59218 63028 59252
rect 62852 59130 63028 59164
rect 67842 59528 68018 59562
rect 67842 59440 68018 59474
rect 67842 59218 68018 59252
rect 67842 59130 68018 59164
rect 72832 59528 73008 59562
rect 72832 59440 73008 59474
rect 72832 59218 73008 59252
rect 72832 59130 73008 59164
rect 77822 59528 77998 59562
rect 77822 59440 77998 59474
rect 77822 59218 77998 59252
rect 77822 59130 77998 59164
rect 2972 57818 3148 57852
rect 2972 57730 3148 57764
rect 2972 57508 3148 57542
rect 2972 57420 3148 57454
rect 7962 57818 8138 57852
rect 7962 57730 8138 57764
rect 7962 57508 8138 57542
rect 7962 57420 8138 57454
rect 12952 57818 13128 57852
rect 12952 57730 13128 57764
rect 12952 57508 13128 57542
rect 12952 57420 13128 57454
rect 17942 57818 18118 57852
rect 17942 57730 18118 57764
rect 17942 57508 18118 57542
rect 17942 57420 18118 57454
rect 22932 57818 23108 57852
rect 22932 57730 23108 57764
rect 22932 57508 23108 57542
rect 22932 57420 23108 57454
rect 27922 57818 28098 57852
rect 27922 57730 28098 57764
rect 27922 57508 28098 57542
rect 27922 57420 28098 57454
rect 32912 57818 33088 57852
rect 32912 57730 33088 57764
rect 32912 57508 33088 57542
rect 32912 57420 33088 57454
rect 37902 57818 38078 57852
rect 37902 57730 38078 57764
rect 37902 57508 38078 57542
rect 37902 57420 38078 57454
rect 42892 57818 43068 57852
rect 42892 57730 43068 57764
rect 42892 57508 43068 57542
rect 42892 57420 43068 57454
rect 47882 57818 48058 57852
rect 47882 57730 48058 57764
rect 47882 57508 48058 57542
rect 47882 57420 48058 57454
rect 52872 57818 53048 57852
rect 52872 57730 53048 57764
rect 52872 57508 53048 57542
rect 52872 57420 53048 57454
rect 57862 57818 58038 57852
rect 57862 57730 58038 57764
rect 57862 57508 58038 57542
rect 57862 57420 58038 57454
rect 62852 57818 63028 57852
rect 62852 57730 63028 57764
rect 62852 57508 63028 57542
rect 62852 57420 63028 57454
rect 67842 57818 68018 57852
rect 67842 57730 68018 57764
rect 67842 57508 68018 57542
rect 67842 57420 68018 57454
rect 72832 57818 73008 57852
rect 72832 57730 73008 57764
rect 72832 57508 73008 57542
rect 72832 57420 73008 57454
rect 77822 57818 77998 57852
rect 77822 57730 77998 57764
rect 77822 57508 77998 57542
rect 77822 57420 77998 57454
rect 2972 56108 3148 56142
rect 2972 56020 3148 56054
rect 2972 55798 3148 55832
rect 2972 55710 3148 55744
rect 7962 56108 8138 56142
rect 7962 56020 8138 56054
rect 7962 55798 8138 55832
rect 7962 55710 8138 55744
rect 12952 56108 13128 56142
rect 12952 56020 13128 56054
rect 12952 55798 13128 55832
rect 12952 55710 13128 55744
rect 17942 56108 18118 56142
rect 17942 56020 18118 56054
rect 17942 55798 18118 55832
rect 17942 55710 18118 55744
rect 22932 56108 23108 56142
rect 22932 56020 23108 56054
rect 22932 55798 23108 55832
rect 22932 55710 23108 55744
rect 27922 56108 28098 56142
rect 27922 56020 28098 56054
rect 27922 55798 28098 55832
rect 27922 55710 28098 55744
rect 32912 56108 33088 56142
rect 32912 56020 33088 56054
rect 32912 55798 33088 55832
rect 32912 55710 33088 55744
rect 37902 56108 38078 56142
rect 37902 56020 38078 56054
rect 37902 55798 38078 55832
rect 37902 55710 38078 55744
rect 42892 56108 43068 56142
rect 42892 56020 43068 56054
rect 42892 55798 43068 55832
rect 42892 55710 43068 55744
rect 47882 56108 48058 56142
rect 47882 56020 48058 56054
rect 47882 55798 48058 55832
rect 47882 55710 48058 55744
rect 52872 56108 53048 56142
rect 52872 56020 53048 56054
rect 52872 55798 53048 55832
rect 52872 55710 53048 55744
rect 57862 56108 58038 56142
rect 57862 56020 58038 56054
rect 57862 55798 58038 55832
rect 57862 55710 58038 55744
rect 62852 56108 63028 56142
rect 62852 56020 63028 56054
rect 62852 55798 63028 55832
rect 62852 55710 63028 55744
rect 67842 56108 68018 56142
rect 67842 56020 68018 56054
rect 67842 55798 68018 55832
rect 67842 55710 68018 55744
rect 72832 56108 73008 56142
rect 72832 56020 73008 56054
rect 72832 55798 73008 55832
rect 72832 55710 73008 55744
rect 77822 56108 77998 56142
rect 77822 56020 77998 56054
rect 77822 55798 77998 55832
rect 77822 55710 77998 55744
rect 2972 54398 3148 54432
rect 2972 54310 3148 54344
rect 2972 54088 3148 54122
rect 2972 54000 3148 54034
rect 7962 54398 8138 54432
rect 7962 54310 8138 54344
rect 7962 54088 8138 54122
rect 7962 54000 8138 54034
rect 12952 54398 13128 54432
rect 12952 54310 13128 54344
rect 12952 54088 13128 54122
rect 12952 54000 13128 54034
rect 17942 54398 18118 54432
rect 17942 54310 18118 54344
rect 17942 54088 18118 54122
rect 17942 54000 18118 54034
rect 22932 54398 23108 54432
rect 22932 54310 23108 54344
rect 22932 54088 23108 54122
rect 22932 54000 23108 54034
rect 27922 54398 28098 54432
rect 27922 54310 28098 54344
rect 27922 54088 28098 54122
rect 27922 54000 28098 54034
rect 32912 54398 33088 54432
rect 32912 54310 33088 54344
rect 32912 54088 33088 54122
rect 32912 54000 33088 54034
rect 37902 54398 38078 54432
rect 37902 54310 38078 54344
rect 37902 54088 38078 54122
rect 37902 54000 38078 54034
rect 42892 54398 43068 54432
rect 42892 54310 43068 54344
rect 42892 54088 43068 54122
rect 42892 54000 43068 54034
rect 47882 54398 48058 54432
rect 47882 54310 48058 54344
rect 47882 54088 48058 54122
rect 47882 54000 48058 54034
rect 52872 54398 53048 54432
rect 52872 54310 53048 54344
rect 52872 54088 53048 54122
rect 52872 54000 53048 54034
rect 57862 54398 58038 54432
rect 57862 54310 58038 54344
rect 57862 54088 58038 54122
rect 57862 54000 58038 54034
rect 62852 54398 63028 54432
rect 62852 54310 63028 54344
rect 62852 54088 63028 54122
rect 62852 54000 63028 54034
rect 67842 54398 68018 54432
rect 67842 54310 68018 54344
rect 67842 54088 68018 54122
rect 67842 54000 68018 54034
rect 72832 54398 73008 54432
rect 72832 54310 73008 54344
rect 72832 54088 73008 54122
rect 72832 54000 73008 54034
rect 77822 54398 77998 54432
rect 77822 54310 77998 54344
rect 77822 54088 77998 54122
rect 77822 54000 77998 54034
rect 2972 52688 3148 52722
rect 2972 52600 3148 52634
rect 2972 52378 3148 52412
rect 2972 52290 3148 52324
rect 7962 52688 8138 52722
rect 7962 52600 8138 52634
rect 7962 52378 8138 52412
rect 7962 52290 8138 52324
rect 12952 52688 13128 52722
rect 12952 52600 13128 52634
rect 12952 52378 13128 52412
rect 12952 52290 13128 52324
rect 17942 52688 18118 52722
rect 17942 52600 18118 52634
rect 17942 52378 18118 52412
rect 17942 52290 18118 52324
rect 22932 52688 23108 52722
rect 22932 52600 23108 52634
rect 22932 52378 23108 52412
rect 22932 52290 23108 52324
rect 27922 52688 28098 52722
rect 27922 52600 28098 52634
rect 27922 52378 28098 52412
rect 27922 52290 28098 52324
rect 32912 52688 33088 52722
rect 32912 52600 33088 52634
rect 32912 52378 33088 52412
rect 32912 52290 33088 52324
rect 37902 52688 38078 52722
rect 37902 52600 38078 52634
rect 37902 52378 38078 52412
rect 37902 52290 38078 52324
rect 42892 52688 43068 52722
rect 42892 52600 43068 52634
rect 42892 52378 43068 52412
rect 42892 52290 43068 52324
rect 47882 52688 48058 52722
rect 47882 52600 48058 52634
rect 47882 52378 48058 52412
rect 47882 52290 48058 52324
rect 52872 52688 53048 52722
rect 52872 52600 53048 52634
rect 52872 52378 53048 52412
rect 52872 52290 53048 52324
rect 57862 52688 58038 52722
rect 57862 52600 58038 52634
rect 57862 52378 58038 52412
rect 57862 52290 58038 52324
rect 62852 52688 63028 52722
rect 62852 52600 63028 52634
rect 62852 52378 63028 52412
rect 62852 52290 63028 52324
rect 67842 52688 68018 52722
rect 67842 52600 68018 52634
rect 67842 52378 68018 52412
rect 67842 52290 68018 52324
rect 72832 52688 73008 52722
rect 72832 52600 73008 52634
rect 72832 52378 73008 52412
rect 72832 52290 73008 52324
rect 77822 52688 77998 52722
rect 77822 52600 77998 52634
rect 77822 52378 77998 52412
rect 77822 52290 77998 52324
rect 2972 50978 3148 51012
rect 2972 50890 3148 50924
rect 2972 50668 3148 50702
rect 2972 50580 3148 50614
rect 7962 50978 8138 51012
rect 7962 50890 8138 50924
rect 7962 50668 8138 50702
rect 7962 50580 8138 50614
rect 12952 50978 13128 51012
rect 12952 50890 13128 50924
rect 12952 50668 13128 50702
rect 12952 50580 13128 50614
rect 17942 50978 18118 51012
rect 17942 50890 18118 50924
rect 17942 50668 18118 50702
rect 17942 50580 18118 50614
rect 22932 50978 23108 51012
rect 22932 50890 23108 50924
rect 22932 50668 23108 50702
rect 22932 50580 23108 50614
rect 27922 50978 28098 51012
rect 27922 50890 28098 50924
rect 27922 50668 28098 50702
rect 27922 50580 28098 50614
rect 32912 50978 33088 51012
rect 32912 50890 33088 50924
rect 32912 50668 33088 50702
rect 32912 50580 33088 50614
rect 37902 50978 38078 51012
rect 37902 50890 38078 50924
rect 37902 50668 38078 50702
rect 37902 50580 38078 50614
rect 42892 50978 43068 51012
rect 42892 50890 43068 50924
rect 42892 50668 43068 50702
rect 42892 50580 43068 50614
rect 47882 50978 48058 51012
rect 47882 50890 48058 50924
rect 47882 50668 48058 50702
rect 47882 50580 48058 50614
rect 52872 50978 53048 51012
rect 52872 50890 53048 50924
rect 52872 50668 53048 50702
rect 52872 50580 53048 50614
rect 57862 50978 58038 51012
rect 57862 50890 58038 50924
rect 57862 50668 58038 50702
rect 57862 50580 58038 50614
rect 62852 50978 63028 51012
rect 62852 50890 63028 50924
rect 62852 50668 63028 50702
rect 62852 50580 63028 50614
rect 67842 50978 68018 51012
rect 67842 50890 68018 50924
rect 67842 50668 68018 50702
rect 67842 50580 68018 50614
rect 72832 50978 73008 51012
rect 72832 50890 73008 50924
rect 72832 50668 73008 50702
rect 72832 50580 73008 50614
rect 77822 50978 77998 51012
rect 77822 50890 77998 50924
rect 77822 50668 77998 50702
rect 77822 50580 77998 50614
rect 2972 49268 3148 49302
rect 2972 49180 3148 49214
rect 2972 48958 3148 48992
rect 2972 48870 3148 48904
rect 7962 49268 8138 49302
rect 7962 49180 8138 49214
rect 7962 48958 8138 48992
rect 7962 48870 8138 48904
rect 12952 49268 13128 49302
rect 12952 49180 13128 49214
rect 12952 48958 13128 48992
rect 12952 48870 13128 48904
rect 17942 49268 18118 49302
rect 17942 49180 18118 49214
rect 17942 48958 18118 48992
rect 17942 48870 18118 48904
rect 22932 49268 23108 49302
rect 22932 49180 23108 49214
rect 22932 48958 23108 48992
rect 22932 48870 23108 48904
rect 27922 49268 28098 49302
rect 27922 49180 28098 49214
rect 27922 48958 28098 48992
rect 27922 48870 28098 48904
rect 32912 49268 33088 49302
rect 32912 49180 33088 49214
rect 32912 48958 33088 48992
rect 32912 48870 33088 48904
rect 37902 49268 38078 49302
rect 37902 49180 38078 49214
rect 37902 48958 38078 48992
rect 37902 48870 38078 48904
rect 42892 49268 43068 49302
rect 42892 49180 43068 49214
rect 42892 48958 43068 48992
rect 42892 48870 43068 48904
rect 47882 49268 48058 49302
rect 47882 49180 48058 49214
rect 47882 48958 48058 48992
rect 47882 48870 48058 48904
rect 52872 49268 53048 49302
rect 52872 49180 53048 49214
rect 52872 48958 53048 48992
rect 52872 48870 53048 48904
rect 57862 49268 58038 49302
rect 57862 49180 58038 49214
rect 57862 48958 58038 48992
rect 57862 48870 58038 48904
rect 62852 49268 63028 49302
rect 62852 49180 63028 49214
rect 62852 48958 63028 48992
rect 62852 48870 63028 48904
rect 67842 49268 68018 49302
rect 67842 49180 68018 49214
rect 67842 48958 68018 48992
rect 67842 48870 68018 48904
rect 72832 49268 73008 49302
rect 72832 49180 73008 49214
rect 72832 48958 73008 48992
rect 72832 48870 73008 48904
rect 77822 49268 77998 49302
rect 77822 49180 77998 49214
rect 77822 48958 77998 48992
rect 77822 48870 77998 48904
rect 2972 47558 3148 47592
rect 2972 47470 3148 47504
rect 2972 47248 3148 47282
rect 2972 47160 3148 47194
rect 7962 47558 8138 47592
rect 7962 47470 8138 47504
rect 7962 47248 8138 47282
rect 7962 47160 8138 47194
rect 12952 47558 13128 47592
rect 12952 47470 13128 47504
rect 12952 47248 13128 47282
rect 12952 47160 13128 47194
rect 17942 47558 18118 47592
rect 17942 47470 18118 47504
rect 17942 47248 18118 47282
rect 17942 47160 18118 47194
rect 22932 47558 23108 47592
rect 22932 47470 23108 47504
rect 22932 47248 23108 47282
rect 22932 47160 23108 47194
rect 27922 47558 28098 47592
rect 27922 47470 28098 47504
rect 27922 47248 28098 47282
rect 27922 47160 28098 47194
rect 32912 47558 33088 47592
rect 32912 47470 33088 47504
rect 32912 47248 33088 47282
rect 32912 47160 33088 47194
rect 37902 47558 38078 47592
rect 37902 47470 38078 47504
rect 37902 47248 38078 47282
rect 37902 47160 38078 47194
rect 42892 47558 43068 47592
rect 42892 47470 43068 47504
rect 42892 47248 43068 47282
rect 42892 47160 43068 47194
rect 47882 47558 48058 47592
rect 47882 47470 48058 47504
rect 47882 47248 48058 47282
rect 47882 47160 48058 47194
rect 52872 47558 53048 47592
rect 52872 47470 53048 47504
rect 52872 47248 53048 47282
rect 52872 47160 53048 47194
rect 57862 47558 58038 47592
rect 57862 47470 58038 47504
rect 57862 47248 58038 47282
rect 57862 47160 58038 47194
rect 62852 47558 63028 47592
rect 62852 47470 63028 47504
rect 62852 47248 63028 47282
rect 62852 47160 63028 47194
rect 67842 47558 68018 47592
rect 67842 47470 68018 47504
rect 67842 47248 68018 47282
rect 67842 47160 68018 47194
rect 72832 47558 73008 47592
rect 72832 47470 73008 47504
rect 72832 47248 73008 47282
rect 72832 47160 73008 47194
rect 77822 47558 77998 47592
rect 77822 47470 77998 47504
rect 77822 47248 77998 47282
rect 77822 47160 77998 47194
rect 2972 45848 3148 45882
rect 2972 45760 3148 45794
rect 2972 45538 3148 45572
rect 2972 45450 3148 45484
rect 7962 45848 8138 45882
rect 7962 45760 8138 45794
rect 7962 45538 8138 45572
rect 7962 45450 8138 45484
rect 12952 45848 13128 45882
rect 12952 45760 13128 45794
rect 12952 45538 13128 45572
rect 12952 45450 13128 45484
rect 17942 45848 18118 45882
rect 17942 45760 18118 45794
rect 17942 45538 18118 45572
rect 17942 45450 18118 45484
rect 22932 45848 23108 45882
rect 22932 45760 23108 45794
rect 22932 45538 23108 45572
rect 22932 45450 23108 45484
rect 27922 45848 28098 45882
rect 27922 45760 28098 45794
rect 27922 45538 28098 45572
rect 27922 45450 28098 45484
rect 32912 45848 33088 45882
rect 32912 45760 33088 45794
rect 32912 45538 33088 45572
rect 32912 45450 33088 45484
rect 37902 45848 38078 45882
rect 37902 45760 38078 45794
rect 37902 45538 38078 45572
rect 37902 45450 38078 45484
rect 42892 45848 43068 45882
rect 42892 45760 43068 45794
rect 42892 45538 43068 45572
rect 42892 45450 43068 45484
rect 47882 45848 48058 45882
rect 47882 45760 48058 45794
rect 47882 45538 48058 45572
rect 47882 45450 48058 45484
rect 52872 45848 53048 45882
rect 52872 45760 53048 45794
rect 52872 45538 53048 45572
rect 52872 45450 53048 45484
rect 57862 45848 58038 45882
rect 57862 45760 58038 45794
rect 57862 45538 58038 45572
rect 57862 45450 58038 45484
rect 62852 45848 63028 45882
rect 62852 45760 63028 45794
rect 62852 45538 63028 45572
rect 62852 45450 63028 45484
rect 67842 45848 68018 45882
rect 67842 45760 68018 45794
rect 67842 45538 68018 45572
rect 67842 45450 68018 45484
rect 72832 45848 73008 45882
rect 72832 45760 73008 45794
rect 72832 45538 73008 45572
rect 72832 45450 73008 45484
rect 77822 45848 77998 45882
rect 77822 45760 77998 45794
rect 77822 45538 77998 45572
rect 77822 45450 77998 45484
rect 2972 44138 3148 44172
rect 2972 44050 3148 44084
rect 2972 43828 3148 43862
rect 2972 43740 3148 43774
rect 7962 44138 8138 44172
rect 7962 44050 8138 44084
rect 7962 43828 8138 43862
rect 7962 43740 8138 43774
rect 12952 44138 13128 44172
rect 12952 44050 13128 44084
rect 12952 43828 13128 43862
rect 12952 43740 13128 43774
rect 17942 44138 18118 44172
rect 17942 44050 18118 44084
rect 17942 43828 18118 43862
rect 17942 43740 18118 43774
rect 22932 44138 23108 44172
rect 22932 44050 23108 44084
rect 22932 43828 23108 43862
rect 22932 43740 23108 43774
rect 27922 44138 28098 44172
rect 27922 44050 28098 44084
rect 27922 43828 28098 43862
rect 27922 43740 28098 43774
rect 32912 44138 33088 44172
rect 32912 44050 33088 44084
rect 32912 43828 33088 43862
rect 32912 43740 33088 43774
rect 37902 44138 38078 44172
rect 37902 44050 38078 44084
rect 37902 43828 38078 43862
rect 37902 43740 38078 43774
rect 42892 44138 43068 44172
rect 42892 44050 43068 44084
rect 42892 43828 43068 43862
rect 42892 43740 43068 43774
rect 47882 44138 48058 44172
rect 47882 44050 48058 44084
rect 47882 43828 48058 43862
rect 47882 43740 48058 43774
rect 52872 44138 53048 44172
rect 52872 44050 53048 44084
rect 52872 43828 53048 43862
rect 52872 43740 53048 43774
rect 57862 44138 58038 44172
rect 57862 44050 58038 44084
rect 57862 43828 58038 43862
rect 57862 43740 58038 43774
rect 62852 44138 63028 44172
rect 62852 44050 63028 44084
rect 62852 43828 63028 43862
rect 62852 43740 63028 43774
rect 67842 44138 68018 44172
rect 67842 44050 68018 44084
rect 67842 43828 68018 43862
rect 67842 43740 68018 43774
rect 72832 44138 73008 44172
rect 72832 44050 73008 44084
rect 72832 43828 73008 43862
rect 72832 43740 73008 43774
rect 77822 44138 77998 44172
rect 77822 44050 77998 44084
rect 77822 43828 77998 43862
rect 77822 43740 77998 43774
rect 2972 42428 3148 42462
rect 2972 42340 3148 42374
rect 2972 42118 3148 42152
rect 2972 42030 3148 42064
rect 7962 42428 8138 42462
rect 7962 42340 8138 42374
rect 7962 42118 8138 42152
rect 7962 42030 8138 42064
rect 12952 42428 13128 42462
rect 12952 42340 13128 42374
rect 12952 42118 13128 42152
rect 12952 42030 13128 42064
rect 17942 42428 18118 42462
rect 17942 42340 18118 42374
rect 17942 42118 18118 42152
rect 17942 42030 18118 42064
rect 22932 42428 23108 42462
rect 22932 42340 23108 42374
rect 22932 42118 23108 42152
rect 22932 42030 23108 42064
rect 27922 42428 28098 42462
rect 27922 42340 28098 42374
rect 27922 42118 28098 42152
rect 27922 42030 28098 42064
rect 32912 42428 33088 42462
rect 32912 42340 33088 42374
rect 32912 42118 33088 42152
rect 32912 42030 33088 42064
rect 37902 42428 38078 42462
rect 37902 42340 38078 42374
rect 37902 42118 38078 42152
rect 37902 42030 38078 42064
rect 42892 42428 43068 42462
rect 42892 42340 43068 42374
rect 42892 42118 43068 42152
rect 42892 42030 43068 42064
rect 47882 42428 48058 42462
rect 47882 42340 48058 42374
rect 47882 42118 48058 42152
rect 47882 42030 48058 42064
rect 52872 42428 53048 42462
rect 52872 42340 53048 42374
rect 52872 42118 53048 42152
rect 52872 42030 53048 42064
rect 57862 42428 58038 42462
rect 57862 42340 58038 42374
rect 57862 42118 58038 42152
rect 57862 42030 58038 42064
rect 62852 42428 63028 42462
rect 62852 42340 63028 42374
rect 62852 42118 63028 42152
rect 62852 42030 63028 42064
rect 67842 42428 68018 42462
rect 67842 42340 68018 42374
rect 67842 42118 68018 42152
rect 67842 42030 68018 42064
rect 72832 42428 73008 42462
rect 72832 42340 73008 42374
rect 72832 42118 73008 42152
rect 72832 42030 73008 42064
rect 77822 42428 77998 42462
rect 77822 42340 77998 42374
rect 77822 42118 77998 42152
rect 77822 42030 77998 42064
rect 2972 40718 3148 40752
rect 2972 40630 3148 40664
rect 2972 40408 3148 40442
rect 2972 40320 3148 40354
rect 7962 40718 8138 40752
rect 7962 40630 8138 40664
rect 7962 40408 8138 40442
rect 7962 40320 8138 40354
rect 12952 40718 13128 40752
rect 12952 40630 13128 40664
rect 12952 40408 13128 40442
rect 12952 40320 13128 40354
rect 17942 40718 18118 40752
rect 17942 40630 18118 40664
rect 17942 40408 18118 40442
rect 17942 40320 18118 40354
rect 22932 40718 23108 40752
rect 22932 40630 23108 40664
rect 22932 40408 23108 40442
rect 22932 40320 23108 40354
rect 27922 40718 28098 40752
rect 27922 40630 28098 40664
rect 27922 40408 28098 40442
rect 27922 40320 28098 40354
rect 32912 40718 33088 40752
rect 32912 40630 33088 40664
rect 32912 40408 33088 40442
rect 32912 40320 33088 40354
rect 37902 40718 38078 40752
rect 37902 40630 38078 40664
rect 37902 40408 38078 40442
rect 37902 40320 38078 40354
rect 42892 40718 43068 40752
rect 42892 40630 43068 40664
rect 42892 40408 43068 40442
rect 42892 40320 43068 40354
rect 47882 40718 48058 40752
rect 47882 40630 48058 40664
rect 47882 40408 48058 40442
rect 47882 40320 48058 40354
rect 52872 40718 53048 40752
rect 52872 40630 53048 40664
rect 52872 40408 53048 40442
rect 52872 40320 53048 40354
rect 57862 40718 58038 40752
rect 57862 40630 58038 40664
rect 57862 40408 58038 40442
rect 57862 40320 58038 40354
rect 62852 40718 63028 40752
rect 62852 40630 63028 40664
rect 62852 40408 63028 40442
rect 62852 40320 63028 40354
rect 67842 40718 68018 40752
rect 67842 40630 68018 40664
rect 67842 40408 68018 40442
rect 67842 40320 68018 40354
rect 72832 40718 73008 40752
rect 72832 40630 73008 40664
rect 72832 40408 73008 40442
rect 72832 40320 73008 40354
rect 77822 40718 77998 40752
rect 77822 40630 77998 40664
rect 77822 40408 77998 40442
rect 77822 40320 77998 40354
<< pdiffc >>
rect 3470 66368 3646 66402
rect 3470 66280 3646 66314
rect 3470 66058 3646 66092
rect 3470 65970 3646 66004
rect 8460 66368 8636 66402
rect 8460 66280 8636 66314
rect 8460 66058 8636 66092
rect 8460 65970 8636 66004
rect 13450 66368 13626 66402
rect 13450 66280 13626 66314
rect 13450 66058 13626 66092
rect 13450 65970 13626 66004
rect 18440 66368 18616 66402
rect 18440 66280 18616 66314
rect 18440 66058 18616 66092
rect 18440 65970 18616 66004
rect 23430 66368 23606 66402
rect 23430 66280 23606 66314
rect 23430 66058 23606 66092
rect 23430 65970 23606 66004
rect 28420 66368 28596 66402
rect 28420 66280 28596 66314
rect 28420 66058 28596 66092
rect 28420 65970 28596 66004
rect 33410 66368 33586 66402
rect 33410 66280 33586 66314
rect 33410 66058 33586 66092
rect 33410 65970 33586 66004
rect 38400 66368 38576 66402
rect 38400 66280 38576 66314
rect 38400 66058 38576 66092
rect 38400 65970 38576 66004
rect 43390 66368 43566 66402
rect 43390 66280 43566 66314
rect 43390 66058 43566 66092
rect 43390 65970 43566 66004
rect 48380 66368 48556 66402
rect 48380 66280 48556 66314
rect 48380 66058 48556 66092
rect 48380 65970 48556 66004
rect 53370 66368 53546 66402
rect 53370 66280 53546 66314
rect 53370 66058 53546 66092
rect 53370 65970 53546 66004
rect 58360 66368 58536 66402
rect 58360 66280 58536 66314
rect 58360 66058 58536 66092
rect 58360 65970 58536 66004
rect 63350 66368 63526 66402
rect 63350 66280 63526 66314
rect 63350 66058 63526 66092
rect 63350 65970 63526 66004
rect 68340 66368 68516 66402
rect 68340 66280 68516 66314
rect 68340 66058 68516 66092
rect 68340 65970 68516 66004
rect 73330 66368 73506 66402
rect 73330 66280 73506 66314
rect 73330 66058 73506 66092
rect 73330 65970 73506 66004
rect 78320 66368 78496 66402
rect 78320 66280 78496 66314
rect 78320 66058 78496 66092
rect 78320 65970 78496 66004
rect 3470 64658 3646 64692
rect 3470 64570 3646 64604
rect 3470 64348 3646 64382
rect 3470 64260 3646 64294
rect 8460 64658 8636 64692
rect 8460 64570 8636 64604
rect 8460 64348 8636 64382
rect 8460 64260 8636 64294
rect 13450 64658 13626 64692
rect 13450 64570 13626 64604
rect 13450 64348 13626 64382
rect 13450 64260 13626 64294
rect 18440 64658 18616 64692
rect 18440 64570 18616 64604
rect 18440 64348 18616 64382
rect 18440 64260 18616 64294
rect 23430 64658 23606 64692
rect 23430 64570 23606 64604
rect 23430 64348 23606 64382
rect 23430 64260 23606 64294
rect 28420 64658 28596 64692
rect 28420 64570 28596 64604
rect 28420 64348 28596 64382
rect 28420 64260 28596 64294
rect 33410 64658 33586 64692
rect 33410 64570 33586 64604
rect 33410 64348 33586 64382
rect 33410 64260 33586 64294
rect 38400 64658 38576 64692
rect 38400 64570 38576 64604
rect 38400 64348 38576 64382
rect 38400 64260 38576 64294
rect 43390 64658 43566 64692
rect 43390 64570 43566 64604
rect 43390 64348 43566 64382
rect 43390 64260 43566 64294
rect 48380 64658 48556 64692
rect 48380 64570 48556 64604
rect 48380 64348 48556 64382
rect 48380 64260 48556 64294
rect 53370 64658 53546 64692
rect 53370 64570 53546 64604
rect 53370 64348 53546 64382
rect 53370 64260 53546 64294
rect 58360 64658 58536 64692
rect 58360 64570 58536 64604
rect 58360 64348 58536 64382
rect 58360 64260 58536 64294
rect 63350 64658 63526 64692
rect 63350 64570 63526 64604
rect 63350 64348 63526 64382
rect 63350 64260 63526 64294
rect 68340 64658 68516 64692
rect 68340 64570 68516 64604
rect 68340 64348 68516 64382
rect 68340 64260 68516 64294
rect 73330 64658 73506 64692
rect 73330 64570 73506 64604
rect 73330 64348 73506 64382
rect 73330 64260 73506 64294
rect 78320 64658 78496 64692
rect 78320 64570 78496 64604
rect 78320 64348 78496 64382
rect 78320 64260 78496 64294
rect 3470 62948 3646 62982
rect 3470 62860 3646 62894
rect 3470 62638 3646 62672
rect 3470 62550 3646 62584
rect 8460 62948 8636 62982
rect 8460 62860 8636 62894
rect 8460 62638 8636 62672
rect 8460 62550 8636 62584
rect 13450 62948 13626 62982
rect 13450 62860 13626 62894
rect 13450 62638 13626 62672
rect 13450 62550 13626 62584
rect 18440 62948 18616 62982
rect 18440 62860 18616 62894
rect 18440 62638 18616 62672
rect 18440 62550 18616 62584
rect 23430 62948 23606 62982
rect 23430 62860 23606 62894
rect 23430 62638 23606 62672
rect 23430 62550 23606 62584
rect 28420 62948 28596 62982
rect 28420 62860 28596 62894
rect 28420 62638 28596 62672
rect 28420 62550 28596 62584
rect 33410 62948 33586 62982
rect 33410 62860 33586 62894
rect 33410 62638 33586 62672
rect 33410 62550 33586 62584
rect 38400 62948 38576 62982
rect 38400 62860 38576 62894
rect 38400 62638 38576 62672
rect 38400 62550 38576 62584
rect 43390 62948 43566 62982
rect 43390 62860 43566 62894
rect 43390 62638 43566 62672
rect 43390 62550 43566 62584
rect 48380 62948 48556 62982
rect 48380 62860 48556 62894
rect 48380 62638 48556 62672
rect 48380 62550 48556 62584
rect 53370 62948 53546 62982
rect 53370 62860 53546 62894
rect 53370 62638 53546 62672
rect 53370 62550 53546 62584
rect 58360 62948 58536 62982
rect 58360 62860 58536 62894
rect 58360 62638 58536 62672
rect 58360 62550 58536 62584
rect 63350 62948 63526 62982
rect 63350 62860 63526 62894
rect 63350 62638 63526 62672
rect 63350 62550 63526 62584
rect 68340 62948 68516 62982
rect 68340 62860 68516 62894
rect 68340 62638 68516 62672
rect 68340 62550 68516 62584
rect 73330 62948 73506 62982
rect 73330 62860 73506 62894
rect 73330 62638 73506 62672
rect 73330 62550 73506 62584
rect 78320 62948 78496 62982
rect 78320 62860 78496 62894
rect 78320 62638 78496 62672
rect 78320 62550 78496 62584
rect 3470 61238 3646 61272
rect 3470 61150 3646 61184
rect 3470 60928 3646 60962
rect 3470 60840 3646 60874
rect 8460 61238 8636 61272
rect 8460 61150 8636 61184
rect 8460 60928 8636 60962
rect 8460 60840 8636 60874
rect 13450 61238 13626 61272
rect 13450 61150 13626 61184
rect 13450 60928 13626 60962
rect 13450 60840 13626 60874
rect 18440 61238 18616 61272
rect 18440 61150 18616 61184
rect 18440 60928 18616 60962
rect 18440 60840 18616 60874
rect 23430 61238 23606 61272
rect 23430 61150 23606 61184
rect 23430 60928 23606 60962
rect 23430 60840 23606 60874
rect 28420 61238 28596 61272
rect 28420 61150 28596 61184
rect 28420 60928 28596 60962
rect 28420 60840 28596 60874
rect 33410 61238 33586 61272
rect 33410 61150 33586 61184
rect 33410 60928 33586 60962
rect 33410 60840 33586 60874
rect 38400 61238 38576 61272
rect 38400 61150 38576 61184
rect 38400 60928 38576 60962
rect 38400 60840 38576 60874
rect 43390 61238 43566 61272
rect 43390 61150 43566 61184
rect 43390 60928 43566 60962
rect 43390 60840 43566 60874
rect 48380 61238 48556 61272
rect 48380 61150 48556 61184
rect 48380 60928 48556 60962
rect 48380 60840 48556 60874
rect 53370 61238 53546 61272
rect 53370 61150 53546 61184
rect 53370 60928 53546 60962
rect 53370 60840 53546 60874
rect 58360 61238 58536 61272
rect 58360 61150 58536 61184
rect 58360 60928 58536 60962
rect 58360 60840 58536 60874
rect 63350 61238 63526 61272
rect 63350 61150 63526 61184
rect 63350 60928 63526 60962
rect 63350 60840 63526 60874
rect 68340 61238 68516 61272
rect 68340 61150 68516 61184
rect 68340 60928 68516 60962
rect 68340 60840 68516 60874
rect 73330 61238 73506 61272
rect 73330 61150 73506 61184
rect 73330 60928 73506 60962
rect 73330 60840 73506 60874
rect 78320 61238 78496 61272
rect 78320 61150 78496 61184
rect 78320 60928 78496 60962
rect 78320 60840 78496 60874
rect 3470 59528 3646 59562
rect 3470 59440 3646 59474
rect 3470 59218 3646 59252
rect 3470 59130 3646 59164
rect 8460 59528 8636 59562
rect 8460 59440 8636 59474
rect 8460 59218 8636 59252
rect 8460 59130 8636 59164
rect 13450 59528 13626 59562
rect 13450 59440 13626 59474
rect 13450 59218 13626 59252
rect 13450 59130 13626 59164
rect 18440 59528 18616 59562
rect 18440 59440 18616 59474
rect 18440 59218 18616 59252
rect 18440 59130 18616 59164
rect 23430 59528 23606 59562
rect 23430 59440 23606 59474
rect 23430 59218 23606 59252
rect 23430 59130 23606 59164
rect 28420 59528 28596 59562
rect 28420 59440 28596 59474
rect 28420 59218 28596 59252
rect 28420 59130 28596 59164
rect 33410 59528 33586 59562
rect 33410 59440 33586 59474
rect 33410 59218 33586 59252
rect 33410 59130 33586 59164
rect 38400 59528 38576 59562
rect 38400 59440 38576 59474
rect 38400 59218 38576 59252
rect 38400 59130 38576 59164
rect 43390 59528 43566 59562
rect 43390 59440 43566 59474
rect 43390 59218 43566 59252
rect 43390 59130 43566 59164
rect 48380 59528 48556 59562
rect 48380 59440 48556 59474
rect 48380 59218 48556 59252
rect 48380 59130 48556 59164
rect 53370 59528 53546 59562
rect 53370 59440 53546 59474
rect 53370 59218 53546 59252
rect 53370 59130 53546 59164
rect 58360 59528 58536 59562
rect 58360 59440 58536 59474
rect 58360 59218 58536 59252
rect 58360 59130 58536 59164
rect 63350 59528 63526 59562
rect 63350 59440 63526 59474
rect 63350 59218 63526 59252
rect 63350 59130 63526 59164
rect 68340 59528 68516 59562
rect 68340 59440 68516 59474
rect 68340 59218 68516 59252
rect 68340 59130 68516 59164
rect 73330 59528 73506 59562
rect 73330 59440 73506 59474
rect 73330 59218 73506 59252
rect 73330 59130 73506 59164
rect 78320 59528 78496 59562
rect 78320 59440 78496 59474
rect 78320 59218 78496 59252
rect 78320 59130 78496 59164
rect 3470 57818 3646 57852
rect 3470 57730 3646 57764
rect 3470 57508 3646 57542
rect 3470 57420 3646 57454
rect 8460 57818 8636 57852
rect 8460 57730 8636 57764
rect 8460 57508 8636 57542
rect 8460 57420 8636 57454
rect 13450 57818 13626 57852
rect 13450 57730 13626 57764
rect 13450 57508 13626 57542
rect 13450 57420 13626 57454
rect 18440 57818 18616 57852
rect 18440 57730 18616 57764
rect 18440 57508 18616 57542
rect 18440 57420 18616 57454
rect 23430 57818 23606 57852
rect 23430 57730 23606 57764
rect 23430 57508 23606 57542
rect 23430 57420 23606 57454
rect 28420 57818 28596 57852
rect 28420 57730 28596 57764
rect 28420 57508 28596 57542
rect 28420 57420 28596 57454
rect 33410 57818 33586 57852
rect 33410 57730 33586 57764
rect 33410 57508 33586 57542
rect 33410 57420 33586 57454
rect 38400 57818 38576 57852
rect 38400 57730 38576 57764
rect 38400 57508 38576 57542
rect 38400 57420 38576 57454
rect 43390 57818 43566 57852
rect 43390 57730 43566 57764
rect 43390 57508 43566 57542
rect 43390 57420 43566 57454
rect 48380 57818 48556 57852
rect 48380 57730 48556 57764
rect 48380 57508 48556 57542
rect 48380 57420 48556 57454
rect 53370 57818 53546 57852
rect 53370 57730 53546 57764
rect 53370 57508 53546 57542
rect 53370 57420 53546 57454
rect 58360 57818 58536 57852
rect 58360 57730 58536 57764
rect 58360 57508 58536 57542
rect 58360 57420 58536 57454
rect 63350 57818 63526 57852
rect 63350 57730 63526 57764
rect 63350 57508 63526 57542
rect 63350 57420 63526 57454
rect 68340 57818 68516 57852
rect 68340 57730 68516 57764
rect 68340 57508 68516 57542
rect 68340 57420 68516 57454
rect 73330 57818 73506 57852
rect 73330 57730 73506 57764
rect 73330 57508 73506 57542
rect 73330 57420 73506 57454
rect 78320 57818 78496 57852
rect 78320 57730 78496 57764
rect 78320 57508 78496 57542
rect 78320 57420 78496 57454
rect 3470 56108 3646 56142
rect 3470 56020 3646 56054
rect 3470 55798 3646 55832
rect 3470 55710 3646 55744
rect 8460 56108 8636 56142
rect 8460 56020 8636 56054
rect 8460 55798 8636 55832
rect 8460 55710 8636 55744
rect 13450 56108 13626 56142
rect 13450 56020 13626 56054
rect 13450 55798 13626 55832
rect 13450 55710 13626 55744
rect 18440 56108 18616 56142
rect 18440 56020 18616 56054
rect 18440 55798 18616 55832
rect 18440 55710 18616 55744
rect 23430 56108 23606 56142
rect 23430 56020 23606 56054
rect 23430 55798 23606 55832
rect 23430 55710 23606 55744
rect 28420 56108 28596 56142
rect 28420 56020 28596 56054
rect 28420 55798 28596 55832
rect 28420 55710 28596 55744
rect 33410 56108 33586 56142
rect 33410 56020 33586 56054
rect 33410 55798 33586 55832
rect 33410 55710 33586 55744
rect 38400 56108 38576 56142
rect 38400 56020 38576 56054
rect 38400 55798 38576 55832
rect 38400 55710 38576 55744
rect 43390 56108 43566 56142
rect 43390 56020 43566 56054
rect 43390 55798 43566 55832
rect 43390 55710 43566 55744
rect 48380 56108 48556 56142
rect 48380 56020 48556 56054
rect 48380 55798 48556 55832
rect 48380 55710 48556 55744
rect 53370 56108 53546 56142
rect 53370 56020 53546 56054
rect 53370 55798 53546 55832
rect 53370 55710 53546 55744
rect 58360 56108 58536 56142
rect 58360 56020 58536 56054
rect 58360 55798 58536 55832
rect 58360 55710 58536 55744
rect 63350 56108 63526 56142
rect 63350 56020 63526 56054
rect 63350 55798 63526 55832
rect 63350 55710 63526 55744
rect 68340 56108 68516 56142
rect 68340 56020 68516 56054
rect 68340 55798 68516 55832
rect 68340 55710 68516 55744
rect 73330 56108 73506 56142
rect 73330 56020 73506 56054
rect 73330 55798 73506 55832
rect 73330 55710 73506 55744
rect 78320 56108 78496 56142
rect 78320 56020 78496 56054
rect 78320 55798 78496 55832
rect 78320 55710 78496 55744
rect 3470 54398 3646 54432
rect 3470 54310 3646 54344
rect 3470 54088 3646 54122
rect 3470 54000 3646 54034
rect 8460 54398 8636 54432
rect 8460 54310 8636 54344
rect 8460 54088 8636 54122
rect 8460 54000 8636 54034
rect 13450 54398 13626 54432
rect 13450 54310 13626 54344
rect 13450 54088 13626 54122
rect 13450 54000 13626 54034
rect 18440 54398 18616 54432
rect 18440 54310 18616 54344
rect 18440 54088 18616 54122
rect 18440 54000 18616 54034
rect 23430 54398 23606 54432
rect 23430 54310 23606 54344
rect 23430 54088 23606 54122
rect 23430 54000 23606 54034
rect 28420 54398 28596 54432
rect 28420 54310 28596 54344
rect 28420 54088 28596 54122
rect 28420 54000 28596 54034
rect 33410 54398 33586 54432
rect 33410 54310 33586 54344
rect 33410 54088 33586 54122
rect 33410 54000 33586 54034
rect 38400 54398 38576 54432
rect 38400 54310 38576 54344
rect 38400 54088 38576 54122
rect 38400 54000 38576 54034
rect 43390 54398 43566 54432
rect 43390 54310 43566 54344
rect 43390 54088 43566 54122
rect 43390 54000 43566 54034
rect 48380 54398 48556 54432
rect 48380 54310 48556 54344
rect 48380 54088 48556 54122
rect 48380 54000 48556 54034
rect 53370 54398 53546 54432
rect 53370 54310 53546 54344
rect 53370 54088 53546 54122
rect 53370 54000 53546 54034
rect 58360 54398 58536 54432
rect 58360 54310 58536 54344
rect 58360 54088 58536 54122
rect 58360 54000 58536 54034
rect 63350 54398 63526 54432
rect 63350 54310 63526 54344
rect 63350 54088 63526 54122
rect 63350 54000 63526 54034
rect 68340 54398 68516 54432
rect 68340 54310 68516 54344
rect 68340 54088 68516 54122
rect 68340 54000 68516 54034
rect 73330 54398 73506 54432
rect 73330 54310 73506 54344
rect 73330 54088 73506 54122
rect 73330 54000 73506 54034
rect 78320 54398 78496 54432
rect 78320 54310 78496 54344
rect 78320 54088 78496 54122
rect 78320 54000 78496 54034
rect 3470 52688 3646 52722
rect 3470 52600 3646 52634
rect 3470 52378 3646 52412
rect 3470 52290 3646 52324
rect 8460 52688 8636 52722
rect 8460 52600 8636 52634
rect 8460 52378 8636 52412
rect 8460 52290 8636 52324
rect 13450 52688 13626 52722
rect 13450 52600 13626 52634
rect 13450 52378 13626 52412
rect 13450 52290 13626 52324
rect 18440 52688 18616 52722
rect 18440 52600 18616 52634
rect 18440 52378 18616 52412
rect 18440 52290 18616 52324
rect 23430 52688 23606 52722
rect 23430 52600 23606 52634
rect 23430 52378 23606 52412
rect 23430 52290 23606 52324
rect 28420 52688 28596 52722
rect 28420 52600 28596 52634
rect 28420 52378 28596 52412
rect 28420 52290 28596 52324
rect 33410 52688 33586 52722
rect 33410 52600 33586 52634
rect 33410 52378 33586 52412
rect 33410 52290 33586 52324
rect 38400 52688 38576 52722
rect 38400 52600 38576 52634
rect 38400 52378 38576 52412
rect 38400 52290 38576 52324
rect 43390 52688 43566 52722
rect 43390 52600 43566 52634
rect 43390 52378 43566 52412
rect 43390 52290 43566 52324
rect 48380 52688 48556 52722
rect 48380 52600 48556 52634
rect 48380 52378 48556 52412
rect 48380 52290 48556 52324
rect 53370 52688 53546 52722
rect 53370 52600 53546 52634
rect 53370 52378 53546 52412
rect 53370 52290 53546 52324
rect 58360 52688 58536 52722
rect 58360 52600 58536 52634
rect 58360 52378 58536 52412
rect 58360 52290 58536 52324
rect 63350 52688 63526 52722
rect 63350 52600 63526 52634
rect 63350 52378 63526 52412
rect 63350 52290 63526 52324
rect 68340 52688 68516 52722
rect 68340 52600 68516 52634
rect 68340 52378 68516 52412
rect 68340 52290 68516 52324
rect 73330 52688 73506 52722
rect 73330 52600 73506 52634
rect 73330 52378 73506 52412
rect 73330 52290 73506 52324
rect 78320 52688 78496 52722
rect 78320 52600 78496 52634
rect 78320 52378 78496 52412
rect 78320 52290 78496 52324
rect 3470 50978 3646 51012
rect 3470 50890 3646 50924
rect 3470 50668 3646 50702
rect 3470 50580 3646 50614
rect 8460 50978 8636 51012
rect 8460 50890 8636 50924
rect 8460 50668 8636 50702
rect 8460 50580 8636 50614
rect 13450 50978 13626 51012
rect 13450 50890 13626 50924
rect 13450 50668 13626 50702
rect 13450 50580 13626 50614
rect 18440 50978 18616 51012
rect 18440 50890 18616 50924
rect 18440 50668 18616 50702
rect 18440 50580 18616 50614
rect 23430 50978 23606 51012
rect 23430 50890 23606 50924
rect 23430 50668 23606 50702
rect 23430 50580 23606 50614
rect 28420 50978 28596 51012
rect 28420 50890 28596 50924
rect 28420 50668 28596 50702
rect 28420 50580 28596 50614
rect 33410 50978 33586 51012
rect 33410 50890 33586 50924
rect 33410 50668 33586 50702
rect 33410 50580 33586 50614
rect 38400 50978 38576 51012
rect 38400 50890 38576 50924
rect 38400 50668 38576 50702
rect 38400 50580 38576 50614
rect 43390 50978 43566 51012
rect 43390 50890 43566 50924
rect 43390 50668 43566 50702
rect 43390 50580 43566 50614
rect 48380 50978 48556 51012
rect 48380 50890 48556 50924
rect 48380 50668 48556 50702
rect 48380 50580 48556 50614
rect 53370 50978 53546 51012
rect 53370 50890 53546 50924
rect 53370 50668 53546 50702
rect 53370 50580 53546 50614
rect 58360 50978 58536 51012
rect 58360 50890 58536 50924
rect 58360 50668 58536 50702
rect 58360 50580 58536 50614
rect 63350 50978 63526 51012
rect 63350 50890 63526 50924
rect 63350 50668 63526 50702
rect 63350 50580 63526 50614
rect 68340 50978 68516 51012
rect 68340 50890 68516 50924
rect 68340 50668 68516 50702
rect 68340 50580 68516 50614
rect 73330 50978 73506 51012
rect 73330 50890 73506 50924
rect 73330 50668 73506 50702
rect 73330 50580 73506 50614
rect 78320 50978 78496 51012
rect 78320 50890 78496 50924
rect 78320 50668 78496 50702
rect 78320 50580 78496 50614
rect 3470 49268 3646 49302
rect 3470 49180 3646 49214
rect 3470 48958 3646 48992
rect 3470 48870 3646 48904
rect 8460 49268 8636 49302
rect 8460 49180 8636 49214
rect 8460 48958 8636 48992
rect 8460 48870 8636 48904
rect 13450 49268 13626 49302
rect 13450 49180 13626 49214
rect 13450 48958 13626 48992
rect 13450 48870 13626 48904
rect 18440 49268 18616 49302
rect 18440 49180 18616 49214
rect 18440 48958 18616 48992
rect 18440 48870 18616 48904
rect 23430 49268 23606 49302
rect 23430 49180 23606 49214
rect 23430 48958 23606 48992
rect 23430 48870 23606 48904
rect 28420 49268 28596 49302
rect 28420 49180 28596 49214
rect 28420 48958 28596 48992
rect 28420 48870 28596 48904
rect 33410 49268 33586 49302
rect 33410 49180 33586 49214
rect 33410 48958 33586 48992
rect 33410 48870 33586 48904
rect 38400 49268 38576 49302
rect 38400 49180 38576 49214
rect 38400 48958 38576 48992
rect 38400 48870 38576 48904
rect 43390 49268 43566 49302
rect 43390 49180 43566 49214
rect 43390 48958 43566 48992
rect 43390 48870 43566 48904
rect 48380 49268 48556 49302
rect 48380 49180 48556 49214
rect 48380 48958 48556 48992
rect 48380 48870 48556 48904
rect 53370 49268 53546 49302
rect 53370 49180 53546 49214
rect 53370 48958 53546 48992
rect 53370 48870 53546 48904
rect 58360 49268 58536 49302
rect 58360 49180 58536 49214
rect 58360 48958 58536 48992
rect 58360 48870 58536 48904
rect 63350 49268 63526 49302
rect 63350 49180 63526 49214
rect 63350 48958 63526 48992
rect 63350 48870 63526 48904
rect 68340 49268 68516 49302
rect 68340 49180 68516 49214
rect 68340 48958 68516 48992
rect 68340 48870 68516 48904
rect 73330 49268 73506 49302
rect 73330 49180 73506 49214
rect 73330 48958 73506 48992
rect 73330 48870 73506 48904
rect 78320 49268 78496 49302
rect 78320 49180 78496 49214
rect 78320 48958 78496 48992
rect 78320 48870 78496 48904
rect 3470 47558 3646 47592
rect 3470 47470 3646 47504
rect 3470 47248 3646 47282
rect 3470 47160 3646 47194
rect 8460 47558 8636 47592
rect 8460 47470 8636 47504
rect 8460 47248 8636 47282
rect 8460 47160 8636 47194
rect 13450 47558 13626 47592
rect 13450 47470 13626 47504
rect 13450 47248 13626 47282
rect 13450 47160 13626 47194
rect 18440 47558 18616 47592
rect 18440 47470 18616 47504
rect 18440 47248 18616 47282
rect 18440 47160 18616 47194
rect 23430 47558 23606 47592
rect 23430 47470 23606 47504
rect 23430 47248 23606 47282
rect 23430 47160 23606 47194
rect 28420 47558 28596 47592
rect 28420 47470 28596 47504
rect 28420 47248 28596 47282
rect 28420 47160 28596 47194
rect 33410 47558 33586 47592
rect 33410 47470 33586 47504
rect 33410 47248 33586 47282
rect 33410 47160 33586 47194
rect 38400 47558 38576 47592
rect 38400 47470 38576 47504
rect 38400 47248 38576 47282
rect 38400 47160 38576 47194
rect 43390 47558 43566 47592
rect 43390 47470 43566 47504
rect 43390 47248 43566 47282
rect 43390 47160 43566 47194
rect 48380 47558 48556 47592
rect 48380 47470 48556 47504
rect 48380 47248 48556 47282
rect 48380 47160 48556 47194
rect 53370 47558 53546 47592
rect 53370 47470 53546 47504
rect 53370 47248 53546 47282
rect 53370 47160 53546 47194
rect 58360 47558 58536 47592
rect 58360 47470 58536 47504
rect 58360 47248 58536 47282
rect 58360 47160 58536 47194
rect 63350 47558 63526 47592
rect 63350 47470 63526 47504
rect 63350 47248 63526 47282
rect 63350 47160 63526 47194
rect 68340 47558 68516 47592
rect 68340 47470 68516 47504
rect 68340 47248 68516 47282
rect 68340 47160 68516 47194
rect 73330 47558 73506 47592
rect 73330 47470 73506 47504
rect 73330 47248 73506 47282
rect 73330 47160 73506 47194
rect 78320 47558 78496 47592
rect 78320 47470 78496 47504
rect 78320 47248 78496 47282
rect 78320 47160 78496 47194
rect 3470 45848 3646 45882
rect 3470 45760 3646 45794
rect 3470 45538 3646 45572
rect 3470 45450 3646 45484
rect 8460 45848 8636 45882
rect 8460 45760 8636 45794
rect 8460 45538 8636 45572
rect 8460 45450 8636 45484
rect 13450 45848 13626 45882
rect 13450 45760 13626 45794
rect 13450 45538 13626 45572
rect 13450 45450 13626 45484
rect 18440 45848 18616 45882
rect 18440 45760 18616 45794
rect 18440 45538 18616 45572
rect 18440 45450 18616 45484
rect 23430 45848 23606 45882
rect 23430 45760 23606 45794
rect 23430 45538 23606 45572
rect 23430 45450 23606 45484
rect 28420 45848 28596 45882
rect 28420 45760 28596 45794
rect 28420 45538 28596 45572
rect 28420 45450 28596 45484
rect 33410 45848 33586 45882
rect 33410 45760 33586 45794
rect 33410 45538 33586 45572
rect 33410 45450 33586 45484
rect 38400 45848 38576 45882
rect 38400 45760 38576 45794
rect 38400 45538 38576 45572
rect 38400 45450 38576 45484
rect 43390 45848 43566 45882
rect 43390 45760 43566 45794
rect 43390 45538 43566 45572
rect 43390 45450 43566 45484
rect 48380 45848 48556 45882
rect 48380 45760 48556 45794
rect 48380 45538 48556 45572
rect 48380 45450 48556 45484
rect 53370 45848 53546 45882
rect 53370 45760 53546 45794
rect 53370 45538 53546 45572
rect 53370 45450 53546 45484
rect 58360 45848 58536 45882
rect 58360 45760 58536 45794
rect 58360 45538 58536 45572
rect 58360 45450 58536 45484
rect 63350 45848 63526 45882
rect 63350 45760 63526 45794
rect 63350 45538 63526 45572
rect 63350 45450 63526 45484
rect 68340 45848 68516 45882
rect 68340 45760 68516 45794
rect 68340 45538 68516 45572
rect 68340 45450 68516 45484
rect 73330 45848 73506 45882
rect 73330 45760 73506 45794
rect 73330 45538 73506 45572
rect 73330 45450 73506 45484
rect 78320 45848 78496 45882
rect 78320 45760 78496 45794
rect 78320 45538 78496 45572
rect 78320 45450 78496 45484
rect 3470 44138 3646 44172
rect 3470 44050 3646 44084
rect 3470 43828 3646 43862
rect 3470 43740 3646 43774
rect 8460 44138 8636 44172
rect 8460 44050 8636 44084
rect 8460 43828 8636 43862
rect 8460 43740 8636 43774
rect 13450 44138 13626 44172
rect 13450 44050 13626 44084
rect 13450 43828 13626 43862
rect 13450 43740 13626 43774
rect 18440 44138 18616 44172
rect 18440 44050 18616 44084
rect 18440 43828 18616 43862
rect 18440 43740 18616 43774
rect 23430 44138 23606 44172
rect 23430 44050 23606 44084
rect 23430 43828 23606 43862
rect 23430 43740 23606 43774
rect 28420 44138 28596 44172
rect 28420 44050 28596 44084
rect 28420 43828 28596 43862
rect 28420 43740 28596 43774
rect 33410 44138 33586 44172
rect 33410 44050 33586 44084
rect 33410 43828 33586 43862
rect 33410 43740 33586 43774
rect 38400 44138 38576 44172
rect 38400 44050 38576 44084
rect 38400 43828 38576 43862
rect 38400 43740 38576 43774
rect 43390 44138 43566 44172
rect 43390 44050 43566 44084
rect 43390 43828 43566 43862
rect 43390 43740 43566 43774
rect 48380 44138 48556 44172
rect 48380 44050 48556 44084
rect 48380 43828 48556 43862
rect 48380 43740 48556 43774
rect 53370 44138 53546 44172
rect 53370 44050 53546 44084
rect 53370 43828 53546 43862
rect 53370 43740 53546 43774
rect 58360 44138 58536 44172
rect 58360 44050 58536 44084
rect 58360 43828 58536 43862
rect 58360 43740 58536 43774
rect 63350 44138 63526 44172
rect 63350 44050 63526 44084
rect 63350 43828 63526 43862
rect 63350 43740 63526 43774
rect 68340 44138 68516 44172
rect 68340 44050 68516 44084
rect 68340 43828 68516 43862
rect 68340 43740 68516 43774
rect 73330 44138 73506 44172
rect 73330 44050 73506 44084
rect 73330 43828 73506 43862
rect 73330 43740 73506 43774
rect 78320 44138 78496 44172
rect 78320 44050 78496 44084
rect 78320 43828 78496 43862
rect 78320 43740 78496 43774
rect 3470 42428 3646 42462
rect 3470 42340 3646 42374
rect 3470 42118 3646 42152
rect 3470 42030 3646 42064
rect 8460 42428 8636 42462
rect 8460 42340 8636 42374
rect 8460 42118 8636 42152
rect 8460 42030 8636 42064
rect 13450 42428 13626 42462
rect 13450 42340 13626 42374
rect 13450 42118 13626 42152
rect 13450 42030 13626 42064
rect 18440 42428 18616 42462
rect 18440 42340 18616 42374
rect 18440 42118 18616 42152
rect 18440 42030 18616 42064
rect 23430 42428 23606 42462
rect 23430 42340 23606 42374
rect 23430 42118 23606 42152
rect 23430 42030 23606 42064
rect 28420 42428 28596 42462
rect 28420 42340 28596 42374
rect 28420 42118 28596 42152
rect 28420 42030 28596 42064
rect 33410 42428 33586 42462
rect 33410 42340 33586 42374
rect 33410 42118 33586 42152
rect 33410 42030 33586 42064
rect 38400 42428 38576 42462
rect 38400 42340 38576 42374
rect 38400 42118 38576 42152
rect 38400 42030 38576 42064
rect 43390 42428 43566 42462
rect 43390 42340 43566 42374
rect 43390 42118 43566 42152
rect 43390 42030 43566 42064
rect 48380 42428 48556 42462
rect 48380 42340 48556 42374
rect 48380 42118 48556 42152
rect 48380 42030 48556 42064
rect 53370 42428 53546 42462
rect 53370 42340 53546 42374
rect 53370 42118 53546 42152
rect 53370 42030 53546 42064
rect 58360 42428 58536 42462
rect 58360 42340 58536 42374
rect 58360 42118 58536 42152
rect 58360 42030 58536 42064
rect 63350 42428 63526 42462
rect 63350 42340 63526 42374
rect 63350 42118 63526 42152
rect 63350 42030 63526 42064
rect 68340 42428 68516 42462
rect 68340 42340 68516 42374
rect 68340 42118 68516 42152
rect 68340 42030 68516 42064
rect 73330 42428 73506 42462
rect 73330 42340 73506 42374
rect 73330 42118 73506 42152
rect 73330 42030 73506 42064
rect 78320 42428 78496 42462
rect 78320 42340 78496 42374
rect 78320 42118 78496 42152
rect 78320 42030 78496 42064
rect 3470 40718 3646 40752
rect 3470 40630 3646 40664
rect 3470 40408 3646 40442
rect 3470 40320 3646 40354
rect 8460 40718 8636 40752
rect 8460 40630 8636 40664
rect 8460 40408 8636 40442
rect 8460 40320 8636 40354
rect 13450 40718 13626 40752
rect 13450 40630 13626 40664
rect 13450 40408 13626 40442
rect 13450 40320 13626 40354
rect 18440 40718 18616 40752
rect 18440 40630 18616 40664
rect 18440 40408 18616 40442
rect 18440 40320 18616 40354
rect 23430 40718 23606 40752
rect 23430 40630 23606 40664
rect 23430 40408 23606 40442
rect 23430 40320 23606 40354
rect 28420 40718 28596 40752
rect 28420 40630 28596 40664
rect 28420 40408 28596 40442
rect 28420 40320 28596 40354
rect 33410 40718 33586 40752
rect 33410 40630 33586 40664
rect 33410 40408 33586 40442
rect 33410 40320 33586 40354
rect 38400 40718 38576 40752
rect 38400 40630 38576 40664
rect 38400 40408 38576 40442
rect 38400 40320 38576 40354
rect 43390 40718 43566 40752
rect 43390 40630 43566 40664
rect 43390 40408 43566 40442
rect 43390 40320 43566 40354
rect 48380 40718 48556 40752
rect 48380 40630 48556 40664
rect 48380 40408 48556 40442
rect 48380 40320 48556 40354
rect 53370 40718 53546 40752
rect 53370 40630 53546 40664
rect 53370 40408 53546 40442
rect 53370 40320 53546 40354
rect 58360 40718 58536 40752
rect 58360 40630 58536 40664
rect 58360 40408 58536 40442
rect 58360 40320 58536 40354
rect 63350 40718 63526 40752
rect 63350 40630 63526 40664
rect 63350 40408 63526 40442
rect 63350 40320 63526 40354
rect 68340 40718 68516 40752
rect 68340 40630 68516 40664
rect 68340 40408 68516 40442
rect 68340 40320 68516 40354
rect 73330 40718 73506 40752
rect 73330 40630 73506 40664
rect 73330 40408 73506 40442
rect 73330 40320 73506 40354
rect 78320 40718 78496 40752
rect 78320 40630 78496 40664
rect 78320 40408 78496 40442
rect 78320 40320 78496 40354
<< psubdiff >>
rect 2786 66482 3272 66516
rect 2786 66420 2820 66482
rect 2786 66206 2820 66262
rect 3238 66206 3272 66482
rect 2786 66166 3272 66206
rect 2786 66110 2820 66166
rect 2786 65890 2820 65952
rect 3238 65890 3272 66166
rect 2786 65856 3272 65890
rect 7776 66482 8262 66516
rect 7776 66420 7810 66482
rect 7776 66206 7810 66262
rect 8228 66206 8262 66482
rect 7776 66166 8262 66206
rect 7776 66110 7810 66166
rect 7776 65890 7810 65952
rect 8228 65890 8262 66166
rect 7776 65856 8262 65890
rect 12766 66482 13252 66516
rect 12766 66420 12800 66482
rect 12766 66206 12800 66262
rect 13218 66206 13252 66482
rect 12766 66166 13252 66206
rect 12766 66110 12800 66166
rect 12766 65890 12800 65952
rect 13218 65890 13252 66166
rect 12766 65856 13252 65890
rect 17756 66482 18242 66516
rect 17756 66420 17790 66482
rect 17756 66206 17790 66262
rect 18208 66206 18242 66482
rect 17756 66166 18242 66206
rect 17756 66110 17790 66166
rect 17756 65890 17790 65952
rect 18208 65890 18242 66166
rect 17756 65856 18242 65890
rect 22746 66482 23232 66516
rect 22746 66420 22780 66482
rect 22746 66206 22780 66262
rect 23198 66206 23232 66482
rect 22746 66166 23232 66206
rect 22746 66110 22780 66166
rect 22746 65890 22780 65952
rect 23198 65890 23232 66166
rect 22746 65856 23232 65890
rect 27736 66482 28222 66516
rect 27736 66420 27770 66482
rect 27736 66206 27770 66262
rect 28188 66206 28222 66482
rect 27736 66166 28222 66206
rect 27736 66110 27770 66166
rect 27736 65890 27770 65952
rect 28188 65890 28222 66166
rect 27736 65856 28222 65890
rect 32726 66482 33212 66516
rect 32726 66420 32760 66482
rect 32726 66206 32760 66262
rect 33178 66206 33212 66482
rect 32726 66166 33212 66206
rect 32726 66110 32760 66166
rect 32726 65890 32760 65952
rect 33178 65890 33212 66166
rect 32726 65856 33212 65890
rect 37716 66482 38202 66516
rect 37716 66420 37750 66482
rect 37716 66206 37750 66262
rect 38168 66206 38202 66482
rect 37716 66166 38202 66206
rect 37716 66110 37750 66166
rect 37716 65890 37750 65952
rect 38168 65890 38202 66166
rect 37716 65856 38202 65890
rect 42706 66482 43192 66516
rect 42706 66420 42740 66482
rect 42706 66206 42740 66262
rect 43158 66206 43192 66482
rect 42706 66166 43192 66206
rect 42706 66110 42740 66166
rect 42706 65890 42740 65952
rect 43158 65890 43192 66166
rect 42706 65856 43192 65890
rect 47696 66482 48182 66516
rect 47696 66420 47730 66482
rect 47696 66206 47730 66262
rect 48148 66206 48182 66482
rect 47696 66166 48182 66206
rect 47696 66110 47730 66166
rect 47696 65890 47730 65952
rect 48148 65890 48182 66166
rect 47696 65856 48182 65890
rect 52686 66482 53172 66516
rect 52686 66420 52720 66482
rect 52686 66206 52720 66262
rect 53138 66206 53172 66482
rect 52686 66166 53172 66206
rect 52686 66110 52720 66166
rect 52686 65890 52720 65952
rect 53138 65890 53172 66166
rect 52686 65856 53172 65890
rect 57676 66482 58162 66516
rect 57676 66420 57710 66482
rect 57676 66206 57710 66262
rect 58128 66206 58162 66482
rect 57676 66166 58162 66206
rect 57676 66110 57710 66166
rect 57676 65890 57710 65952
rect 58128 65890 58162 66166
rect 57676 65856 58162 65890
rect 62666 66482 63152 66516
rect 62666 66420 62700 66482
rect 62666 66206 62700 66262
rect 63118 66206 63152 66482
rect 62666 66166 63152 66206
rect 62666 66110 62700 66166
rect 62666 65890 62700 65952
rect 63118 65890 63152 66166
rect 62666 65856 63152 65890
rect 67656 66482 68142 66516
rect 67656 66420 67690 66482
rect 67656 66206 67690 66262
rect 68108 66206 68142 66482
rect 67656 66166 68142 66206
rect 67656 66110 67690 66166
rect 67656 65890 67690 65952
rect 68108 65890 68142 66166
rect 67656 65856 68142 65890
rect 72646 66482 73132 66516
rect 72646 66420 72680 66482
rect 72646 66206 72680 66262
rect 73098 66206 73132 66482
rect 72646 66166 73132 66206
rect 72646 66110 72680 66166
rect 72646 65890 72680 65952
rect 73098 65890 73132 66166
rect 72646 65856 73132 65890
rect 77636 66482 78122 66516
rect 77636 66420 77670 66482
rect 77636 66206 77670 66262
rect 78088 66206 78122 66482
rect 77636 66166 78122 66206
rect 77636 66110 77670 66166
rect 77636 65890 77670 65952
rect 78088 65890 78122 66166
rect 77636 65856 78122 65890
rect 2786 64772 3272 64806
rect 2786 64710 2820 64772
rect 2786 64496 2820 64552
rect 3238 64496 3272 64772
rect 2786 64456 3272 64496
rect 2786 64400 2820 64456
rect 2786 64180 2820 64242
rect 3238 64180 3272 64456
rect 2786 64146 3272 64180
rect 7776 64772 8262 64806
rect 7776 64710 7810 64772
rect 7776 64496 7810 64552
rect 8228 64496 8262 64772
rect 7776 64456 8262 64496
rect 7776 64400 7810 64456
rect 7776 64180 7810 64242
rect 8228 64180 8262 64456
rect 7776 64146 8262 64180
rect 12766 64772 13252 64806
rect 12766 64710 12800 64772
rect 12766 64496 12800 64552
rect 13218 64496 13252 64772
rect 12766 64456 13252 64496
rect 12766 64400 12800 64456
rect 12766 64180 12800 64242
rect 13218 64180 13252 64456
rect 12766 64146 13252 64180
rect 17756 64772 18242 64806
rect 17756 64710 17790 64772
rect 17756 64496 17790 64552
rect 18208 64496 18242 64772
rect 17756 64456 18242 64496
rect 17756 64400 17790 64456
rect 17756 64180 17790 64242
rect 18208 64180 18242 64456
rect 17756 64146 18242 64180
rect 22746 64772 23232 64806
rect 22746 64710 22780 64772
rect 22746 64496 22780 64552
rect 23198 64496 23232 64772
rect 22746 64456 23232 64496
rect 22746 64400 22780 64456
rect 22746 64180 22780 64242
rect 23198 64180 23232 64456
rect 22746 64146 23232 64180
rect 27736 64772 28222 64806
rect 27736 64710 27770 64772
rect 27736 64496 27770 64552
rect 28188 64496 28222 64772
rect 27736 64456 28222 64496
rect 27736 64400 27770 64456
rect 27736 64180 27770 64242
rect 28188 64180 28222 64456
rect 27736 64146 28222 64180
rect 32726 64772 33212 64806
rect 32726 64710 32760 64772
rect 32726 64496 32760 64552
rect 33178 64496 33212 64772
rect 32726 64456 33212 64496
rect 32726 64400 32760 64456
rect 32726 64180 32760 64242
rect 33178 64180 33212 64456
rect 32726 64146 33212 64180
rect 37716 64772 38202 64806
rect 37716 64710 37750 64772
rect 37716 64496 37750 64552
rect 38168 64496 38202 64772
rect 37716 64456 38202 64496
rect 37716 64400 37750 64456
rect 37716 64180 37750 64242
rect 38168 64180 38202 64456
rect 37716 64146 38202 64180
rect 42706 64772 43192 64806
rect 42706 64710 42740 64772
rect 42706 64496 42740 64552
rect 43158 64496 43192 64772
rect 42706 64456 43192 64496
rect 42706 64400 42740 64456
rect 42706 64180 42740 64242
rect 43158 64180 43192 64456
rect 42706 64146 43192 64180
rect 47696 64772 48182 64806
rect 47696 64710 47730 64772
rect 47696 64496 47730 64552
rect 48148 64496 48182 64772
rect 47696 64456 48182 64496
rect 47696 64400 47730 64456
rect 47696 64180 47730 64242
rect 48148 64180 48182 64456
rect 47696 64146 48182 64180
rect 52686 64772 53172 64806
rect 52686 64710 52720 64772
rect 52686 64496 52720 64552
rect 53138 64496 53172 64772
rect 52686 64456 53172 64496
rect 52686 64400 52720 64456
rect 52686 64180 52720 64242
rect 53138 64180 53172 64456
rect 52686 64146 53172 64180
rect 57676 64772 58162 64806
rect 57676 64710 57710 64772
rect 57676 64496 57710 64552
rect 58128 64496 58162 64772
rect 57676 64456 58162 64496
rect 57676 64400 57710 64456
rect 57676 64180 57710 64242
rect 58128 64180 58162 64456
rect 57676 64146 58162 64180
rect 62666 64772 63152 64806
rect 62666 64710 62700 64772
rect 62666 64496 62700 64552
rect 63118 64496 63152 64772
rect 62666 64456 63152 64496
rect 62666 64400 62700 64456
rect 62666 64180 62700 64242
rect 63118 64180 63152 64456
rect 62666 64146 63152 64180
rect 67656 64772 68142 64806
rect 67656 64710 67690 64772
rect 67656 64496 67690 64552
rect 68108 64496 68142 64772
rect 67656 64456 68142 64496
rect 67656 64400 67690 64456
rect 67656 64180 67690 64242
rect 68108 64180 68142 64456
rect 67656 64146 68142 64180
rect 72646 64772 73132 64806
rect 72646 64710 72680 64772
rect 72646 64496 72680 64552
rect 73098 64496 73132 64772
rect 72646 64456 73132 64496
rect 72646 64400 72680 64456
rect 72646 64180 72680 64242
rect 73098 64180 73132 64456
rect 72646 64146 73132 64180
rect 77636 64772 78122 64806
rect 77636 64710 77670 64772
rect 77636 64496 77670 64552
rect 78088 64496 78122 64772
rect 77636 64456 78122 64496
rect 77636 64400 77670 64456
rect 77636 64180 77670 64242
rect 78088 64180 78122 64456
rect 77636 64146 78122 64180
rect 2786 63062 3272 63096
rect 2786 63000 2820 63062
rect 2786 62786 2820 62842
rect 3238 62786 3272 63062
rect 2786 62746 3272 62786
rect 2786 62690 2820 62746
rect 2786 62470 2820 62532
rect 3238 62470 3272 62746
rect 2786 62436 3272 62470
rect 7776 63062 8262 63096
rect 7776 63000 7810 63062
rect 7776 62786 7810 62842
rect 8228 62786 8262 63062
rect 7776 62746 8262 62786
rect 7776 62690 7810 62746
rect 7776 62470 7810 62532
rect 8228 62470 8262 62746
rect 7776 62436 8262 62470
rect 12766 63062 13252 63096
rect 12766 63000 12800 63062
rect 12766 62786 12800 62842
rect 13218 62786 13252 63062
rect 12766 62746 13252 62786
rect 12766 62690 12800 62746
rect 12766 62470 12800 62532
rect 13218 62470 13252 62746
rect 12766 62436 13252 62470
rect 17756 63062 18242 63096
rect 17756 63000 17790 63062
rect 17756 62786 17790 62842
rect 18208 62786 18242 63062
rect 17756 62746 18242 62786
rect 17756 62690 17790 62746
rect 17756 62470 17790 62532
rect 18208 62470 18242 62746
rect 17756 62436 18242 62470
rect 22746 63062 23232 63096
rect 22746 63000 22780 63062
rect 22746 62786 22780 62842
rect 23198 62786 23232 63062
rect 22746 62746 23232 62786
rect 22746 62690 22780 62746
rect 22746 62470 22780 62532
rect 23198 62470 23232 62746
rect 22746 62436 23232 62470
rect 27736 63062 28222 63096
rect 27736 63000 27770 63062
rect 27736 62786 27770 62842
rect 28188 62786 28222 63062
rect 27736 62746 28222 62786
rect 27736 62690 27770 62746
rect 27736 62470 27770 62532
rect 28188 62470 28222 62746
rect 27736 62436 28222 62470
rect 32726 63062 33212 63096
rect 32726 63000 32760 63062
rect 32726 62786 32760 62842
rect 33178 62786 33212 63062
rect 32726 62746 33212 62786
rect 32726 62690 32760 62746
rect 32726 62470 32760 62532
rect 33178 62470 33212 62746
rect 32726 62436 33212 62470
rect 37716 63062 38202 63096
rect 37716 63000 37750 63062
rect 37716 62786 37750 62842
rect 38168 62786 38202 63062
rect 37716 62746 38202 62786
rect 37716 62690 37750 62746
rect 37716 62470 37750 62532
rect 38168 62470 38202 62746
rect 37716 62436 38202 62470
rect 42706 63062 43192 63096
rect 42706 63000 42740 63062
rect 42706 62786 42740 62842
rect 43158 62786 43192 63062
rect 42706 62746 43192 62786
rect 42706 62690 42740 62746
rect 42706 62470 42740 62532
rect 43158 62470 43192 62746
rect 42706 62436 43192 62470
rect 47696 63062 48182 63096
rect 47696 63000 47730 63062
rect 47696 62786 47730 62842
rect 48148 62786 48182 63062
rect 47696 62746 48182 62786
rect 47696 62690 47730 62746
rect 47696 62470 47730 62532
rect 48148 62470 48182 62746
rect 47696 62436 48182 62470
rect 52686 63062 53172 63096
rect 52686 63000 52720 63062
rect 52686 62786 52720 62842
rect 53138 62786 53172 63062
rect 52686 62746 53172 62786
rect 52686 62690 52720 62746
rect 52686 62470 52720 62532
rect 53138 62470 53172 62746
rect 52686 62436 53172 62470
rect 57676 63062 58162 63096
rect 57676 63000 57710 63062
rect 57676 62786 57710 62842
rect 58128 62786 58162 63062
rect 57676 62746 58162 62786
rect 57676 62690 57710 62746
rect 57676 62470 57710 62532
rect 58128 62470 58162 62746
rect 57676 62436 58162 62470
rect 62666 63062 63152 63096
rect 62666 63000 62700 63062
rect 62666 62786 62700 62842
rect 63118 62786 63152 63062
rect 62666 62746 63152 62786
rect 62666 62690 62700 62746
rect 62666 62470 62700 62532
rect 63118 62470 63152 62746
rect 62666 62436 63152 62470
rect 67656 63062 68142 63096
rect 67656 63000 67690 63062
rect 67656 62786 67690 62842
rect 68108 62786 68142 63062
rect 67656 62746 68142 62786
rect 67656 62690 67690 62746
rect 67656 62470 67690 62532
rect 68108 62470 68142 62746
rect 67656 62436 68142 62470
rect 72646 63062 73132 63096
rect 72646 63000 72680 63062
rect 72646 62786 72680 62842
rect 73098 62786 73132 63062
rect 72646 62746 73132 62786
rect 72646 62690 72680 62746
rect 72646 62470 72680 62532
rect 73098 62470 73132 62746
rect 72646 62436 73132 62470
rect 77636 63062 78122 63096
rect 77636 63000 77670 63062
rect 77636 62786 77670 62842
rect 78088 62786 78122 63062
rect 77636 62746 78122 62786
rect 77636 62690 77670 62746
rect 77636 62470 77670 62532
rect 78088 62470 78122 62746
rect 77636 62436 78122 62470
rect 2786 61352 3272 61386
rect 2786 61290 2820 61352
rect 2786 61076 2820 61132
rect 3238 61076 3272 61352
rect 2786 61036 3272 61076
rect 2786 60980 2820 61036
rect 2786 60760 2820 60822
rect 3238 60760 3272 61036
rect 2786 60726 3272 60760
rect 7776 61352 8262 61386
rect 7776 61290 7810 61352
rect 7776 61076 7810 61132
rect 8228 61076 8262 61352
rect 7776 61036 8262 61076
rect 7776 60980 7810 61036
rect 7776 60760 7810 60822
rect 8228 60760 8262 61036
rect 7776 60726 8262 60760
rect 12766 61352 13252 61386
rect 12766 61290 12800 61352
rect 12766 61076 12800 61132
rect 13218 61076 13252 61352
rect 12766 61036 13252 61076
rect 12766 60980 12800 61036
rect 12766 60760 12800 60822
rect 13218 60760 13252 61036
rect 12766 60726 13252 60760
rect 17756 61352 18242 61386
rect 17756 61290 17790 61352
rect 17756 61076 17790 61132
rect 18208 61076 18242 61352
rect 17756 61036 18242 61076
rect 17756 60980 17790 61036
rect 17756 60760 17790 60822
rect 18208 60760 18242 61036
rect 17756 60726 18242 60760
rect 22746 61352 23232 61386
rect 22746 61290 22780 61352
rect 22746 61076 22780 61132
rect 23198 61076 23232 61352
rect 22746 61036 23232 61076
rect 22746 60980 22780 61036
rect 22746 60760 22780 60822
rect 23198 60760 23232 61036
rect 22746 60726 23232 60760
rect 27736 61352 28222 61386
rect 27736 61290 27770 61352
rect 27736 61076 27770 61132
rect 28188 61076 28222 61352
rect 27736 61036 28222 61076
rect 27736 60980 27770 61036
rect 27736 60760 27770 60822
rect 28188 60760 28222 61036
rect 27736 60726 28222 60760
rect 32726 61352 33212 61386
rect 32726 61290 32760 61352
rect 32726 61076 32760 61132
rect 33178 61076 33212 61352
rect 32726 61036 33212 61076
rect 32726 60980 32760 61036
rect 32726 60760 32760 60822
rect 33178 60760 33212 61036
rect 32726 60726 33212 60760
rect 37716 61352 38202 61386
rect 37716 61290 37750 61352
rect 37716 61076 37750 61132
rect 38168 61076 38202 61352
rect 37716 61036 38202 61076
rect 37716 60980 37750 61036
rect 37716 60760 37750 60822
rect 38168 60760 38202 61036
rect 37716 60726 38202 60760
rect 42706 61352 43192 61386
rect 42706 61290 42740 61352
rect 42706 61076 42740 61132
rect 43158 61076 43192 61352
rect 42706 61036 43192 61076
rect 42706 60980 42740 61036
rect 42706 60760 42740 60822
rect 43158 60760 43192 61036
rect 42706 60726 43192 60760
rect 47696 61352 48182 61386
rect 47696 61290 47730 61352
rect 47696 61076 47730 61132
rect 48148 61076 48182 61352
rect 47696 61036 48182 61076
rect 47696 60980 47730 61036
rect 47696 60760 47730 60822
rect 48148 60760 48182 61036
rect 47696 60726 48182 60760
rect 52686 61352 53172 61386
rect 52686 61290 52720 61352
rect 52686 61076 52720 61132
rect 53138 61076 53172 61352
rect 52686 61036 53172 61076
rect 52686 60980 52720 61036
rect 52686 60760 52720 60822
rect 53138 60760 53172 61036
rect 52686 60726 53172 60760
rect 57676 61352 58162 61386
rect 57676 61290 57710 61352
rect 57676 61076 57710 61132
rect 58128 61076 58162 61352
rect 57676 61036 58162 61076
rect 57676 60980 57710 61036
rect 57676 60760 57710 60822
rect 58128 60760 58162 61036
rect 57676 60726 58162 60760
rect 62666 61352 63152 61386
rect 62666 61290 62700 61352
rect 62666 61076 62700 61132
rect 63118 61076 63152 61352
rect 62666 61036 63152 61076
rect 62666 60980 62700 61036
rect 62666 60760 62700 60822
rect 63118 60760 63152 61036
rect 62666 60726 63152 60760
rect 67656 61352 68142 61386
rect 67656 61290 67690 61352
rect 67656 61076 67690 61132
rect 68108 61076 68142 61352
rect 67656 61036 68142 61076
rect 67656 60980 67690 61036
rect 67656 60760 67690 60822
rect 68108 60760 68142 61036
rect 67656 60726 68142 60760
rect 72646 61352 73132 61386
rect 72646 61290 72680 61352
rect 72646 61076 72680 61132
rect 73098 61076 73132 61352
rect 72646 61036 73132 61076
rect 72646 60980 72680 61036
rect 72646 60760 72680 60822
rect 73098 60760 73132 61036
rect 72646 60726 73132 60760
rect 77636 61352 78122 61386
rect 77636 61290 77670 61352
rect 77636 61076 77670 61132
rect 78088 61076 78122 61352
rect 77636 61036 78122 61076
rect 77636 60980 77670 61036
rect 77636 60760 77670 60822
rect 78088 60760 78122 61036
rect 77636 60726 78122 60760
rect 2786 59642 3272 59676
rect 2786 59580 2820 59642
rect 2786 59366 2820 59422
rect 3238 59366 3272 59642
rect 2786 59326 3272 59366
rect 2786 59270 2820 59326
rect 2786 59050 2820 59112
rect 3238 59050 3272 59326
rect 2786 59016 3272 59050
rect 7776 59642 8262 59676
rect 7776 59580 7810 59642
rect 7776 59366 7810 59422
rect 8228 59366 8262 59642
rect 7776 59326 8262 59366
rect 7776 59270 7810 59326
rect 7776 59050 7810 59112
rect 8228 59050 8262 59326
rect 7776 59016 8262 59050
rect 12766 59642 13252 59676
rect 12766 59580 12800 59642
rect 12766 59366 12800 59422
rect 13218 59366 13252 59642
rect 12766 59326 13252 59366
rect 12766 59270 12800 59326
rect 12766 59050 12800 59112
rect 13218 59050 13252 59326
rect 12766 59016 13252 59050
rect 17756 59642 18242 59676
rect 17756 59580 17790 59642
rect 17756 59366 17790 59422
rect 18208 59366 18242 59642
rect 17756 59326 18242 59366
rect 17756 59270 17790 59326
rect 17756 59050 17790 59112
rect 18208 59050 18242 59326
rect 17756 59016 18242 59050
rect 22746 59642 23232 59676
rect 22746 59580 22780 59642
rect 22746 59366 22780 59422
rect 23198 59366 23232 59642
rect 22746 59326 23232 59366
rect 22746 59270 22780 59326
rect 22746 59050 22780 59112
rect 23198 59050 23232 59326
rect 22746 59016 23232 59050
rect 27736 59642 28222 59676
rect 27736 59580 27770 59642
rect 27736 59366 27770 59422
rect 28188 59366 28222 59642
rect 27736 59326 28222 59366
rect 27736 59270 27770 59326
rect 27736 59050 27770 59112
rect 28188 59050 28222 59326
rect 27736 59016 28222 59050
rect 32726 59642 33212 59676
rect 32726 59580 32760 59642
rect 32726 59366 32760 59422
rect 33178 59366 33212 59642
rect 32726 59326 33212 59366
rect 32726 59270 32760 59326
rect 32726 59050 32760 59112
rect 33178 59050 33212 59326
rect 32726 59016 33212 59050
rect 37716 59642 38202 59676
rect 37716 59580 37750 59642
rect 37716 59366 37750 59422
rect 38168 59366 38202 59642
rect 37716 59326 38202 59366
rect 37716 59270 37750 59326
rect 37716 59050 37750 59112
rect 38168 59050 38202 59326
rect 37716 59016 38202 59050
rect 42706 59642 43192 59676
rect 42706 59580 42740 59642
rect 42706 59366 42740 59422
rect 43158 59366 43192 59642
rect 42706 59326 43192 59366
rect 42706 59270 42740 59326
rect 42706 59050 42740 59112
rect 43158 59050 43192 59326
rect 42706 59016 43192 59050
rect 47696 59642 48182 59676
rect 47696 59580 47730 59642
rect 47696 59366 47730 59422
rect 48148 59366 48182 59642
rect 47696 59326 48182 59366
rect 47696 59270 47730 59326
rect 47696 59050 47730 59112
rect 48148 59050 48182 59326
rect 47696 59016 48182 59050
rect 52686 59642 53172 59676
rect 52686 59580 52720 59642
rect 52686 59366 52720 59422
rect 53138 59366 53172 59642
rect 52686 59326 53172 59366
rect 52686 59270 52720 59326
rect 52686 59050 52720 59112
rect 53138 59050 53172 59326
rect 52686 59016 53172 59050
rect 57676 59642 58162 59676
rect 57676 59580 57710 59642
rect 57676 59366 57710 59422
rect 58128 59366 58162 59642
rect 57676 59326 58162 59366
rect 57676 59270 57710 59326
rect 57676 59050 57710 59112
rect 58128 59050 58162 59326
rect 57676 59016 58162 59050
rect 62666 59642 63152 59676
rect 62666 59580 62700 59642
rect 62666 59366 62700 59422
rect 63118 59366 63152 59642
rect 62666 59326 63152 59366
rect 62666 59270 62700 59326
rect 62666 59050 62700 59112
rect 63118 59050 63152 59326
rect 62666 59016 63152 59050
rect 67656 59642 68142 59676
rect 67656 59580 67690 59642
rect 67656 59366 67690 59422
rect 68108 59366 68142 59642
rect 67656 59326 68142 59366
rect 67656 59270 67690 59326
rect 67656 59050 67690 59112
rect 68108 59050 68142 59326
rect 67656 59016 68142 59050
rect 72646 59642 73132 59676
rect 72646 59580 72680 59642
rect 72646 59366 72680 59422
rect 73098 59366 73132 59642
rect 72646 59326 73132 59366
rect 72646 59270 72680 59326
rect 72646 59050 72680 59112
rect 73098 59050 73132 59326
rect 72646 59016 73132 59050
rect 77636 59642 78122 59676
rect 77636 59580 77670 59642
rect 77636 59366 77670 59422
rect 78088 59366 78122 59642
rect 77636 59326 78122 59366
rect 77636 59270 77670 59326
rect 77636 59050 77670 59112
rect 78088 59050 78122 59326
rect 77636 59016 78122 59050
rect 2786 57932 3272 57966
rect 2786 57870 2820 57932
rect 2786 57656 2820 57712
rect 3238 57656 3272 57932
rect 2786 57616 3272 57656
rect 2786 57560 2820 57616
rect 2786 57340 2820 57402
rect 3238 57340 3272 57616
rect 2786 57306 3272 57340
rect 7776 57932 8262 57966
rect 7776 57870 7810 57932
rect 7776 57656 7810 57712
rect 8228 57656 8262 57932
rect 7776 57616 8262 57656
rect 7776 57560 7810 57616
rect 7776 57340 7810 57402
rect 8228 57340 8262 57616
rect 7776 57306 8262 57340
rect 12766 57932 13252 57966
rect 12766 57870 12800 57932
rect 12766 57656 12800 57712
rect 13218 57656 13252 57932
rect 12766 57616 13252 57656
rect 12766 57560 12800 57616
rect 12766 57340 12800 57402
rect 13218 57340 13252 57616
rect 12766 57306 13252 57340
rect 17756 57932 18242 57966
rect 17756 57870 17790 57932
rect 17756 57656 17790 57712
rect 18208 57656 18242 57932
rect 17756 57616 18242 57656
rect 17756 57560 17790 57616
rect 17756 57340 17790 57402
rect 18208 57340 18242 57616
rect 17756 57306 18242 57340
rect 22746 57932 23232 57966
rect 22746 57870 22780 57932
rect 22746 57656 22780 57712
rect 23198 57656 23232 57932
rect 22746 57616 23232 57656
rect 22746 57560 22780 57616
rect 22746 57340 22780 57402
rect 23198 57340 23232 57616
rect 22746 57306 23232 57340
rect 27736 57932 28222 57966
rect 27736 57870 27770 57932
rect 27736 57656 27770 57712
rect 28188 57656 28222 57932
rect 27736 57616 28222 57656
rect 27736 57560 27770 57616
rect 27736 57340 27770 57402
rect 28188 57340 28222 57616
rect 27736 57306 28222 57340
rect 32726 57932 33212 57966
rect 32726 57870 32760 57932
rect 32726 57656 32760 57712
rect 33178 57656 33212 57932
rect 32726 57616 33212 57656
rect 32726 57560 32760 57616
rect 32726 57340 32760 57402
rect 33178 57340 33212 57616
rect 32726 57306 33212 57340
rect 37716 57932 38202 57966
rect 37716 57870 37750 57932
rect 37716 57656 37750 57712
rect 38168 57656 38202 57932
rect 37716 57616 38202 57656
rect 37716 57560 37750 57616
rect 37716 57340 37750 57402
rect 38168 57340 38202 57616
rect 37716 57306 38202 57340
rect 42706 57932 43192 57966
rect 42706 57870 42740 57932
rect 42706 57656 42740 57712
rect 43158 57656 43192 57932
rect 42706 57616 43192 57656
rect 42706 57560 42740 57616
rect 42706 57340 42740 57402
rect 43158 57340 43192 57616
rect 42706 57306 43192 57340
rect 47696 57932 48182 57966
rect 47696 57870 47730 57932
rect 47696 57656 47730 57712
rect 48148 57656 48182 57932
rect 47696 57616 48182 57656
rect 47696 57560 47730 57616
rect 47696 57340 47730 57402
rect 48148 57340 48182 57616
rect 47696 57306 48182 57340
rect 52686 57932 53172 57966
rect 52686 57870 52720 57932
rect 52686 57656 52720 57712
rect 53138 57656 53172 57932
rect 52686 57616 53172 57656
rect 52686 57560 52720 57616
rect 52686 57340 52720 57402
rect 53138 57340 53172 57616
rect 52686 57306 53172 57340
rect 57676 57932 58162 57966
rect 57676 57870 57710 57932
rect 57676 57656 57710 57712
rect 58128 57656 58162 57932
rect 57676 57616 58162 57656
rect 57676 57560 57710 57616
rect 57676 57340 57710 57402
rect 58128 57340 58162 57616
rect 57676 57306 58162 57340
rect 62666 57932 63152 57966
rect 62666 57870 62700 57932
rect 62666 57656 62700 57712
rect 63118 57656 63152 57932
rect 62666 57616 63152 57656
rect 62666 57560 62700 57616
rect 62666 57340 62700 57402
rect 63118 57340 63152 57616
rect 62666 57306 63152 57340
rect 67656 57932 68142 57966
rect 67656 57870 67690 57932
rect 67656 57656 67690 57712
rect 68108 57656 68142 57932
rect 67656 57616 68142 57656
rect 67656 57560 67690 57616
rect 67656 57340 67690 57402
rect 68108 57340 68142 57616
rect 67656 57306 68142 57340
rect 72646 57932 73132 57966
rect 72646 57870 72680 57932
rect 72646 57656 72680 57712
rect 73098 57656 73132 57932
rect 72646 57616 73132 57656
rect 72646 57560 72680 57616
rect 72646 57340 72680 57402
rect 73098 57340 73132 57616
rect 72646 57306 73132 57340
rect 77636 57932 78122 57966
rect 77636 57870 77670 57932
rect 77636 57656 77670 57712
rect 78088 57656 78122 57932
rect 77636 57616 78122 57656
rect 77636 57560 77670 57616
rect 77636 57340 77670 57402
rect 78088 57340 78122 57616
rect 77636 57306 78122 57340
rect 2786 56222 3272 56256
rect 2786 56160 2820 56222
rect 2786 55946 2820 56002
rect 3238 55946 3272 56222
rect 2786 55906 3272 55946
rect 2786 55850 2820 55906
rect 2786 55630 2820 55692
rect 3238 55630 3272 55906
rect 2786 55596 3272 55630
rect 7776 56222 8262 56256
rect 7776 56160 7810 56222
rect 7776 55946 7810 56002
rect 8228 55946 8262 56222
rect 7776 55906 8262 55946
rect 7776 55850 7810 55906
rect 7776 55630 7810 55692
rect 8228 55630 8262 55906
rect 7776 55596 8262 55630
rect 12766 56222 13252 56256
rect 12766 56160 12800 56222
rect 12766 55946 12800 56002
rect 13218 55946 13252 56222
rect 12766 55906 13252 55946
rect 12766 55850 12800 55906
rect 12766 55630 12800 55692
rect 13218 55630 13252 55906
rect 12766 55596 13252 55630
rect 17756 56222 18242 56256
rect 17756 56160 17790 56222
rect 17756 55946 17790 56002
rect 18208 55946 18242 56222
rect 17756 55906 18242 55946
rect 17756 55850 17790 55906
rect 17756 55630 17790 55692
rect 18208 55630 18242 55906
rect 17756 55596 18242 55630
rect 22746 56222 23232 56256
rect 22746 56160 22780 56222
rect 22746 55946 22780 56002
rect 23198 55946 23232 56222
rect 22746 55906 23232 55946
rect 22746 55850 22780 55906
rect 22746 55630 22780 55692
rect 23198 55630 23232 55906
rect 22746 55596 23232 55630
rect 27736 56222 28222 56256
rect 27736 56160 27770 56222
rect 27736 55946 27770 56002
rect 28188 55946 28222 56222
rect 27736 55906 28222 55946
rect 27736 55850 27770 55906
rect 27736 55630 27770 55692
rect 28188 55630 28222 55906
rect 27736 55596 28222 55630
rect 32726 56222 33212 56256
rect 32726 56160 32760 56222
rect 32726 55946 32760 56002
rect 33178 55946 33212 56222
rect 32726 55906 33212 55946
rect 32726 55850 32760 55906
rect 32726 55630 32760 55692
rect 33178 55630 33212 55906
rect 32726 55596 33212 55630
rect 37716 56222 38202 56256
rect 37716 56160 37750 56222
rect 37716 55946 37750 56002
rect 38168 55946 38202 56222
rect 37716 55906 38202 55946
rect 37716 55850 37750 55906
rect 37716 55630 37750 55692
rect 38168 55630 38202 55906
rect 37716 55596 38202 55630
rect 42706 56222 43192 56256
rect 42706 56160 42740 56222
rect 42706 55946 42740 56002
rect 43158 55946 43192 56222
rect 42706 55906 43192 55946
rect 42706 55850 42740 55906
rect 42706 55630 42740 55692
rect 43158 55630 43192 55906
rect 42706 55596 43192 55630
rect 47696 56222 48182 56256
rect 47696 56160 47730 56222
rect 47696 55946 47730 56002
rect 48148 55946 48182 56222
rect 47696 55906 48182 55946
rect 47696 55850 47730 55906
rect 47696 55630 47730 55692
rect 48148 55630 48182 55906
rect 47696 55596 48182 55630
rect 52686 56222 53172 56256
rect 52686 56160 52720 56222
rect 52686 55946 52720 56002
rect 53138 55946 53172 56222
rect 52686 55906 53172 55946
rect 52686 55850 52720 55906
rect 52686 55630 52720 55692
rect 53138 55630 53172 55906
rect 52686 55596 53172 55630
rect 57676 56222 58162 56256
rect 57676 56160 57710 56222
rect 57676 55946 57710 56002
rect 58128 55946 58162 56222
rect 57676 55906 58162 55946
rect 57676 55850 57710 55906
rect 57676 55630 57710 55692
rect 58128 55630 58162 55906
rect 57676 55596 58162 55630
rect 62666 56222 63152 56256
rect 62666 56160 62700 56222
rect 62666 55946 62700 56002
rect 63118 55946 63152 56222
rect 62666 55906 63152 55946
rect 62666 55850 62700 55906
rect 62666 55630 62700 55692
rect 63118 55630 63152 55906
rect 62666 55596 63152 55630
rect 67656 56222 68142 56256
rect 67656 56160 67690 56222
rect 67656 55946 67690 56002
rect 68108 55946 68142 56222
rect 67656 55906 68142 55946
rect 67656 55850 67690 55906
rect 67656 55630 67690 55692
rect 68108 55630 68142 55906
rect 67656 55596 68142 55630
rect 72646 56222 73132 56256
rect 72646 56160 72680 56222
rect 72646 55946 72680 56002
rect 73098 55946 73132 56222
rect 72646 55906 73132 55946
rect 72646 55850 72680 55906
rect 72646 55630 72680 55692
rect 73098 55630 73132 55906
rect 72646 55596 73132 55630
rect 77636 56222 78122 56256
rect 77636 56160 77670 56222
rect 77636 55946 77670 56002
rect 78088 55946 78122 56222
rect 77636 55906 78122 55946
rect 77636 55850 77670 55906
rect 77636 55630 77670 55692
rect 78088 55630 78122 55906
rect 77636 55596 78122 55630
rect 2786 54512 3272 54546
rect 2786 54450 2820 54512
rect 2786 54236 2820 54292
rect 3238 54236 3272 54512
rect 2786 54196 3272 54236
rect 2786 54140 2820 54196
rect 2786 53920 2820 53982
rect 3238 53920 3272 54196
rect 2786 53886 3272 53920
rect 7776 54512 8262 54546
rect 7776 54450 7810 54512
rect 7776 54236 7810 54292
rect 8228 54236 8262 54512
rect 7776 54196 8262 54236
rect 7776 54140 7810 54196
rect 7776 53920 7810 53982
rect 8228 53920 8262 54196
rect 7776 53886 8262 53920
rect 12766 54512 13252 54546
rect 12766 54450 12800 54512
rect 12766 54236 12800 54292
rect 13218 54236 13252 54512
rect 12766 54196 13252 54236
rect 12766 54140 12800 54196
rect 12766 53920 12800 53982
rect 13218 53920 13252 54196
rect 12766 53886 13252 53920
rect 17756 54512 18242 54546
rect 17756 54450 17790 54512
rect 17756 54236 17790 54292
rect 18208 54236 18242 54512
rect 17756 54196 18242 54236
rect 17756 54140 17790 54196
rect 17756 53920 17790 53982
rect 18208 53920 18242 54196
rect 17756 53886 18242 53920
rect 22746 54512 23232 54546
rect 22746 54450 22780 54512
rect 22746 54236 22780 54292
rect 23198 54236 23232 54512
rect 22746 54196 23232 54236
rect 22746 54140 22780 54196
rect 22746 53920 22780 53982
rect 23198 53920 23232 54196
rect 22746 53886 23232 53920
rect 27736 54512 28222 54546
rect 27736 54450 27770 54512
rect 27736 54236 27770 54292
rect 28188 54236 28222 54512
rect 27736 54196 28222 54236
rect 27736 54140 27770 54196
rect 27736 53920 27770 53982
rect 28188 53920 28222 54196
rect 27736 53886 28222 53920
rect 32726 54512 33212 54546
rect 32726 54450 32760 54512
rect 32726 54236 32760 54292
rect 33178 54236 33212 54512
rect 32726 54196 33212 54236
rect 32726 54140 32760 54196
rect 32726 53920 32760 53982
rect 33178 53920 33212 54196
rect 32726 53886 33212 53920
rect 37716 54512 38202 54546
rect 37716 54450 37750 54512
rect 37716 54236 37750 54292
rect 38168 54236 38202 54512
rect 37716 54196 38202 54236
rect 37716 54140 37750 54196
rect 37716 53920 37750 53982
rect 38168 53920 38202 54196
rect 37716 53886 38202 53920
rect 42706 54512 43192 54546
rect 42706 54450 42740 54512
rect 42706 54236 42740 54292
rect 43158 54236 43192 54512
rect 42706 54196 43192 54236
rect 42706 54140 42740 54196
rect 42706 53920 42740 53982
rect 43158 53920 43192 54196
rect 42706 53886 43192 53920
rect 47696 54512 48182 54546
rect 47696 54450 47730 54512
rect 47696 54236 47730 54292
rect 48148 54236 48182 54512
rect 47696 54196 48182 54236
rect 47696 54140 47730 54196
rect 47696 53920 47730 53982
rect 48148 53920 48182 54196
rect 47696 53886 48182 53920
rect 52686 54512 53172 54546
rect 52686 54450 52720 54512
rect 52686 54236 52720 54292
rect 53138 54236 53172 54512
rect 52686 54196 53172 54236
rect 52686 54140 52720 54196
rect 52686 53920 52720 53982
rect 53138 53920 53172 54196
rect 52686 53886 53172 53920
rect 57676 54512 58162 54546
rect 57676 54450 57710 54512
rect 57676 54236 57710 54292
rect 58128 54236 58162 54512
rect 57676 54196 58162 54236
rect 57676 54140 57710 54196
rect 57676 53920 57710 53982
rect 58128 53920 58162 54196
rect 57676 53886 58162 53920
rect 62666 54512 63152 54546
rect 62666 54450 62700 54512
rect 62666 54236 62700 54292
rect 63118 54236 63152 54512
rect 62666 54196 63152 54236
rect 62666 54140 62700 54196
rect 62666 53920 62700 53982
rect 63118 53920 63152 54196
rect 62666 53886 63152 53920
rect 67656 54512 68142 54546
rect 67656 54450 67690 54512
rect 67656 54236 67690 54292
rect 68108 54236 68142 54512
rect 67656 54196 68142 54236
rect 67656 54140 67690 54196
rect 67656 53920 67690 53982
rect 68108 53920 68142 54196
rect 67656 53886 68142 53920
rect 72646 54512 73132 54546
rect 72646 54450 72680 54512
rect 72646 54236 72680 54292
rect 73098 54236 73132 54512
rect 72646 54196 73132 54236
rect 72646 54140 72680 54196
rect 72646 53920 72680 53982
rect 73098 53920 73132 54196
rect 72646 53886 73132 53920
rect 77636 54512 78122 54546
rect 77636 54450 77670 54512
rect 77636 54236 77670 54292
rect 78088 54236 78122 54512
rect 77636 54196 78122 54236
rect 77636 54140 77670 54196
rect 77636 53920 77670 53982
rect 78088 53920 78122 54196
rect 77636 53886 78122 53920
rect 2786 52802 3272 52836
rect 2786 52740 2820 52802
rect 2786 52526 2820 52582
rect 3238 52526 3272 52802
rect 2786 52486 3272 52526
rect 2786 52430 2820 52486
rect 2786 52210 2820 52272
rect 3238 52210 3272 52486
rect 2786 52176 3272 52210
rect 7776 52802 8262 52836
rect 7776 52740 7810 52802
rect 7776 52526 7810 52582
rect 8228 52526 8262 52802
rect 7776 52486 8262 52526
rect 7776 52430 7810 52486
rect 7776 52210 7810 52272
rect 8228 52210 8262 52486
rect 7776 52176 8262 52210
rect 12766 52802 13252 52836
rect 12766 52740 12800 52802
rect 12766 52526 12800 52582
rect 13218 52526 13252 52802
rect 12766 52486 13252 52526
rect 12766 52430 12800 52486
rect 12766 52210 12800 52272
rect 13218 52210 13252 52486
rect 12766 52176 13252 52210
rect 17756 52802 18242 52836
rect 17756 52740 17790 52802
rect 17756 52526 17790 52582
rect 18208 52526 18242 52802
rect 17756 52486 18242 52526
rect 17756 52430 17790 52486
rect 17756 52210 17790 52272
rect 18208 52210 18242 52486
rect 17756 52176 18242 52210
rect 22746 52802 23232 52836
rect 22746 52740 22780 52802
rect 22746 52526 22780 52582
rect 23198 52526 23232 52802
rect 22746 52486 23232 52526
rect 22746 52430 22780 52486
rect 22746 52210 22780 52272
rect 23198 52210 23232 52486
rect 22746 52176 23232 52210
rect 27736 52802 28222 52836
rect 27736 52740 27770 52802
rect 27736 52526 27770 52582
rect 28188 52526 28222 52802
rect 27736 52486 28222 52526
rect 27736 52430 27770 52486
rect 27736 52210 27770 52272
rect 28188 52210 28222 52486
rect 27736 52176 28222 52210
rect 32726 52802 33212 52836
rect 32726 52740 32760 52802
rect 32726 52526 32760 52582
rect 33178 52526 33212 52802
rect 32726 52486 33212 52526
rect 32726 52430 32760 52486
rect 32726 52210 32760 52272
rect 33178 52210 33212 52486
rect 32726 52176 33212 52210
rect 37716 52802 38202 52836
rect 37716 52740 37750 52802
rect 37716 52526 37750 52582
rect 38168 52526 38202 52802
rect 37716 52486 38202 52526
rect 37716 52430 37750 52486
rect 37716 52210 37750 52272
rect 38168 52210 38202 52486
rect 37716 52176 38202 52210
rect 42706 52802 43192 52836
rect 42706 52740 42740 52802
rect 42706 52526 42740 52582
rect 43158 52526 43192 52802
rect 42706 52486 43192 52526
rect 42706 52430 42740 52486
rect 42706 52210 42740 52272
rect 43158 52210 43192 52486
rect 42706 52176 43192 52210
rect 47696 52802 48182 52836
rect 47696 52740 47730 52802
rect 47696 52526 47730 52582
rect 48148 52526 48182 52802
rect 47696 52486 48182 52526
rect 47696 52430 47730 52486
rect 47696 52210 47730 52272
rect 48148 52210 48182 52486
rect 47696 52176 48182 52210
rect 52686 52802 53172 52836
rect 52686 52740 52720 52802
rect 52686 52526 52720 52582
rect 53138 52526 53172 52802
rect 52686 52486 53172 52526
rect 52686 52430 52720 52486
rect 52686 52210 52720 52272
rect 53138 52210 53172 52486
rect 52686 52176 53172 52210
rect 57676 52802 58162 52836
rect 57676 52740 57710 52802
rect 57676 52526 57710 52582
rect 58128 52526 58162 52802
rect 57676 52486 58162 52526
rect 57676 52430 57710 52486
rect 57676 52210 57710 52272
rect 58128 52210 58162 52486
rect 57676 52176 58162 52210
rect 62666 52802 63152 52836
rect 62666 52740 62700 52802
rect 62666 52526 62700 52582
rect 63118 52526 63152 52802
rect 62666 52486 63152 52526
rect 62666 52430 62700 52486
rect 62666 52210 62700 52272
rect 63118 52210 63152 52486
rect 62666 52176 63152 52210
rect 67656 52802 68142 52836
rect 67656 52740 67690 52802
rect 67656 52526 67690 52582
rect 68108 52526 68142 52802
rect 67656 52486 68142 52526
rect 67656 52430 67690 52486
rect 67656 52210 67690 52272
rect 68108 52210 68142 52486
rect 67656 52176 68142 52210
rect 72646 52802 73132 52836
rect 72646 52740 72680 52802
rect 72646 52526 72680 52582
rect 73098 52526 73132 52802
rect 72646 52486 73132 52526
rect 72646 52430 72680 52486
rect 72646 52210 72680 52272
rect 73098 52210 73132 52486
rect 72646 52176 73132 52210
rect 77636 52802 78122 52836
rect 77636 52740 77670 52802
rect 77636 52526 77670 52582
rect 78088 52526 78122 52802
rect 77636 52486 78122 52526
rect 77636 52430 77670 52486
rect 77636 52210 77670 52272
rect 78088 52210 78122 52486
rect 77636 52176 78122 52210
rect 2786 51092 3272 51126
rect 2786 51030 2820 51092
rect 2786 50816 2820 50872
rect 3238 50816 3272 51092
rect 2786 50776 3272 50816
rect 2786 50720 2820 50776
rect 2786 50500 2820 50562
rect 3238 50500 3272 50776
rect 2786 50466 3272 50500
rect 7776 51092 8262 51126
rect 7776 51030 7810 51092
rect 7776 50816 7810 50872
rect 8228 50816 8262 51092
rect 7776 50776 8262 50816
rect 7776 50720 7810 50776
rect 7776 50500 7810 50562
rect 8228 50500 8262 50776
rect 7776 50466 8262 50500
rect 12766 51092 13252 51126
rect 12766 51030 12800 51092
rect 12766 50816 12800 50872
rect 13218 50816 13252 51092
rect 12766 50776 13252 50816
rect 12766 50720 12800 50776
rect 12766 50500 12800 50562
rect 13218 50500 13252 50776
rect 12766 50466 13252 50500
rect 17756 51092 18242 51126
rect 17756 51030 17790 51092
rect 17756 50816 17790 50872
rect 18208 50816 18242 51092
rect 17756 50776 18242 50816
rect 17756 50720 17790 50776
rect 17756 50500 17790 50562
rect 18208 50500 18242 50776
rect 17756 50466 18242 50500
rect 22746 51092 23232 51126
rect 22746 51030 22780 51092
rect 22746 50816 22780 50872
rect 23198 50816 23232 51092
rect 22746 50776 23232 50816
rect 22746 50720 22780 50776
rect 22746 50500 22780 50562
rect 23198 50500 23232 50776
rect 22746 50466 23232 50500
rect 27736 51092 28222 51126
rect 27736 51030 27770 51092
rect 27736 50816 27770 50872
rect 28188 50816 28222 51092
rect 27736 50776 28222 50816
rect 27736 50720 27770 50776
rect 27736 50500 27770 50562
rect 28188 50500 28222 50776
rect 27736 50466 28222 50500
rect 32726 51092 33212 51126
rect 32726 51030 32760 51092
rect 32726 50816 32760 50872
rect 33178 50816 33212 51092
rect 32726 50776 33212 50816
rect 32726 50720 32760 50776
rect 32726 50500 32760 50562
rect 33178 50500 33212 50776
rect 32726 50466 33212 50500
rect 37716 51092 38202 51126
rect 37716 51030 37750 51092
rect 37716 50816 37750 50872
rect 38168 50816 38202 51092
rect 37716 50776 38202 50816
rect 37716 50720 37750 50776
rect 37716 50500 37750 50562
rect 38168 50500 38202 50776
rect 37716 50466 38202 50500
rect 42706 51092 43192 51126
rect 42706 51030 42740 51092
rect 42706 50816 42740 50872
rect 43158 50816 43192 51092
rect 42706 50776 43192 50816
rect 42706 50720 42740 50776
rect 42706 50500 42740 50562
rect 43158 50500 43192 50776
rect 42706 50466 43192 50500
rect 47696 51092 48182 51126
rect 47696 51030 47730 51092
rect 47696 50816 47730 50872
rect 48148 50816 48182 51092
rect 47696 50776 48182 50816
rect 47696 50720 47730 50776
rect 47696 50500 47730 50562
rect 48148 50500 48182 50776
rect 47696 50466 48182 50500
rect 52686 51092 53172 51126
rect 52686 51030 52720 51092
rect 52686 50816 52720 50872
rect 53138 50816 53172 51092
rect 52686 50776 53172 50816
rect 52686 50720 52720 50776
rect 52686 50500 52720 50562
rect 53138 50500 53172 50776
rect 52686 50466 53172 50500
rect 57676 51092 58162 51126
rect 57676 51030 57710 51092
rect 57676 50816 57710 50872
rect 58128 50816 58162 51092
rect 57676 50776 58162 50816
rect 57676 50720 57710 50776
rect 57676 50500 57710 50562
rect 58128 50500 58162 50776
rect 57676 50466 58162 50500
rect 62666 51092 63152 51126
rect 62666 51030 62700 51092
rect 62666 50816 62700 50872
rect 63118 50816 63152 51092
rect 62666 50776 63152 50816
rect 62666 50720 62700 50776
rect 62666 50500 62700 50562
rect 63118 50500 63152 50776
rect 62666 50466 63152 50500
rect 67656 51092 68142 51126
rect 67656 51030 67690 51092
rect 67656 50816 67690 50872
rect 68108 50816 68142 51092
rect 67656 50776 68142 50816
rect 67656 50720 67690 50776
rect 67656 50500 67690 50562
rect 68108 50500 68142 50776
rect 67656 50466 68142 50500
rect 72646 51092 73132 51126
rect 72646 51030 72680 51092
rect 72646 50816 72680 50872
rect 73098 50816 73132 51092
rect 72646 50776 73132 50816
rect 72646 50720 72680 50776
rect 72646 50500 72680 50562
rect 73098 50500 73132 50776
rect 72646 50466 73132 50500
rect 77636 51092 78122 51126
rect 77636 51030 77670 51092
rect 77636 50816 77670 50872
rect 78088 50816 78122 51092
rect 77636 50776 78122 50816
rect 77636 50720 77670 50776
rect 77636 50500 77670 50562
rect 78088 50500 78122 50776
rect 77636 50466 78122 50500
rect 2786 49382 3272 49416
rect 2786 49320 2820 49382
rect 2786 49106 2820 49162
rect 3238 49106 3272 49382
rect 2786 49066 3272 49106
rect 2786 49010 2820 49066
rect 2786 48790 2820 48852
rect 3238 48790 3272 49066
rect 2786 48756 3272 48790
rect 7776 49382 8262 49416
rect 7776 49320 7810 49382
rect 7776 49106 7810 49162
rect 8228 49106 8262 49382
rect 7776 49066 8262 49106
rect 7776 49010 7810 49066
rect 7776 48790 7810 48852
rect 8228 48790 8262 49066
rect 7776 48756 8262 48790
rect 12766 49382 13252 49416
rect 12766 49320 12800 49382
rect 12766 49106 12800 49162
rect 13218 49106 13252 49382
rect 12766 49066 13252 49106
rect 12766 49010 12800 49066
rect 12766 48790 12800 48852
rect 13218 48790 13252 49066
rect 12766 48756 13252 48790
rect 17756 49382 18242 49416
rect 17756 49320 17790 49382
rect 17756 49106 17790 49162
rect 18208 49106 18242 49382
rect 17756 49066 18242 49106
rect 17756 49010 17790 49066
rect 17756 48790 17790 48852
rect 18208 48790 18242 49066
rect 17756 48756 18242 48790
rect 22746 49382 23232 49416
rect 22746 49320 22780 49382
rect 22746 49106 22780 49162
rect 23198 49106 23232 49382
rect 22746 49066 23232 49106
rect 22746 49010 22780 49066
rect 22746 48790 22780 48852
rect 23198 48790 23232 49066
rect 22746 48756 23232 48790
rect 27736 49382 28222 49416
rect 27736 49320 27770 49382
rect 27736 49106 27770 49162
rect 28188 49106 28222 49382
rect 27736 49066 28222 49106
rect 27736 49010 27770 49066
rect 27736 48790 27770 48852
rect 28188 48790 28222 49066
rect 27736 48756 28222 48790
rect 32726 49382 33212 49416
rect 32726 49320 32760 49382
rect 32726 49106 32760 49162
rect 33178 49106 33212 49382
rect 32726 49066 33212 49106
rect 32726 49010 32760 49066
rect 32726 48790 32760 48852
rect 33178 48790 33212 49066
rect 32726 48756 33212 48790
rect 37716 49382 38202 49416
rect 37716 49320 37750 49382
rect 37716 49106 37750 49162
rect 38168 49106 38202 49382
rect 37716 49066 38202 49106
rect 37716 49010 37750 49066
rect 37716 48790 37750 48852
rect 38168 48790 38202 49066
rect 37716 48756 38202 48790
rect 42706 49382 43192 49416
rect 42706 49320 42740 49382
rect 42706 49106 42740 49162
rect 43158 49106 43192 49382
rect 42706 49066 43192 49106
rect 42706 49010 42740 49066
rect 42706 48790 42740 48852
rect 43158 48790 43192 49066
rect 42706 48756 43192 48790
rect 47696 49382 48182 49416
rect 47696 49320 47730 49382
rect 47696 49106 47730 49162
rect 48148 49106 48182 49382
rect 47696 49066 48182 49106
rect 47696 49010 47730 49066
rect 47696 48790 47730 48852
rect 48148 48790 48182 49066
rect 47696 48756 48182 48790
rect 52686 49382 53172 49416
rect 52686 49320 52720 49382
rect 52686 49106 52720 49162
rect 53138 49106 53172 49382
rect 52686 49066 53172 49106
rect 52686 49010 52720 49066
rect 52686 48790 52720 48852
rect 53138 48790 53172 49066
rect 52686 48756 53172 48790
rect 57676 49382 58162 49416
rect 57676 49320 57710 49382
rect 57676 49106 57710 49162
rect 58128 49106 58162 49382
rect 57676 49066 58162 49106
rect 57676 49010 57710 49066
rect 57676 48790 57710 48852
rect 58128 48790 58162 49066
rect 57676 48756 58162 48790
rect 62666 49382 63152 49416
rect 62666 49320 62700 49382
rect 62666 49106 62700 49162
rect 63118 49106 63152 49382
rect 62666 49066 63152 49106
rect 62666 49010 62700 49066
rect 62666 48790 62700 48852
rect 63118 48790 63152 49066
rect 62666 48756 63152 48790
rect 67656 49382 68142 49416
rect 67656 49320 67690 49382
rect 67656 49106 67690 49162
rect 68108 49106 68142 49382
rect 67656 49066 68142 49106
rect 67656 49010 67690 49066
rect 67656 48790 67690 48852
rect 68108 48790 68142 49066
rect 67656 48756 68142 48790
rect 72646 49382 73132 49416
rect 72646 49320 72680 49382
rect 72646 49106 72680 49162
rect 73098 49106 73132 49382
rect 72646 49066 73132 49106
rect 72646 49010 72680 49066
rect 72646 48790 72680 48852
rect 73098 48790 73132 49066
rect 72646 48756 73132 48790
rect 77636 49382 78122 49416
rect 77636 49320 77670 49382
rect 77636 49106 77670 49162
rect 78088 49106 78122 49382
rect 77636 49066 78122 49106
rect 77636 49010 77670 49066
rect 77636 48790 77670 48852
rect 78088 48790 78122 49066
rect 77636 48756 78122 48790
rect 2786 47672 3272 47706
rect 2786 47610 2820 47672
rect 2786 47396 2820 47452
rect 3238 47396 3272 47672
rect 2786 47356 3272 47396
rect 2786 47300 2820 47356
rect 2786 47080 2820 47142
rect 3238 47080 3272 47356
rect 2786 47046 3272 47080
rect 7776 47672 8262 47706
rect 7776 47610 7810 47672
rect 7776 47396 7810 47452
rect 8228 47396 8262 47672
rect 7776 47356 8262 47396
rect 7776 47300 7810 47356
rect 7776 47080 7810 47142
rect 8228 47080 8262 47356
rect 7776 47046 8262 47080
rect 12766 47672 13252 47706
rect 12766 47610 12800 47672
rect 12766 47396 12800 47452
rect 13218 47396 13252 47672
rect 12766 47356 13252 47396
rect 12766 47300 12800 47356
rect 12766 47080 12800 47142
rect 13218 47080 13252 47356
rect 12766 47046 13252 47080
rect 17756 47672 18242 47706
rect 17756 47610 17790 47672
rect 17756 47396 17790 47452
rect 18208 47396 18242 47672
rect 17756 47356 18242 47396
rect 17756 47300 17790 47356
rect 17756 47080 17790 47142
rect 18208 47080 18242 47356
rect 17756 47046 18242 47080
rect 22746 47672 23232 47706
rect 22746 47610 22780 47672
rect 22746 47396 22780 47452
rect 23198 47396 23232 47672
rect 22746 47356 23232 47396
rect 22746 47300 22780 47356
rect 22746 47080 22780 47142
rect 23198 47080 23232 47356
rect 22746 47046 23232 47080
rect 27736 47672 28222 47706
rect 27736 47610 27770 47672
rect 27736 47396 27770 47452
rect 28188 47396 28222 47672
rect 27736 47356 28222 47396
rect 27736 47300 27770 47356
rect 27736 47080 27770 47142
rect 28188 47080 28222 47356
rect 27736 47046 28222 47080
rect 32726 47672 33212 47706
rect 32726 47610 32760 47672
rect 32726 47396 32760 47452
rect 33178 47396 33212 47672
rect 32726 47356 33212 47396
rect 32726 47300 32760 47356
rect 32726 47080 32760 47142
rect 33178 47080 33212 47356
rect 32726 47046 33212 47080
rect 37716 47672 38202 47706
rect 37716 47610 37750 47672
rect 37716 47396 37750 47452
rect 38168 47396 38202 47672
rect 37716 47356 38202 47396
rect 37716 47300 37750 47356
rect 37716 47080 37750 47142
rect 38168 47080 38202 47356
rect 37716 47046 38202 47080
rect 42706 47672 43192 47706
rect 42706 47610 42740 47672
rect 42706 47396 42740 47452
rect 43158 47396 43192 47672
rect 42706 47356 43192 47396
rect 42706 47300 42740 47356
rect 42706 47080 42740 47142
rect 43158 47080 43192 47356
rect 42706 47046 43192 47080
rect 47696 47672 48182 47706
rect 47696 47610 47730 47672
rect 47696 47396 47730 47452
rect 48148 47396 48182 47672
rect 47696 47356 48182 47396
rect 47696 47300 47730 47356
rect 47696 47080 47730 47142
rect 48148 47080 48182 47356
rect 47696 47046 48182 47080
rect 52686 47672 53172 47706
rect 52686 47610 52720 47672
rect 52686 47396 52720 47452
rect 53138 47396 53172 47672
rect 52686 47356 53172 47396
rect 52686 47300 52720 47356
rect 52686 47080 52720 47142
rect 53138 47080 53172 47356
rect 52686 47046 53172 47080
rect 57676 47672 58162 47706
rect 57676 47610 57710 47672
rect 57676 47396 57710 47452
rect 58128 47396 58162 47672
rect 57676 47356 58162 47396
rect 57676 47300 57710 47356
rect 57676 47080 57710 47142
rect 58128 47080 58162 47356
rect 57676 47046 58162 47080
rect 62666 47672 63152 47706
rect 62666 47610 62700 47672
rect 62666 47396 62700 47452
rect 63118 47396 63152 47672
rect 62666 47356 63152 47396
rect 62666 47300 62700 47356
rect 62666 47080 62700 47142
rect 63118 47080 63152 47356
rect 62666 47046 63152 47080
rect 67656 47672 68142 47706
rect 67656 47610 67690 47672
rect 67656 47396 67690 47452
rect 68108 47396 68142 47672
rect 67656 47356 68142 47396
rect 67656 47300 67690 47356
rect 67656 47080 67690 47142
rect 68108 47080 68142 47356
rect 67656 47046 68142 47080
rect 72646 47672 73132 47706
rect 72646 47610 72680 47672
rect 72646 47396 72680 47452
rect 73098 47396 73132 47672
rect 72646 47356 73132 47396
rect 72646 47300 72680 47356
rect 72646 47080 72680 47142
rect 73098 47080 73132 47356
rect 72646 47046 73132 47080
rect 77636 47672 78122 47706
rect 77636 47610 77670 47672
rect 77636 47396 77670 47452
rect 78088 47396 78122 47672
rect 77636 47356 78122 47396
rect 77636 47300 77670 47356
rect 77636 47080 77670 47142
rect 78088 47080 78122 47356
rect 77636 47046 78122 47080
rect 2786 45962 3272 45996
rect 2786 45900 2820 45962
rect 2786 45686 2820 45742
rect 3238 45686 3272 45962
rect 2786 45646 3272 45686
rect 2786 45590 2820 45646
rect 2786 45370 2820 45432
rect 3238 45370 3272 45646
rect 2786 45336 3272 45370
rect 7776 45962 8262 45996
rect 7776 45900 7810 45962
rect 7776 45686 7810 45742
rect 8228 45686 8262 45962
rect 7776 45646 8262 45686
rect 7776 45590 7810 45646
rect 7776 45370 7810 45432
rect 8228 45370 8262 45646
rect 7776 45336 8262 45370
rect 12766 45962 13252 45996
rect 12766 45900 12800 45962
rect 12766 45686 12800 45742
rect 13218 45686 13252 45962
rect 12766 45646 13252 45686
rect 12766 45590 12800 45646
rect 12766 45370 12800 45432
rect 13218 45370 13252 45646
rect 12766 45336 13252 45370
rect 17756 45962 18242 45996
rect 17756 45900 17790 45962
rect 17756 45686 17790 45742
rect 18208 45686 18242 45962
rect 17756 45646 18242 45686
rect 17756 45590 17790 45646
rect 17756 45370 17790 45432
rect 18208 45370 18242 45646
rect 17756 45336 18242 45370
rect 22746 45962 23232 45996
rect 22746 45900 22780 45962
rect 22746 45686 22780 45742
rect 23198 45686 23232 45962
rect 22746 45646 23232 45686
rect 22746 45590 22780 45646
rect 22746 45370 22780 45432
rect 23198 45370 23232 45646
rect 22746 45336 23232 45370
rect 27736 45962 28222 45996
rect 27736 45900 27770 45962
rect 27736 45686 27770 45742
rect 28188 45686 28222 45962
rect 27736 45646 28222 45686
rect 27736 45590 27770 45646
rect 27736 45370 27770 45432
rect 28188 45370 28222 45646
rect 27736 45336 28222 45370
rect 32726 45962 33212 45996
rect 32726 45900 32760 45962
rect 32726 45686 32760 45742
rect 33178 45686 33212 45962
rect 32726 45646 33212 45686
rect 32726 45590 32760 45646
rect 32726 45370 32760 45432
rect 33178 45370 33212 45646
rect 32726 45336 33212 45370
rect 37716 45962 38202 45996
rect 37716 45900 37750 45962
rect 37716 45686 37750 45742
rect 38168 45686 38202 45962
rect 37716 45646 38202 45686
rect 37716 45590 37750 45646
rect 37716 45370 37750 45432
rect 38168 45370 38202 45646
rect 37716 45336 38202 45370
rect 42706 45962 43192 45996
rect 42706 45900 42740 45962
rect 42706 45686 42740 45742
rect 43158 45686 43192 45962
rect 42706 45646 43192 45686
rect 42706 45590 42740 45646
rect 42706 45370 42740 45432
rect 43158 45370 43192 45646
rect 42706 45336 43192 45370
rect 47696 45962 48182 45996
rect 47696 45900 47730 45962
rect 47696 45686 47730 45742
rect 48148 45686 48182 45962
rect 47696 45646 48182 45686
rect 47696 45590 47730 45646
rect 47696 45370 47730 45432
rect 48148 45370 48182 45646
rect 47696 45336 48182 45370
rect 52686 45962 53172 45996
rect 52686 45900 52720 45962
rect 52686 45686 52720 45742
rect 53138 45686 53172 45962
rect 52686 45646 53172 45686
rect 52686 45590 52720 45646
rect 52686 45370 52720 45432
rect 53138 45370 53172 45646
rect 52686 45336 53172 45370
rect 57676 45962 58162 45996
rect 57676 45900 57710 45962
rect 57676 45686 57710 45742
rect 58128 45686 58162 45962
rect 57676 45646 58162 45686
rect 57676 45590 57710 45646
rect 57676 45370 57710 45432
rect 58128 45370 58162 45646
rect 57676 45336 58162 45370
rect 62666 45962 63152 45996
rect 62666 45900 62700 45962
rect 62666 45686 62700 45742
rect 63118 45686 63152 45962
rect 62666 45646 63152 45686
rect 62666 45590 62700 45646
rect 62666 45370 62700 45432
rect 63118 45370 63152 45646
rect 62666 45336 63152 45370
rect 67656 45962 68142 45996
rect 67656 45900 67690 45962
rect 67656 45686 67690 45742
rect 68108 45686 68142 45962
rect 67656 45646 68142 45686
rect 67656 45590 67690 45646
rect 67656 45370 67690 45432
rect 68108 45370 68142 45646
rect 67656 45336 68142 45370
rect 72646 45962 73132 45996
rect 72646 45900 72680 45962
rect 72646 45686 72680 45742
rect 73098 45686 73132 45962
rect 72646 45646 73132 45686
rect 72646 45590 72680 45646
rect 72646 45370 72680 45432
rect 73098 45370 73132 45646
rect 72646 45336 73132 45370
rect 77636 45962 78122 45996
rect 77636 45900 77670 45962
rect 77636 45686 77670 45742
rect 78088 45686 78122 45962
rect 77636 45646 78122 45686
rect 77636 45590 77670 45646
rect 77636 45370 77670 45432
rect 78088 45370 78122 45646
rect 77636 45336 78122 45370
rect 2786 44252 3272 44286
rect 2786 44190 2820 44252
rect 2786 43976 2820 44032
rect 3238 43976 3272 44252
rect 2786 43936 3272 43976
rect 2786 43880 2820 43936
rect 2786 43660 2820 43722
rect 3238 43660 3272 43936
rect 2786 43626 3272 43660
rect 7776 44252 8262 44286
rect 7776 44190 7810 44252
rect 7776 43976 7810 44032
rect 8228 43976 8262 44252
rect 7776 43936 8262 43976
rect 7776 43880 7810 43936
rect 7776 43660 7810 43722
rect 8228 43660 8262 43936
rect 7776 43626 8262 43660
rect 12766 44252 13252 44286
rect 12766 44190 12800 44252
rect 12766 43976 12800 44032
rect 13218 43976 13252 44252
rect 12766 43936 13252 43976
rect 12766 43880 12800 43936
rect 12766 43660 12800 43722
rect 13218 43660 13252 43936
rect 12766 43626 13252 43660
rect 17756 44252 18242 44286
rect 17756 44190 17790 44252
rect 17756 43976 17790 44032
rect 18208 43976 18242 44252
rect 17756 43936 18242 43976
rect 17756 43880 17790 43936
rect 17756 43660 17790 43722
rect 18208 43660 18242 43936
rect 17756 43626 18242 43660
rect 22746 44252 23232 44286
rect 22746 44190 22780 44252
rect 22746 43976 22780 44032
rect 23198 43976 23232 44252
rect 22746 43936 23232 43976
rect 22746 43880 22780 43936
rect 22746 43660 22780 43722
rect 23198 43660 23232 43936
rect 22746 43626 23232 43660
rect 27736 44252 28222 44286
rect 27736 44190 27770 44252
rect 27736 43976 27770 44032
rect 28188 43976 28222 44252
rect 27736 43936 28222 43976
rect 27736 43880 27770 43936
rect 27736 43660 27770 43722
rect 28188 43660 28222 43936
rect 27736 43626 28222 43660
rect 32726 44252 33212 44286
rect 32726 44190 32760 44252
rect 32726 43976 32760 44032
rect 33178 43976 33212 44252
rect 32726 43936 33212 43976
rect 32726 43880 32760 43936
rect 32726 43660 32760 43722
rect 33178 43660 33212 43936
rect 32726 43626 33212 43660
rect 37716 44252 38202 44286
rect 37716 44190 37750 44252
rect 37716 43976 37750 44032
rect 38168 43976 38202 44252
rect 37716 43936 38202 43976
rect 37716 43880 37750 43936
rect 37716 43660 37750 43722
rect 38168 43660 38202 43936
rect 37716 43626 38202 43660
rect 42706 44252 43192 44286
rect 42706 44190 42740 44252
rect 42706 43976 42740 44032
rect 43158 43976 43192 44252
rect 42706 43936 43192 43976
rect 42706 43880 42740 43936
rect 42706 43660 42740 43722
rect 43158 43660 43192 43936
rect 42706 43626 43192 43660
rect 47696 44252 48182 44286
rect 47696 44190 47730 44252
rect 47696 43976 47730 44032
rect 48148 43976 48182 44252
rect 47696 43936 48182 43976
rect 47696 43880 47730 43936
rect 47696 43660 47730 43722
rect 48148 43660 48182 43936
rect 47696 43626 48182 43660
rect 52686 44252 53172 44286
rect 52686 44190 52720 44252
rect 52686 43976 52720 44032
rect 53138 43976 53172 44252
rect 52686 43936 53172 43976
rect 52686 43880 52720 43936
rect 52686 43660 52720 43722
rect 53138 43660 53172 43936
rect 52686 43626 53172 43660
rect 57676 44252 58162 44286
rect 57676 44190 57710 44252
rect 57676 43976 57710 44032
rect 58128 43976 58162 44252
rect 57676 43936 58162 43976
rect 57676 43880 57710 43936
rect 57676 43660 57710 43722
rect 58128 43660 58162 43936
rect 57676 43626 58162 43660
rect 62666 44252 63152 44286
rect 62666 44190 62700 44252
rect 62666 43976 62700 44032
rect 63118 43976 63152 44252
rect 62666 43936 63152 43976
rect 62666 43880 62700 43936
rect 62666 43660 62700 43722
rect 63118 43660 63152 43936
rect 62666 43626 63152 43660
rect 67656 44252 68142 44286
rect 67656 44190 67690 44252
rect 67656 43976 67690 44032
rect 68108 43976 68142 44252
rect 67656 43936 68142 43976
rect 67656 43880 67690 43936
rect 67656 43660 67690 43722
rect 68108 43660 68142 43936
rect 67656 43626 68142 43660
rect 72646 44252 73132 44286
rect 72646 44190 72680 44252
rect 72646 43976 72680 44032
rect 73098 43976 73132 44252
rect 72646 43936 73132 43976
rect 72646 43880 72680 43936
rect 72646 43660 72680 43722
rect 73098 43660 73132 43936
rect 72646 43626 73132 43660
rect 77636 44252 78122 44286
rect 77636 44190 77670 44252
rect 77636 43976 77670 44032
rect 78088 43976 78122 44252
rect 77636 43936 78122 43976
rect 77636 43880 77670 43936
rect 77636 43660 77670 43722
rect 78088 43660 78122 43936
rect 77636 43626 78122 43660
rect 2786 42542 3272 42576
rect 2786 42480 2820 42542
rect 2786 42266 2820 42322
rect 3238 42266 3272 42542
rect 2786 42226 3272 42266
rect 2786 42170 2820 42226
rect 2786 41950 2820 42012
rect 3238 41950 3272 42226
rect 2786 41916 3272 41950
rect 7776 42542 8262 42576
rect 7776 42480 7810 42542
rect 7776 42266 7810 42322
rect 8228 42266 8262 42542
rect 7776 42226 8262 42266
rect 7776 42170 7810 42226
rect 7776 41950 7810 42012
rect 8228 41950 8262 42226
rect 7776 41916 8262 41950
rect 12766 42542 13252 42576
rect 12766 42480 12800 42542
rect 12766 42266 12800 42322
rect 13218 42266 13252 42542
rect 12766 42226 13252 42266
rect 12766 42170 12800 42226
rect 12766 41950 12800 42012
rect 13218 41950 13252 42226
rect 12766 41916 13252 41950
rect 17756 42542 18242 42576
rect 17756 42480 17790 42542
rect 17756 42266 17790 42322
rect 18208 42266 18242 42542
rect 17756 42226 18242 42266
rect 17756 42170 17790 42226
rect 17756 41950 17790 42012
rect 18208 41950 18242 42226
rect 17756 41916 18242 41950
rect 22746 42542 23232 42576
rect 22746 42480 22780 42542
rect 22746 42266 22780 42322
rect 23198 42266 23232 42542
rect 22746 42226 23232 42266
rect 22746 42170 22780 42226
rect 22746 41950 22780 42012
rect 23198 41950 23232 42226
rect 22746 41916 23232 41950
rect 27736 42542 28222 42576
rect 27736 42480 27770 42542
rect 27736 42266 27770 42322
rect 28188 42266 28222 42542
rect 27736 42226 28222 42266
rect 27736 42170 27770 42226
rect 27736 41950 27770 42012
rect 28188 41950 28222 42226
rect 27736 41916 28222 41950
rect 32726 42542 33212 42576
rect 32726 42480 32760 42542
rect 32726 42266 32760 42322
rect 33178 42266 33212 42542
rect 32726 42226 33212 42266
rect 32726 42170 32760 42226
rect 32726 41950 32760 42012
rect 33178 41950 33212 42226
rect 32726 41916 33212 41950
rect 37716 42542 38202 42576
rect 37716 42480 37750 42542
rect 37716 42266 37750 42322
rect 38168 42266 38202 42542
rect 37716 42226 38202 42266
rect 37716 42170 37750 42226
rect 37716 41950 37750 42012
rect 38168 41950 38202 42226
rect 37716 41916 38202 41950
rect 42706 42542 43192 42576
rect 42706 42480 42740 42542
rect 42706 42266 42740 42322
rect 43158 42266 43192 42542
rect 42706 42226 43192 42266
rect 42706 42170 42740 42226
rect 42706 41950 42740 42012
rect 43158 41950 43192 42226
rect 42706 41916 43192 41950
rect 47696 42542 48182 42576
rect 47696 42480 47730 42542
rect 47696 42266 47730 42322
rect 48148 42266 48182 42542
rect 47696 42226 48182 42266
rect 47696 42170 47730 42226
rect 47696 41950 47730 42012
rect 48148 41950 48182 42226
rect 47696 41916 48182 41950
rect 52686 42542 53172 42576
rect 52686 42480 52720 42542
rect 52686 42266 52720 42322
rect 53138 42266 53172 42542
rect 52686 42226 53172 42266
rect 52686 42170 52720 42226
rect 52686 41950 52720 42012
rect 53138 41950 53172 42226
rect 52686 41916 53172 41950
rect 57676 42542 58162 42576
rect 57676 42480 57710 42542
rect 57676 42266 57710 42322
rect 58128 42266 58162 42542
rect 57676 42226 58162 42266
rect 57676 42170 57710 42226
rect 57676 41950 57710 42012
rect 58128 41950 58162 42226
rect 57676 41916 58162 41950
rect 62666 42542 63152 42576
rect 62666 42480 62700 42542
rect 62666 42266 62700 42322
rect 63118 42266 63152 42542
rect 62666 42226 63152 42266
rect 62666 42170 62700 42226
rect 62666 41950 62700 42012
rect 63118 41950 63152 42226
rect 62666 41916 63152 41950
rect 67656 42542 68142 42576
rect 67656 42480 67690 42542
rect 67656 42266 67690 42322
rect 68108 42266 68142 42542
rect 67656 42226 68142 42266
rect 67656 42170 67690 42226
rect 67656 41950 67690 42012
rect 68108 41950 68142 42226
rect 67656 41916 68142 41950
rect 72646 42542 73132 42576
rect 72646 42480 72680 42542
rect 72646 42266 72680 42322
rect 73098 42266 73132 42542
rect 72646 42226 73132 42266
rect 72646 42170 72680 42226
rect 72646 41950 72680 42012
rect 73098 41950 73132 42226
rect 72646 41916 73132 41950
rect 77636 42542 78122 42576
rect 77636 42480 77670 42542
rect 77636 42266 77670 42322
rect 78088 42266 78122 42542
rect 77636 42226 78122 42266
rect 77636 42170 77670 42226
rect 77636 41950 77670 42012
rect 78088 41950 78122 42226
rect 77636 41916 78122 41950
rect 2786 40832 3272 40866
rect 2786 40770 2820 40832
rect 2786 40556 2820 40612
rect 3238 40556 3272 40832
rect 2786 40516 3272 40556
rect 2786 40460 2820 40516
rect 2786 40240 2820 40302
rect 3238 40240 3272 40516
rect 2786 40206 3272 40240
rect 7776 40832 8262 40866
rect 7776 40770 7810 40832
rect 7776 40556 7810 40612
rect 8228 40556 8262 40832
rect 7776 40516 8262 40556
rect 7776 40460 7810 40516
rect 7776 40240 7810 40302
rect 8228 40240 8262 40516
rect 7776 40206 8262 40240
rect 12766 40832 13252 40866
rect 12766 40770 12800 40832
rect 12766 40556 12800 40612
rect 13218 40556 13252 40832
rect 12766 40516 13252 40556
rect 12766 40460 12800 40516
rect 12766 40240 12800 40302
rect 13218 40240 13252 40516
rect 12766 40206 13252 40240
rect 17756 40832 18242 40866
rect 17756 40770 17790 40832
rect 17756 40556 17790 40612
rect 18208 40556 18242 40832
rect 17756 40516 18242 40556
rect 17756 40460 17790 40516
rect 17756 40240 17790 40302
rect 18208 40240 18242 40516
rect 17756 40206 18242 40240
rect 22746 40832 23232 40866
rect 22746 40770 22780 40832
rect 22746 40556 22780 40612
rect 23198 40556 23232 40832
rect 22746 40516 23232 40556
rect 22746 40460 22780 40516
rect 22746 40240 22780 40302
rect 23198 40240 23232 40516
rect 22746 40206 23232 40240
rect 27736 40832 28222 40866
rect 27736 40770 27770 40832
rect 27736 40556 27770 40612
rect 28188 40556 28222 40832
rect 27736 40516 28222 40556
rect 27736 40460 27770 40516
rect 27736 40240 27770 40302
rect 28188 40240 28222 40516
rect 27736 40206 28222 40240
rect 32726 40832 33212 40866
rect 32726 40770 32760 40832
rect 32726 40556 32760 40612
rect 33178 40556 33212 40832
rect 32726 40516 33212 40556
rect 32726 40460 32760 40516
rect 32726 40240 32760 40302
rect 33178 40240 33212 40516
rect 32726 40206 33212 40240
rect 37716 40832 38202 40866
rect 37716 40770 37750 40832
rect 37716 40556 37750 40612
rect 38168 40556 38202 40832
rect 37716 40516 38202 40556
rect 37716 40460 37750 40516
rect 37716 40240 37750 40302
rect 38168 40240 38202 40516
rect 37716 40206 38202 40240
rect 42706 40832 43192 40866
rect 42706 40770 42740 40832
rect 42706 40556 42740 40612
rect 43158 40556 43192 40832
rect 42706 40516 43192 40556
rect 42706 40460 42740 40516
rect 42706 40240 42740 40302
rect 43158 40240 43192 40516
rect 42706 40206 43192 40240
rect 47696 40832 48182 40866
rect 47696 40770 47730 40832
rect 47696 40556 47730 40612
rect 48148 40556 48182 40832
rect 47696 40516 48182 40556
rect 47696 40460 47730 40516
rect 47696 40240 47730 40302
rect 48148 40240 48182 40516
rect 47696 40206 48182 40240
rect 52686 40832 53172 40866
rect 52686 40770 52720 40832
rect 52686 40556 52720 40612
rect 53138 40556 53172 40832
rect 52686 40516 53172 40556
rect 52686 40460 52720 40516
rect 52686 40240 52720 40302
rect 53138 40240 53172 40516
rect 52686 40206 53172 40240
rect 57676 40832 58162 40866
rect 57676 40770 57710 40832
rect 57676 40556 57710 40612
rect 58128 40556 58162 40832
rect 57676 40516 58162 40556
rect 57676 40460 57710 40516
rect 57676 40240 57710 40302
rect 58128 40240 58162 40516
rect 57676 40206 58162 40240
rect 62666 40832 63152 40866
rect 62666 40770 62700 40832
rect 62666 40556 62700 40612
rect 63118 40556 63152 40832
rect 62666 40516 63152 40556
rect 62666 40460 62700 40516
rect 62666 40240 62700 40302
rect 63118 40240 63152 40516
rect 62666 40206 63152 40240
rect 67656 40832 68142 40866
rect 67656 40770 67690 40832
rect 67656 40556 67690 40612
rect 68108 40556 68142 40832
rect 67656 40516 68142 40556
rect 67656 40460 67690 40516
rect 67656 40240 67690 40302
rect 68108 40240 68142 40516
rect 67656 40206 68142 40240
rect 72646 40832 73132 40866
rect 72646 40770 72680 40832
rect 72646 40556 72680 40612
rect 73098 40556 73132 40832
rect 72646 40516 73132 40556
rect 72646 40460 72680 40516
rect 72646 40240 72680 40302
rect 73098 40240 73132 40516
rect 72646 40206 73132 40240
rect 77636 40832 78122 40866
rect 77636 40770 77670 40832
rect 77636 40556 77670 40612
rect 78088 40556 78122 40832
rect 77636 40516 78122 40556
rect 77636 40460 77670 40516
rect 77636 40240 77670 40302
rect 78088 40240 78122 40516
rect 77636 40206 78122 40240
<< nsubdiff >>
rect 3346 66482 3842 66516
rect 3346 66206 3380 66482
rect 3808 66420 3842 66482
rect 3808 66206 3842 66262
rect 3346 66166 3842 66206
rect 3346 65890 3380 66166
rect 3808 66110 3842 66166
rect 3808 65890 3842 65952
rect 3346 65856 3842 65890
rect 8336 66482 8832 66516
rect 8336 66206 8370 66482
rect 8798 66420 8832 66482
rect 8798 66206 8832 66262
rect 8336 66166 8832 66206
rect 8336 65890 8370 66166
rect 8798 66110 8832 66166
rect 8798 65890 8832 65952
rect 8336 65856 8832 65890
rect 13326 66482 13822 66516
rect 13326 66206 13360 66482
rect 13788 66420 13822 66482
rect 13788 66206 13822 66262
rect 13326 66166 13822 66206
rect 13326 65890 13360 66166
rect 13788 66110 13822 66166
rect 13788 65890 13822 65952
rect 13326 65856 13822 65890
rect 18316 66482 18812 66516
rect 18316 66206 18350 66482
rect 18778 66420 18812 66482
rect 18778 66206 18812 66262
rect 18316 66166 18812 66206
rect 18316 65890 18350 66166
rect 18778 66110 18812 66166
rect 18778 65890 18812 65952
rect 18316 65856 18812 65890
rect 23306 66482 23802 66516
rect 23306 66206 23340 66482
rect 23768 66420 23802 66482
rect 23768 66206 23802 66262
rect 23306 66166 23802 66206
rect 23306 65890 23340 66166
rect 23768 66110 23802 66166
rect 23768 65890 23802 65952
rect 23306 65856 23802 65890
rect 28296 66482 28792 66516
rect 28296 66206 28330 66482
rect 28758 66420 28792 66482
rect 28758 66206 28792 66262
rect 28296 66166 28792 66206
rect 28296 65890 28330 66166
rect 28758 66110 28792 66166
rect 28758 65890 28792 65952
rect 28296 65856 28792 65890
rect 33286 66482 33782 66516
rect 33286 66206 33320 66482
rect 33748 66420 33782 66482
rect 33748 66206 33782 66262
rect 33286 66166 33782 66206
rect 33286 65890 33320 66166
rect 33748 66110 33782 66166
rect 33748 65890 33782 65952
rect 33286 65856 33782 65890
rect 38276 66482 38772 66516
rect 38276 66206 38310 66482
rect 38738 66420 38772 66482
rect 38738 66206 38772 66262
rect 38276 66166 38772 66206
rect 38276 65890 38310 66166
rect 38738 66110 38772 66166
rect 38738 65890 38772 65952
rect 38276 65856 38772 65890
rect 43266 66482 43762 66516
rect 43266 66206 43300 66482
rect 43728 66420 43762 66482
rect 43728 66206 43762 66262
rect 43266 66166 43762 66206
rect 43266 65890 43300 66166
rect 43728 66110 43762 66166
rect 43728 65890 43762 65952
rect 43266 65856 43762 65890
rect 48256 66482 48752 66516
rect 48256 66206 48290 66482
rect 48718 66420 48752 66482
rect 48718 66206 48752 66262
rect 48256 66166 48752 66206
rect 48256 65890 48290 66166
rect 48718 66110 48752 66166
rect 48718 65890 48752 65952
rect 48256 65856 48752 65890
rect 53246 66482 53742 66516
rect 53246 66206 53280 66482
rect 53708 66420 53742 66482
rect 53708 66206 53742 66262
rect 53246 66166 53742 66206
rect 53246 65890 53280 66166
rect 53708 66110 53742 66166
rect 53708 65890 53742 65952
rect 53246 65856 53742 65890
rect 58236 66482 58732 66516
rect 58236 66206 58270 66482
rect 58698 66420 58732 66482
rect 58698 66206 58732 66262
rect 58236 66166 58732 66206
rect 58236 65890 58270 66166
rect 58698 66110 58732 66166
rect 58698 65890 58732 65952
rect 58236 65856 58732 65890
rect 63226 66482 63722 66516
rect 63226 66206 63260 66482
rect 63688 66420 63722 66482
rect 63688 66206 63722 66262
rect 63226 66166 63722 66206
rect 63226 65890 63260 66166
rect 63688 66110 63722 66166
rect 63688 65890 63722 65952
rect 63226 65856 63722 65890
rect 68216 66482 68712 66516
rect 68216 66206 68250 66482
rect 68678 66420 68712 66482
rect 68678 66206 68712 66262
rect 68216 66166 68712 66206
rect 68216 65890 68250 66166
rect 68678 66110 68712 66166
rect 68678 65890 68712 65952
rect 68216 65856 68712 65890
rect 73206 66482 73702 66516
rect 73206 66206 73240 66482
rect 73668 66420 73702 66482
rect 73668 66206 73702 66262
rect 73206 66166 73702 66206
rect 73206 65890 73240 66166
rect 73668 66110 73702 66166
rect 73668 65890 73702 65952
rect 73206 65856 73702 65890
rect 78196 66482 78692 66516
rect 78196 66206 78230 66482
rect 78658 66420 78692 66482
rect 78658 66206 78692 66262
rect 78196 66166 78692 66206
rect 78196 65890 78230 66166
rect 78658 66110 78692 66166
rect 78658 65890 78692 65952
rect 78196 65856 78692 65890
rect 3346 64772 3842 64806
rect 3346 64496 3380 64772
rect 3808 64710 3842 64772
rect 3808 64496 3842 64552
rect 3346 64456 3842 64496
rect 3346 64180 3380 64456
rect 3808 64400 3842 64456
rect 3808 64180 3842 64242
rect 3346 64146 3842 64180
rect 8336 64772 8832 64806
rect 8336 64496 8370 64772
rect 8798 64710 8832 64772
rect 8798 64496 8832 64552
rect 8336 64456 8832 64496
rect 8336 64180 8370 64456
rect 8798 64400 8832 64456
rect 8798 64180 8832 64242
rect 8336 64146 8832 64180
rect 13326 64772 13822 64806
rect 13326 64496 13360 64772
rect 13788 64710 13822 64772
rect 13788 64496 13822 64552
rect 13326 64456 13822 64496
rect 13326 64180 13360 64456
rect 13788 64400 13822 64456
rect 13788 64180 13822 64242
rect 13326 64146 13822 64180
rect 18316 64772 18812 64806
rect 18316 64496 18350 64772
rect 18778 64710 18812 64772
rect 18778 64496 18812 64552
rect 18316 64456 18812 64496
rect 18316 64180 18350 64456
rect 18778 64400 18812 64456
rect 18778 64180 18812 64242
rect 18316 64146 18812 64180
rect 23306 64772 23802 64806
rect 23306 64496 23340 64772
rect 23768 64710 23802 64772
rect 23768 64496 23802 64552
rect 23306 64456 23802 64496
rect 23306 64180 23340 64456
rect 23768 64400 23802 64456
rect 23768 64180 23802 64242
rect 23306 64146 23802 64180
rect 28296 64772 28792 64806
rect 28296 64496 28330 64772
rect 28758 64710 28792 64772
rect 28758 64496 28792 64552
rect 28296 64456 28792 64496
rect 28296 64180 28330 64456
rect 28758 64400 28792 64456
rect 28758 64180 28792 64242
rect 28296 64146 28792 64180
rect 33286 64772 33782 64806
rect 33286 64496 33320 64772
rect 33748 64710 33782 64772
rect 33748 64496 33782 64552
rect 33286 64456 33782 64496
rect 33286 64180 33320 64456
rect 33748 64400 33782 64456
rect 33748 64180 33782 64242
rect 33286 64146 33782 64180
rect 38276 64772 38772 64806
rect 38276 64496 38310 64772
rect 38738 64710 38772 64772
rect 38738 64496 38772 64552
rect 38276 64456 38772 64496
rect 38276 64180 38310 64456
rect 38738 64400 38772 64456
rect 38738 64180 38772 64242
rect 38276 64146 38772 64180
rect 43266 64772 43762 64806
rect 43266 64496 43300 64772
rect 43728 64710 43762 64772
rect 43728 64496 43762 64552
rect 43266 64456 43762 64496
rect 43266 64180 43300 64456
rect 43728 64400 43762 64456
rect 43728 64180 43762 64242
rect 43266 64146 43762 64180
rect 48256 64772 48752 64806
rect 48256 64496 48290 64772
rect 48718 64710 48752 64772
rect 48718 64496 48752 64552
rect 48256 64456 48752 64496
rect 48256 64180 48290 64456
rect 48718 64400 48752 64456
rect 48718 64180 48752 64242
rect 48256 64146 48752 64180
rect 53246 64772 53742 64806
rect 53246 64496 53280 64772
rect 53708 64710 53742 64772
rect 53708 64496 53742 64552
rect 53246 64456 53742 64496
rect 53246 64180 53280 64456
rect 53708 64400 53742 64456
rect 53708 64180 53742 64242
rect 53246 64146 53742 64180
rect 58236 64772 58732 64806
rect 58236 64496 58270 64772
rect 58698 64710 58732 64772
rect 58698 64496 58732 64552
rect 58236 64456 58732 64496
rect 58236 64180 58270 64456
rect 58698 64400 58732 64456
rect 58698 64180 58732 64242
rect 58236 64146 58732 64180
rect 63226 64772 63722 64806
rect 63226 64496 63260 64772
rect 63688 64710 63722 64772
rect 63688 64496 63722 64552
rect 63226 64456 63722 64496
rect 63226 64180 63260 64456
rect 63688 64400 63722 64456
rect 63688 64180 63722 64242
rect 63226 64146 63722 64180
rect 68216 64772 68712 64806
rect 68216 64496 68250 64772
rect 68678 64710 68712 64772
rect 68678 64496 68712 64552
rect 68216 64456 68712 64496
rect 68216 64180 68250 64456
rect 68678 64400 68712 64456
rect 68678 64180 68712 64242
rect 68216 64146 68712 64180
rect 73206 64772 73702 64806
rect 73206 64496 73240 64772
rect 73668 64710 73702 64772
rect 73668 64496 73702 64552
rect 73206 64456 73702 64496
rect 73206 64180 73240 64456
rect 73668 64400 73702 64456
rect 73668 64180 73702 64242
rect 73206 64146 73702 64180
rect 78196 64772 78692 64806
rect 78196 64496 78230 64772
rect 78658 64710 78692 64772
rect 78658 64496 78692 64552
rect 78196 64456 78692 64496
rect 78196 64180 78230 64456
rect 78658 64400 78692 64456
rect 78658 64180 78692 64242
rect 78196 64146 78692 64180
rect 3346 63062 3842 63096
rect 3346 62786 3380 63062
rect 3808 63000 3842 63062
rect 3808 62786 3842 62842
rect 3346 62746 3842 62786
rect 3346 62470 3380 62746
rect 3808 62690 3842 62746
rect 3808 62470 3842 62532
rect 3346 62436 3842 62470
rect 8336 63062 8832 63096
rect 8336 62786 8370 63062
rect 8798 63000 8832 63062
rect 8798 62786 8832 62842
rect 8336 62746 8832 62786
rect 8336 62470 8370 62746
rect 8798 62690 8832 62746
rect 8798 62470 8832 62532
rect 8336 62436 8832 62470
rect 13326 63062 13822 63096
rect 13326 62786 13360 63062
rect 13788 63000 13822 63062
rect 13788 62786 13822 62842
rect 13326 62746 13822 62786
rect 13326 62470 13360 62746
rect 13788 62690 13822 62746
rect 13788 62470 13822 62532
rect 13326 62436 13822 62470
rect 18316 63062 18812 63096
rect 18316 62786 18350 63062
rect 18778 63000 18812 63062
rect 18778 62786 18812 62842
rect 18316 62746 18812 62786
rect 18316 62470 18350 62746
rect 18778 62690 18812 62746
rect 18778 62470 18812 62532
rect 18316 62436 18812 62470
rect 23306 63062 23802 63096
rect 23306 62786 23340 63062
rect 23768 63000 23802 63062
rect 23768 62786 23802 62842
rect 23306 62746 23802 62786
rect 23306 62470 23340 62746
rect 23768 62690 23802 62746
rect 23768 62470 23802 62532
rect 23306 62436 23802 62470
rect 28296 63062 28792 63096
rect 28296 62786 28330 63062
rect 28758 63000 28792 63062
rect 28758 62786 28792 62842
rect 28296 62746 28792 62786
rect 28296 62470 28330 62746
rect 28758 62690 28792 62746
rect 28758 62470 28792 62532
rect 28296 62436 28792 62470
rect 33286 63062 33782 63096
rect 33286 62786 33320 63062
rect 33748 63000 33782 63062
rect 33748 62786 33782 62842
rect 33286 62746 33782 62786
rect 33286 62470 33320 62746
rect 33748 62690 33782 62746
rect 33748 62470 33782 62532
rect 33286 62436 33782 62470
rect 38276 63062 38772 63096
rect 38276 62786 38310 63062
rect 38738 63000 38772 63062
rect 38738 62786 38772 62842
rect 38276 62746 38772 62786
rect 38276 62470 38310 62746
rect 38738 62690 38772 62746
rect 38738 62470 38772 62532
rect 38276 62436 38772 62470
rect 43266 63062 43762 63096
rect 43266 62786 43300 63062
rect 43728 63000 43762 63062
rect 43728 62786 43762 62842
rect 43266 62746 43762 62786
rect 43266 62470 43300 62746
rect 43728 62690 43762 62746
rect 43728 62470 43762 62532
rect 43266 62436 43762 62470
rect 48256 63062 48752 63096
rect 48256 62786 48290 63062
rect 48718 63000 48752 63062
rect 48718 62786 48752 62842
rect 48256 62746 48752 62786
rect 48256 62470 48290 62746
rect 48718 62690 48752 62746
rect 48718 62470 48752 62532
rect 48256 62436 48752 62470
rect 53246 63062 53742 63096
rect 53246 62786 53280 63062
rect 53708 63000 53742 63062
rect 53708 62786 53742 62842
rect 53246 62746 53742 62786
rect 53246 62470 53280 62746
rect 53708 62690 53742 62746
rect 53708 62470 53742 62532
rect 53246 62436 53742 62470
rect 58236 63062 58732 63096
rect 58236 62786 58270 63062
rect 58698 63000 58732 63062
rect 58698 62786 58732 62842
rect 58236 62746 58732 62786
rect 58236 62470 58270 62746
rect 58698 62690 58732 62746
rect 58698 62470 58732 62532
rect 58236 62436 58732 62470
rect 63226 63062 63722 63096
rect 63226 62786 63260 63062
rect 63688 63000 63722 63062
rect 63688 62786 63722 62842
rect 63226 62746 63722 62786
rect 63226 62470 63260 62746
rect 63688 62690 63722 62746
rect 63688 62470 63722 62532
rect 63226 62436 63722 62470
rect 68216 63062 68712 63096
rect 68216 62786 68250 63062
rect 68678 63000 68712 63062
rect 68678 62786 68712 62842
rect 68216 62746 68712 62786
rect 68216 62470 68250 62746
rect 68678 62690 68712 62746
rect 68678 62470 68712 62532
rect 68216 62436 68712 62470
rect 73206 63062 73702 63096
rect 73206 62786 73240 63062
rect 73668 63000 73702 63062
rect 73668 62786 73702 62842
rect 73206 62746 73702 62786
rect 73206 62470 73240 62746
rect 73668 62690 73702 62746
rect 73668 62470 73702 62532
rect 73206 62436 73702 62470
rect 78196 63062 78692 63096
rect 78196 62786 78230 63062
rect 78658 63000 78692 63062
rect 78658 62786 78692 62842
rect 78196 62746 78692 62786
rect 78196 62470 78230 62746
rect 78658 62690 78692 62746
rect 78658 62470 78692 62532
rect 78196 62436 78692 62470
rect 3346 61352 3842 61386
rect 3346 61076 3380 61352
rect 3808 61290 3842 61352
rect 3808 61076 3842 61132
rect 3346 61036 3842 61076
rect 3346 60760 3380 61036
rect 3808 60980 3842 61036
rect 3808 60760 3842 60822
rect 3346 60726 3842 60760
rect 8336 61352 8832 61386
rect 8336 61076 8370 61352
rect 8798 61290 8832 61352
rect 8798 61076 8832 61132
rect 8336 61036 8832 61076
rect 8336 60760 8370 61036
rect 8798 60980 8832 61036
rect 8798 60760 8832 60822
rect 8336 60726 8832 60760
rect 13326 61352 13822 61386
rect 13326 61076 13360 61352
rect 13788 61290 13822 61352
rect 13788 61076 13822 61132
rect 13326 61036 13822 61076
rect 13326 60760 13360 61036
rect 13788 60980 13822 61036
rect 13788 60760 13822 60822
rect 13326 60726 13822 60760
rect 18316 61352 18812 61386
rect 18316 61076 18350 61352
rect 18778 61290 18812 61352
rect 18778 61076 18812 61132
rect 18316 61036 18812 61076
rect 18316 60760 18350 61036
rect 18778 60980 18812 61036
rect 18778 60760 18812 60822
rect 18316 60726 18812 60760
rect 23306 61352 23802 61386
rect 23306 61076 23340 61352
rect 23768 61290 23802 61352
rect 23768 61076 23802 61132
rect 23306 61036 23802 61076
rect 23306 60760 23340 61036
rect 23768 60980 23802 61036
rect 23768 60760 23802 60822
rect 23306 60726 23802 60760
rect 28296 61352 28792 61386
rect 28296 61076 28330 61352
rect 28758 61290 28792 61352
rect 28758 61076 28792 61132
rect 28296 61036 28792 61076
rect 28296 60760 28330 61036
rect 28758 60980 28792 61036
rect 28758 60760 28792 60822
rect 28296 60726 28792 60760
rect 33286 61352 33782 61386
rect 33286 61076 33320 61352
rect 33748 61290 33782 61352
rect 33748 61076 33782 61132
rect 33286 61036 33782 61076
rect 33286 60760 33320 61036
rect 33748 60980 33782 61036
rect 33748 60760 33782 60822
rect 33286 60726 33782 60760
rect 38276 61352 38772 61386
rect 38276 61076 38310 61352
rect 38738 61290 38772 61352
rect 38738 61076 38772 61132
rect 38276 61036 38772 61076
rect 38276 60760 38310 61036
rect 38738 60980 38772 61036
rect 38738 60760 38772 60822
rect 38276 60726 38772 60760
rect 43266 61352 43762 61386
rect 43266 61076 43300 61352
rect 43728 61290 43762 61352
rect 43728 61076 43762 61132
rect 43266 61036 43762 61076
rect 43266 60760 43300 61036
rect 43728 60980 43762 61036
rect 43728 60760 43762 60822
rect 43266 60726 43762 60760
rect 48256 61352 48752 61386
rect 48256 61076 48290 61352
rect 48718 61290 48752 61352
rect 48718 61076 48752 61132
rect 48256 61036 48752 61076
rect 48256 60760 48290 61036
rect 48718 60980 48752 61036
rect 48718 60760 48752 60822
rect 48256 60726 48752 60760
rect 53246 61352 53742 61386
rect 53246 61076 53280 61352
rect 53708 61290 53742 61352
rect 53708 61076 53742 61132
rect 53246 61036 53742 61076
rect 53246 60760 53280 61036
rect 53708 60980 53742 61036
rect 53708 60760 53742 60822
rect 53246 60726 53742 60760
rect 58236 61352 58732 61386
rect 58236 61076 58270 61352
rect 58698 61290 58732 61352
rect 58698 61076 58732 61132
rect 58236 61036 58732 61076
rect 58236 60760 58270 61036
rect 58698 60980 58732 61036
rect 58698 60760 58732 60822
rect 58236 60726 58732 60760
rect 63226 61352 63722 61386
rect 63226 61076 63260 61352
rect 63688 61290 63722 61352
rect 63688 61076 63722 61132
rect 63226 61036 63722 61076
rect 63226 60760 63260 61036
rect 63688 60980 63722 61036
rect 63688 60760 63722 60822
rect 63226 60726 63722 60760
rect 68216 61352 68712 61386
rect 68216 61076 68250 61352
rect 68678 61290 68712 61352
rect 68678 61076 68712 61132
rect 68216 61036 68712 61076
rect 68216 60760 68250 61036
rect 68678 60980 68712 61036
rect 68678 60760 68712 60822
rect 68216 60726 68712 60760
rect 73206 61352 73702 61386
rect 73206 61076 73240 61352
rect 73668 61290 73702 61352
rect 73668 61076 73702 61132
rect 73206 61036 73702 61076
rect 73206 60760 73240 61036
rect 73668 60980 73702 61036
rect 73668 60760 73702 60822
rect 73206 60726 73702 60760
rect 78196 61352 78692 61386
rect 78196 61076 78230 61352
rect 78658 61290 78692 61352
rect 78658 61076 78692 61132
rect 78196 61036 78692 61076
rect 78196 60760 78230 61036
rect 78658 60980 78692 61036
rect 78658 60760 78692 60822
rect 78196 60726 78692 60760
rect 3346 59642 3842 59676
rect 3346 59366 3380 59642
rect 3808 59580 3842 59642
rect 3808 59366 3842 59422
rect 3346 59326 3842 59366
rect 3346 59050 3380 59326
rect 3808 59270 3842 59326
rect 3808 59050 3842 59112
rect 3346 59016 3842 59050
rect 8336 59642 8832 59676
rect 8336 59366 8370 59642
rect 8798 59580 8832 59642
rect 8798 59366 8832 59422
rect 8336 59326 8832 59366
rect 8336 59050 8370 59326
rect 8798 59270 8832 59326
rect 8798 59050 8832 59112
rect 8336 59016 8832 59050
rect 13326 59642 13822 59676
rect 13326 59366 13360 59642
rect 13788 59580 13822 59642
rect 13788 59366 13822 59422
rect 13326 59326 13822 59366
rect 13326 59050 13360 59326
rect 13788 59270 13822 59326
rect 13788 59050 13822 59112
rect 13326 59016 13822 59050
rect 18316 59642 18812 59676
rect 18316 59366 18350 59642
rect 18778 59580 18812 59642
rect 18778 59366 18812 59422
rect 18316 59326 18812 59366
rect 18316 59050 18350 59326
rect 18778 59270 18812 59326
rect 18778 59050 18812 59112
rect 18316 59016 18812 59050
rect 23306 59642 23802 59676
rect 23306 59366 23340 59642
rect 23768 59580 23802 59642
rect 23768 59366 23802 59422
rect 23306 59326 23802 59366
rect 23306 59050 23340 59326
rect 23768 59270 23802 59326
rect 23768 59050 23802 59112
rect 23306 59016 23802 59050
rect 28296 59642 28792 59676
rect 28296 59366 28330 59642
rect 28758 59580 28792 59642
rect 28758 59366 28792 59422
rect 28296 59326 28792 59366
rect 28296 59050 28330 59326
rect 28758 59270 28792 59326
rect 28758 59050 28792 59112
rect 28296 59016 28792 59050
rect 33286 59642 33782 59676
rect 33286 59366 33320 59642
rect 33748 59580 33782 59642
rect 33748 59366 33782 59422
rect 33286 59326 33782 59366
rect 33286 59050 33320 59326
rect 33748 59270 33782 59326
rect 33748 59050 33782 59112
rect 33286 59016 33782 59050
rect 38276 59642 38772 59676
rect 38276 59366 38310 59642
rect 38738 59580 38772 59642
rect 38738 59366 38772 59422
rect 38276 59326 38772 59366
rect 38276 59050 38310 59326
rect 38738 59270 38772 59326
rect 38738 59050 38772 59112
rect 38276 59016 38772 59050
rect 43266 59642 43762 59676
rect 43266 59366 43300 59642
rect 43728 59580 43762 59642
rect 43728 59366 43762 59422
rect 43266 59326 43762 59366
rect 43266 59050 43300 59326
rect 43728 59270 43762 59326
rect 43728 59050 43762 59112
rect 43266 59016 43762 59050
rect 48256 59642 48752 59676
rect 48256 59366 48290 59642
rect 48718 59580 48752 59642
rect 48718 59366 48752 59422
rect 48256 59326 48752 59366
rect 48256 59050 48290 59326
rect 48718 59270 48752 59326
rect 48718 59050 48752 59112
rect 48256 59016 48752 59050
rect 53246 59642 53742 59676
rect 53246 59366 53280 59642
rect 53708 59580 53742 59642
rect 53708 59366 53742 59422
rect 53246 59326 53742 59366
rect 53246 59050 53280 59326
rect 53708 59270 53742 59326
rect 53708 59050 53742 59112
rect 53246 59016 53742 59050
rect 58236 59642 58732 59676
rect 58236 59366 58270 59642
rect 58698 59580 58732 59642
rect 58698 59366 58732 59422
rect 58236 59326 58732 59366
rect 58236 59050 58270 59326
rect 58698 59270 58732 59326
rect 58698 59050 58732 59112
rect 58236 59016 58732 59050
rect 63226 59642 63722 59676
rect 63226 59366 63260 59642
rect 63688 59580 63722 59642
rect 63688 59366 63722 59422
rect 63226 59326 63722 59366
rect 63226 59050 63260 59326
rect 63688 59270 63722 59326
rect 63688 59050 63722 59112
rect 63226 59016 63722 59050
rect 68216 59642 68712 59676
rect 68216 59366 68250 59642
rect 68678 59580 68712 59642
rect 68678 59366 68712 59422
rect 68216 59326 68712 59366
rect 68216 59050 68250 59326
rect 68678 59270 68712 59326
rect 68678 59050 68712 59112
rect 68216 59016 68712 59050
rect 73206 59642 73702 59676
rect 73206 59366 73240 59642
rect 73668 59580 73702 59642
rect 73668 59366 73702 59422
rect 73206 59326 73702 59366
rect 73206 59050 73240 59326
rect 73668 59270 73702 59326
rect 73668 59050 73702 59112
rect 73206 59016 73702 59050
rect 78196 59642 78692 59676
rect 78196 59366 78230 59642
rect 78658 59580 78692 59642
rect 78658 59366 78692 59422
rect 78196 59326 78692 59366
rect 78196 59050 78230 59326
rect 78658 59270 78692 59326
rect 78658 59050 78692 59112
rect 78196 59016 78692 59050
rect 3346 57932 3842 57966
rect 3346 57656 3380 57932
rect 3808 57870 3842 57932
rect 3808 57656 3842 57712
rect 3346 57616 3842 57656
rect 3346 57340 3380 57616
rect 3808 57560 3842 57616
rect 3808 57340 3842 57402
rect 3346 57306 3842 57340
rect 8336 57932 8832 57966
rect 8336 57656 8370 57932
rect 8798 57870 8832 57932
rect 8798 57656 8832 57712
rect 8336 57616 8832 57656
rect 8336 57340 8370 57616
rect 8798 57560 8832 57616
rect 8798 57340 8832 57402
rect 8336 57306 8832 57340
rect 13326 57932 13822 57966
rect 13326 57656 13360 57932
rect 13788 57870 13822 57932
rect 13788 57656 13822 57712
rect 13326 57616 13822 57656
rect 13326 57340 13360 57616
rect 13788 57560 13822 57616
rect 13788 57340 13822 57402
rect 13326 57306 13822 57340
rect 18316 57932 18812 57966
rect 18316 57656 18350 57932
rect 18778 57870 18812 57932
rect 18778 57656 18812 57712
rect 18316 57616 18812 57656
rect 18316 57340 18350 57616
rect 18778 57560 18812 57616
rect 18778 57340 18812 57402
rect 18316 57306 18812 57340
rect 23306 57932 23802 57966
rect 23306 57656 23340 57932
rect 23768 57870 23802 57932
rect 23768 57656 23802 57712
rect 23306 57616 23802 57656
rect 23306 57340 23340 57616
rect 23768 57560 23802 57616
rect 23768 57340 23802 57402
rect 23306 57306 23802 57340
rect 28296 57932 28792 57966
rect 28296 57656 28330 57932
rect 28758 57870 28792 57932
rect 28758 57656 28792 57712
rect 28296 57616 28792 57656
rect 28296 57340 28330 57616
rect 28758 57560 28792 57616
rect 28758 57340 28792 57402
rect 28296 57306 28792 57340
rect 33286 57932 33782 57966
rect 33286 57656 33320 57932
rect 33748 57870 33782 57932
rect 33748 57656 33782 57712
rect 33286 57616 33782 57656
rect 33286 57340 33320 57616
rect 33748 57560 33782 57616
rect 33748 57340 33782 57402
rect 33286 57306 33782 57340
rect 38276 57932 38772 57966
rect 38276 57656 38310 57932
rect 38738 57870 38772 57932
rect 38738 57656 38772 57712
rect 38276 57616 38772 57656
rect 38276 57340 38310 57616
rect 38738 57560 38772 57616
rect 38738 57340 38772 57402
rect 38276 57306 38772 57340
rect 43266 57932 43762 57966
rect 43266 57656 43300 57932
rect 43728 57870 43762 57932
rect 43728 57656 43762 57712
rect 43266 57616 43762 57656
rect 43266 57340 43300 57616
rect 43728 57560 43762 57616
rect 43728 57340 43762 57402
rect 43266 57306 43762 57340
rect 48256 57932 48752 57966
rect 48256 57656 48290 57932
rect 48718 57870 48752 57932
rect 48718 57656 48752 57712
rect 48256 57616 48752 57656
rect 48256 57340 48290 57616
rect 48718 57560 48752 57616
rect 48718 57340 48752 57402
rect 48256 57306 48752 57340
rect 53246 57932 53742 57966
rect 53246 57656 53280 57932
rect 53708 57870 53742 57932
rect 53708 57656 53742 57712
rect 53246 57616 53742 57656
rect 53246 57340 53280 57616
rect 53708 57560 53742 57616
rect 53708 57340 53742 57402
rect 53246 57306 53742 57340
rect 58236 57932 58732 57966
rect 58236 57656 58270 57932
rect 58698 57870 58732 57932
rect 58698 57656 58732 57712
rect 58236 57616 58732 57656
rect 58236 57340 58270 57616
rect 58698 57560 58732 57616
rect 58698 57340 58732 57402
rect 58236 57306 58732 57340
rect 63226 57932 63722 57966
rect 63226 57656 63260 57932
rect 63688 57870 63722 57932
rect 63688 57656 63722 57712
rect 63226 57616 63722 57656
rect 63226 57340 63260 57616
rect 63688 57560 63722 57616
rect 63688 57340 63722 57402
rect 63226 57306 63722 57340
rect 68216 57932 68712 57966
rect 68216 57656 68250 57932
rect 68678 57870 68712 57932
rect 68678 57656 68712 57712
rect 68216 57616 68712 57656
rect 68216 57340 68250 57616
rect 68678 57560 68712 57616
rect 68678 57340 68712 57402
rect 68216 57306 68712 57340
rect 73206 57932 73702 57966
rect 73206 57656 73240 57932
rect 73668 57870 73702 57932
rect 73668 57656 73702 57712
rect 73206 57616 73702 57656
rect 73206 57340 73240 57616
rect 73668 57560 73702 57616
rect 73668 57340 73702 57402
rect 73206 57306 73702 57340
rect 78196 57932 78692 57966
rect 78196 57656 78230 57932
rect 78658 57870 78692 57932
rect 78658 57656 78692 57712
rect 78196 57616 78692 57656
rect 78196 57340 78230 57616
rect 78658 57560 78692 57616
rect 78658 57340 78692 57402
rect 78196 57306 78692 57340
rect 3346 56222 3842 56256
rect 3346 55946 3380 56222
rect 3808 56160 3842 56222
rect 3808 55946 3842 56002
rect 3346 55906 3842 55946
rect 3346 55630 3380 55906
rect 3808 55850 3842 55906
rect 3808 55630 3842 55692
rect 3346 55596 3842 55630
rect 8336 56222 8832 56256
rect 8336 55946 8370 56222
rect 8798 56160 8832 56222
rect 8798 55946 8832 56002
rect 8336 55906 8832 55946
rect 8336 55630 8370 55906
rect 8798 55850 8832 55906
rect 8798 55630 8832 55692
rect 8336 55596 8832 55630
rect 13326 56222 13822 56256
rect 13326 55946 13360 56222
rect 13788 56160 13822 56222
rect 13788 55946 13822 56002
rect 13326 55906 13822 55946
rect 13326 55630 13360 55906
rect 13788 55850 13822 55906
rect 13788 55630 13822 55692
rect 13326 55596 13822 55630
rect 18316 56222 18812 56256
rect 18316 55946 18350 56222
rect 18778 56160 18812 56222
rect 18778 55946 18812 56002
rect 18316 55906 18812 55946
rect 18316 55630 18350 55906
rect 18778 55850 18812 55906
rect 18778 55630 18812 55692
rect 18316 55596 18812 55630
rect 23306 56222 23802 56256
rect 23306 55946 23340 56222
rect 23768 56160 23802 56222
rect 23768 55946 23802 56002
rect 23306 55906 23802 55946
rect 23306 55630 23340 55906
rect 23768 55850 23802 55906
rect 23768 55630 23802 55692
rect 23306 55596 23802 55630
rect 28296 56222 28792 56256
rect 28296 55946 28330 56222
rect 28758 56160 28792 56222
rect 28758 55946 28792 56002
rect 28296 55906 28792 55946
rect 28296 55630 28330 55906
rect 28758 55850 28792 55906
rect 28758 55630 28792 55692
rect 28296 55596 28792 55630
rect 33286 56222 33782 56256
rect 33286 55946 33320 56222
rect 33748 56160 33782 56222
rect 33748 55946 33782 56002
rect 33286 55906 33782 55946
rect 33286 55630 33320 55906
rect 33748 55850 33782 55906
rect 33748 55630 33782 55692
rect 33286 55596 33782 55630
rect 38276 56222 38772 56256
rect 38276 55946 38310 56222
rect 38738 56160 38772 56222
rect 38738 55946 38772 56002
rect 38276 55906 38772 55946
rect 38276 55630 38310 55906
rect 38738 55850 38772 55906
rect 38738 55630 38772 55692
rect 38276 55596 38772 55630
rect 43266 56222 43762 56256
rect 43266 55946 43300 56222
rect 43728 56160 43762 56222
rect 43728 55946 43762 56002
rect 43266 55906 43762 55946
rect 43266 55630 43300 55906
rect 43728 55850 43762 55906
rect 43728 55630 43762 55692
rect 43266 55596 43762 55630
rect 48256 56222 48752 56256
rect 48256 55946 48290 56222
rect 48718 56160 48752 56222
rect 48718 55946 48752 56002
rect 48256 55906 48752 55946
rect 48256 55630 48290 55906
rect 48718 55850 48752 55906
rect 48718 55630 48752 55692
rect 48256 55596 48752 55630
rect 53246 56222 53742 56256
rect 53246 55946 53280 56222
rect 53708 56160 53742 56222
rect 53708 55946 53742 56002
rect 53246 55906 53742 55946
rect 53246 55630 53280 55906
rect 53708 55850 53742 55906
rect 53708 55630 53742 55692
rect 53246 55596 53742 55630
rect 58236 56222 58732 56256
rect 58236 55946 58270 56222
rect 58698 56160 58732 56222
rect 58698 55946 58732 56002
rect 58236 55906 58732 55946
rect 58236 55630 58270 55906
rect 58698 55850 58732 55906
rect 58698 55630 58732 55692
rect 58236 55596 58732 55630
rect 63226 56222 63722 56256
rect 63226 55946 63260 56222
rect 63688 56160 63722 56222
rect 63688 55946 63722 56002
rect 63226 55906 63722 55946
rect 63226 55630 63260 55906
rect 63688 55850 63722 55906
rect 63688 55630 63722 55692
rect 63226 55596 63722 55630
rect 68216 56222 68712 56256
rect 68216 55946 68250 56222
rect 68678 56160 68712 56222
rect 68678 55946 68712 56002
rect 68216 55906 68712 55946
rect 68216 55630 68250 55906
rect 68678 55850 68712 55906
rect 68678 55630 68712 55692
rect 68216 55596 68712 55630
rect 73206 56222 73702 56256
rect 73206 55946 73240 56222
rect 73668 56160 73702 56222
rect 73668 55946 73702 56002
rect 73206 55906 73702 55946
rect 73206 55630 73240 55906
rect 73668 55850 73702 55906
rect 73668 55630 73702 55692
rect 73206 55596 73702 55630
rect 78196 56222 78692 56256
rect 78196 55946 78230 56222
rect 78658 56160 78692 56222
rect 78658 55946 78692 56002
rect 78196 55906 78692 55946
rect 78196 55630 78230 55906
rect 78658 55850 78692 55906
rect 78658 55630 78692 55692
rect 78196 55596 78692 55630
rect 3346 54512 3842 54546
rect 3346 54236 3380 54512
rect 3808 54450 3842 54512
rect 3808 54236 3842 54292
rect 3346 54196 3842 54236
rect 3346 53920 3380 54196
rect 3808 54140 3842 54196
rect 3808 53920 3842 53982
rect 3346 53886 3842 53920
rect 8336 54512 8832 54546
rect 8336 54236 8370 54512
rect 8798 54450 8832 54512
rect 8798 54236 8832 54292
rect 8336 54196 8832 54236
rect 8336 53920 8370 54196
rect 8798 54140 8832 54196
rect 8798 53920 8832 53982
rect 8336 53886 8832 53920
rect 13326 54512 13822 54546
rect 13326 54236 13360 54512
rect 13788 54450 13822 54512
rect 13788 54236 13822 54292
rect 13326 54196 13822 54236
rect 13326 53920 13360 54196
rect 13788 54140 13822 54196
rect 13788 53920 13822 53982
rect 13326 53886 13822 53920
rect 18316 54512 18812 54546
rect 18316 54236 18350 54512
rect 18778 54450 18812 54512
rect 18778 54236 18812 54292
rect 18316 54196 18812 54236
rect 18316 53920 18350 54196
rect 18778 54140 18812 54196
rect 18778 53920 18812 53982
rect 18316 53886 18812 53920
rect 23306 54512 23802 54546
rect 23306 54236 23340 54512
rect 23768 54450 23802 54512
rect 23768 54236 23802 54292
rect 23306 54196 23802 54236
rect 23306 53920 23340 54196
rect 23768 54140 23802 54196
rect 23768 53920 23802 53982
rect 23306 53886 23802 53920
rect 28296 54512 28792 54546
rect 28296 54236 28330 54512
rect 28758 54450 28792 54512
rect 28758 54236 28792 54292
rect 28296 54196 28792 54236
rect 28296 53920 28330 54196
rect 28758 54140 28792 54196
rect 28758 53920 28792 53982
rect 28296 53886 28792 53920
rect 33286 54512 33782 54546
rect 33286 54236 33320 54512
rect 33748 54450 33782 54512
rect 33748 54236 33782 54292
rect 33286 54196 33782 54236
rect 33286 53920 33320 54196
rect 33748 54140 33782 54196
rect 33748 53920 33782 53982
rect 33286 53886 33782 53920
rect 38276 54512 38772 54546
rect 38276 54236 38310 54512
rect 38738 54450 38772 54512
rect 38738 54236 38772 54292
rect 38276 54196 38772 54236
rect 38276 53920 38310 54196
rect 38738 54140 38772 54196
rect 38738 53920 38772 53982
rect 38276 53886 38772 53920
rect 43266 54512 43762 54546
rect 43266 54236 43300 54512
rect 43728 54450 43762 54512
rect 43728 54236 43762 54292
rect 43266 54196 43762 54236
rect 43266 53920 43300 54196
rect 43728 54140 43762 54196
rect 43728 53920 43762 53982
rect 43266 53886 43762 53920
rect 48256 54512 48752 54546
rect 48256 54236 48290 54512
rect 48718 54450 48752 54512
rect 48718 54236 48752 54292
rect 48256 54196 48752 54236
rect 48256 53920 48290 54196
rect 48718 54140 48752 54196
rect 48718 53920 48752 53982
rect 48256 53886 48752 53920
rect 53246 54512 53742 54546
rect 53246 54236 53280 54512
rect 53708 54450 53742 54512
rect 53708 54236 53742 54292
rect 53246 54196 53742 54236
rect 53246 53920 53280 54196
rect 53708 54140 53742 54196
rect 53708 53920 53742 53982
rect 53246 53886 53742 53920
rect 58236 54512 58732 54546
rect 58236 54236 58270 54512
rect 58698 54450 58732 54512
rect 58698 54236 58732 54292
rect 58236 54196 58732 54236
rect 58236 53920 58270 54196
rect 58698 54140 58732 54196
rect 58698 53920 58732 53982
rect 58236 53886 58732 53920
rect 63226 54512 63722 54546
rect 63226 54236 63260 54512
rect 63688 54450 63722 54512
rect 63688 54236 63722 54292
rect 63226 54196 63722 54236
rect 63226 53920 63260 54196
rect 63688 54140 63722 54196
rect 63688 53920 63722 53982
rect 63226 53886 63722 53920
rect 68216 54512 68712 54546
rect 68216 54236 68250 54512
rect 68678 54450 68712 54512
rect 68678 54236 68712 54292
rect 68216 54196 68712 54236
rect 68216 53920 68250 54196
rect 68678 54140 68712 54196
rect 68678 53920 68712 53982
rect 68216 53886 68712 53920
rect 73206 54512 73702 54546
rect 73206 54236 73240 54512
rect 73668 54450 73702 54512
rect 73668 54236 73702 54292
rect 73206 54196 73702 54236
rect 73206 53920 73240 54196
rect 73668 54140 73702 54196
rect 73668 53920 73702 53982
rect 73206 53886 73702 53920
rect 78196 54512 78692 54546
rect 78196 54236 78230 54512
rect 78658 54450 78692 54512
rect 78658 54236 78692 54292
rect 78196 54196 78692 54236
rect 78196 53920 78230 54196
rect 78658 54140 78692 54196
rect 78658 53920 78692 53982
rect 78196 53886 78692 53920
rect 3346 52802 3842 52836
rect 3346 52526 3380 52802
rect 3808 52740 3842 52802
rect 3808 52526 3842 52582
rect 3346 52486 3842 52526
rect 3346 52210 3380 52486
rect 3808 52430 3842 52486
rect 3808 52210 3842 52272
rect 3346 52176 3842 52210
rect 8336 52802 8832 52836
rect 8336 52526 8370 52802
rect 8798 52740 8832 52802
rect 8798 52526 8832 52582
rect 8336 52486 8832 52526
rect 8336 52210 8370 52486
rect 8798 52430 8832 52486
rect 8798 52210 8832 52272
rect 8336 52176 8832 52210
rect 13326 52802 13822 52836
rect 13326 52526 13360 52802
rect 13788 52740 13822 52802
rect 13788 52526 13822 52582
rect 13326 52486 13822 52526
rect 13326 52210 13360 52486
rect 13788 52430 13822 52486
rect 13788 52210 13822 52272
rect 13326 52176 13822 52210
rect 18316 52802 18812 52836
rect 18316 52526 18350 52802
rect 18778 52740 18812 52802
rect 18778 52526 18812 52582
rect 18316 52486 18812 52526
rect 18316 52210 18350 52486
rect 18778 52430 18812 52486
rect 18778 52210 18812 52272
rect 18316 52176 18812 52210
rect 23306 52802 23802 52836
rect 23306 52526 23340 52802
rect 23768 52740 23802 52802
rect 23768 52526 23802 52582
rect 23306 52486 23802 52526
rect 23306 52210 23340 52486
rect 23768 52430 23802 52486
rect 23768 52210 23802 52272
rect 23306 52176 23802 52210
rect 28296 52802 28792 52836
rect 28296 52526 28330 52802
rect 28758 52740 28792 52802
rect 28758 52526 28792 52582
rect 28296 52486 28792 52526
rect 28296 52210 28330 52486
rect 28758 52430 28792 52486
rect 28758 52210 28792 52272
rect 28296 52176 28792 52210
rect 33286 52802 33782 52836
rect 33286 52526 33320 52802
rect 33748 52740 33782 52802
rect 33748 52526 33782 52582
rect 33286 52486 33782 52526
rect 33286 52210 33320 52486
rect 33748 52430 33782 52486
rect 33748 52210 33782 52272
rect 33286 52176 33782 52210
rect 38276 52802 38772 52836
rect 38276 52526 38310 52802
rect 38738 52740 38772 52802
rect 38738 52526 38772 52582
rect 38276 52486 38772 52526
rect 38276 52210 38310 52486
rect 38738 52430 38772 52486
rect 38738 52210 38772 52272
rect 38276 52176 38772 52210
rect 43266 52802 43762 52836
rect 43266 52526 43300 52802
rect 43728 52740 43762 52802
rect 43728 52526 43762 52582
rect 43266 52486 43762 52526
rect 43266 52210 43300 52486
rect 43728 52430 43762 52486
rect 43728 52210 43762 52272
rect 43266 52176 43762 52210
rect 48256 52802 48752 52836
rect 48256 52526 48290 52802
rect 48718 52740 48752 52802
rect 48718 52526 48752 52582
rect 48256 52486 48752 52526
rect 48256 52210 48290 52486
rect 48718 52430 48752 52486
rect 48718 52210 48752 52272
rect 48256 52176 48752 52210
rect 53246 52802 53742 52836
rect 53246 52526 53280 52802
rect 53708 52740 53742 52802
rect 53708 52526 53742 52582
rect 53246 52486 53742 52526
rect 53246 52210 53280 52486
rect 53708 52430 53742 52486
rect 53708 52210 53742 52272
rect 53246 52176 53742 52210
rect 58236 52802 58732 52836
rect 58236 52526 58270 52802
rect 58698 52740 58732 52802
rect 58698 52526 58732 52582
rect 58236 52486 58732 52526
rect 58236 52210 58270 52486
rect 58698 52430 58732 52486
rect 58698 52210 58732 52272
rect 58236 52176 58732 52210
rect 63226 52802 63722 52836
rect 63226 52526 63260 52802
rect 63688 52740 63722 52802
rect 63688 52526 63722 52582
rect 63226 52486 63722 52526
rect 63226 52210 63260 52486
rect 63688 52430 63722 52486
rect 63688 52210 63722 52272
rect 63226 52176 63722 52210
rect 68216 52802 68712 52836
rect 68216 52526 68250 52802
rect 68678 52740 68712 52802
rect 68678 52526 68712 52582
rect 68216 52486 68712 52526
rect 68216 52210 68250 52486
rect 68678 52430 68712 52486
rect 68678 52210 68712 52272
rect 68216 52176 68712 52210
rect 73206 52802 73702 52836
rect 73206 52526 73240 52802
rect 73668 52740 73702 52802
rect 73668 52526 73702 52582
rect 73206 52486 73702 52526
rect 73206 52210 73240 52486
rect 73668 52430 73702 52486
rect 73668 52210 73702 52272
rect 73206 52176 73702 52210
rect 78196 52802 78692 52836
rect 78196 52526 78230 52802
rect 78658 52740 78692 52802
rect 78658 52526 78692 52582
rect 78196 52486 78692 52526
rect 78196 52210 78230 52486
rect 78658 52430 78692 52486
rect 78658 52210 78692 52272
rect 78196 52176 78692 52210
rect 3346 51092 3842 51126
rect 3346 50816 3380 51092
rect 3808 51030 3842 51092
rect 3808 50816 3842 50872
rect 3346 50776 3842 50816
rect 3346 50500 3380 50776
rect 3808 50720 3842 50776
rect 3808 50500 3842 50562
rect 3346 50466 3842 50500
rect 8336 51092 8832 51126
rect 8336 50816 8370 51092
rect 8798 51030 8832 51092
rect 8798 50816 8832 50872
rect 8336 50776 8832 50816
rect 8336 50500 8370 50776
rect 8798 50720 8832 50776
rect 8798 50500 8832 50562
rect 8336 50466 8832 50500
rect 13326 51092 13822 51126
rect 13326 50816 13360 51092
rect 13788 51030 13822 51092
rect 13788 50816 13822 50872
rect 13326 50776 13822 50816
rect 13326 50500 13360 50776
rect 13788 50720 13822 50776
rect 13788 50500 13822 50562
rect 13326 50466 13822 50500
rect 18316 51092 18812 51126
rect 18316 50816 18350 51092
rect 18778 51030 18812 51092
rect 18778 50816 18812 50872
rect 18316 50776 18812 50816
rect 18316 50500 18350 50776
rect 18778 50720 18812 50776
rect 18778 50500 18812 50562
rect 18316 50466 18812 50500
rect 23306 51092 23802 51126
rect 23306 50816 23340 51092
rect 23768 51030 23802 51092
rect 23768 50816 23802 50872
rect 23306 50776 23802 50816
rect 23306 50500 23340 50776
rect 23768 50720 23802 50776
rect 23768 50500 23802 50562
rect 23306 50466 23802 50500
rect 28296 51092 28792 51126
rect 28296 50816 28330 51092
rect 28758 51030 28792 51092
rect 28758 50816 28792 50872
rect 28296 50776 28792 50816
rect 28296 50500 28330 50776
rect 28758 50720 28792 50776
rect 28758 50500 28792 50562
rect 28296 50466 28792 50500
rect 33286 51092 33782 51126
rect 33286 50816 33320 51092
rect 33748 51030 33782 51092
rect 33748 50816 33782 50872
rect 33286 50776 33782 50816
rect 33286 50500 33320 50776
rect 33748 50720 33782 50776
rect 33748 50500 33782 50562
rect 33286 50466 33782 50500
rect 38276 51092 38772 51126
rect 38276 50816 38310 51092
rect 38738 51030 38772 51092
rect 38738 50816 38772 50872
rect 38276 50776 38772 50816
rect 38276 50500 38310 50776
rect 38738 50720 38772 50776
rect 38738 50500 38772 50562
rect 38276 50466 38772 50500
rect 43266 51092 43762 51126
rect 43266 50816 43300 51092
rect 43728 51030 43762 51092
rect 43728 50816 43762 50872
rect 43266 50776 43762 50816
rect 43266 50500 43300 50776
rect 43728 50720 43762 50776
rect 43728 50500 43762 50562
rect 43266 50466 43762 50500
rect 48256 51092 48752 51126
rect 48256 50816 48290 51092
rect 48718 51030 48752 51092
rect 48718 50816 48752 50872
rect 48256 50776 48752 50816
rect 48256 50500 48290 50776
rect 48718 50720 48752 50776
rect 48718 50500 48752 50562
rect 48256 50466 48752 50500
rect 53246 51092 53742 51126
rect 53246 50816 53280 51092
rect 53708 51030 53742 51092
rect 53708 50816 53742 50872
rect 53246 50776 53742 50816
rect 53246 50500 53280 50776
rect 53708 50720 53742 50776
rect 53708 50500 53742 50562
rect 53246 50466 53742 50500
rect 58236 51092 58732 51126
rect 58236 50816 58270 51092
rect 58698 51030 58732 51092
rect 58698 50816 58732 50872
rect 58236 50776 58732 50816
rect 58236 50500 58270 50776
rect 58698 50720 58732 50776
rect 58698 50500 58732 50562
rect 58236 50466 58732 50500
rect 63226 51092 63722 51126
rect 63226 50816 63260 51092
rect 63688 51030 63722 51092
rect 63688 50816 63722 50872
rect 63226 50776 63722 50816
rect 63226 50500 63260 50776
rect 63688 50720 63722 50776
rect 63688 50500 63722 50562
rect 63226 50466 63722 50500
rect 68216 51092 68712 51126
rect 68216 50816 68250 51092
rect 68678 51030 68712 51092
rect 68678 50816 68712 50872
rect 68216 50776 68712 50816
rect 68216 50500 68250 50776
rect 68678 50720 68712 50776
rect 68678 50500 68712 50562
rect 68216 50466 68712 50500
rect 73206 51092 73702 51126
rect 73206 50816 73240 51092
rect 73668 51030 73702 51092
rect 73668 50816 73702 50872
rect 73206 50776 73702 50816
rect 73206 50500 73240 50776
rect 73668 50720 73702 50776
rect 73668 50500 73702 50562
rect 73206 50466 73702 50500
rect 78196 51092 78692 51126
rect 78196 50816 78230 51092
rect 78658 51030 78692 51092
rect 78658 50816 78692 50872
rect 78196 50776 78692 50816
rect 78196 50500 78230 50776
rect 78658 50720 78692 50776
rect 78658 50500 78692 50562
rect 78196 50466 78692 50500
rect 3346 49382 3842 49416
rect 3346 49106 3380 49382
rect 3808 49320 3842 49382
rect 3808 49106 3842 49162
rect 3346 49066 3842 49106
rect 3346 48790 3380 49066
rect 3808 49010 3842 49066
rect 3808 48790 3842 48852
rect 3346 48756 3842 48790
rect 8336 49382 8832 49416
rect 8336 49106 8370 49382
rect 8798 49320 8832 49382
rect 8798 49106 8832 49162
rect 8336 49066 8832 49106
rect 8336 48790 8370 49066
rect 8798 49010 8832 49066
rect 8798 48790 8832 48852
rect 8336 48756 8832 48790
rect 13326 49382 13822 49416
rect 13326 49106 13360 49382
rect 13788 49320 13822 49382
rect 13788 49106 13822 49162
rect 13326 49066 13822 49106
rect 13326 48790 13360 49066
rect 13788 49010 13822 49066
rect 13788 48790 13822 48852
rect 13326 48756 13822 48790
rect 18316 49382 18812 49416
rect 18316 49106 18350 49382
rect 18778 49320 18812 49382
rect 18778 49106 18812 49162
rect 18316 49066 18812 49106
rect 18316 48790 18350 49066
rect 18778 49010 18812 49066
rect 18778 48790 18812 48852
rect 18316 48756 18812 48790
rect 23306 49382 23802 49416
rect 23306 49106 23340 49382
rect 23768 49320 23802 49382
rect 23768 49106 23802 49162
rect 23306 49066 23802 49106
rect 23306 48790 23340 49066
rect 23768 49010 23802 49066
rect 23768 48790 23802 48852
rect 23306 48756 23802 48790
rect 28296 49382 28792 49416
rect 28296 49106 28330 49382
rect 28758 49320 28792 49382
rect 28758 49106 28792 49162
rect 28296 49066 28792 49106
rect 28296 48790 28330 49066
rect 28758 49010 28792 49066
rect 28758 48790 28792 48852
rect 28296 48756 28792 48790
rect 33286 49382 33782 49416
rect 33286 49106 33320 49382
rect 33748 49320 33782 49382
rect 33748 49106 33782 49162
rect 33286 49066 33782 49106
rect 33286 48790 33320 49066
rect 33748 49010 33782 49066
rect 33748 48790 33782 48852
rect 33286 48756 33782 48790
rect 38276 49382 38772 49416
rect 38276 49106 38310 49382
rect 38738 49320 38772 49382
rect 38738 49106 38772 49162
rect 38276 49066 38772 49106
rect 38276 48790 38310 49066
rect 38738 49010 38772 49066
rect 38738 48790 38772 48852
rect 38276 48756 38772 48790
rect 43266 49382 43762 49416
rect 43266 49106 43300 49382
rect 43728 49320 43762 49382
rect 43728 49106 43762 49162
rect 43266 49066 43762 49106
rect 43266 48790 43300 49066
rect 43728 49010 43762 49066
rect 43728 48790 43762 48852
rect 43266 48756 43762 48790
rect 48256 49382 48752 49416
rect 48256 49106 48290 49382
rect 48718 49320 48752 49382
rect 48718 49106 48752 49162
rect 48256 49066 48752 49106
rect 48256 48790 48290 49066
rect 48718 49010 48752 49066
rect 48718 48790 48752 48852
rect 48256 48756 48752 48790
rect 53246 49382 53742 49416
rect 53246 49106 53280 49382
rect 53708 49320 53742 49382
rect 53708 49106 53742 49162
rect 53246 49066 53742 49106
rect 53246 48790 53280 49066
rect 53708 49010 53742 49066
rect 53708 48790 53742 48852
rect 53246 48756 53742 48790
rect 58236 49382 58732 49416
rect 58236 49106 58270 49382
rect 58698 49320 58732 49382
rect 58698 49106 58732 49162
rect 58236 49066 58732 49106
rect 58236 48790 58270 49066
rect 58698 49010 58732 49066
rect 58698 48790 58732 48852
rect 58236 48756 58732 48790
rect 63226 49382 63722 49416
rect 63226 49106 63260 49382
rect 63688 49320 63722 49382
rect 63688 49106 63722 49162
rect 63226 49066 63722 49106
rect 63226 48790 63260 49066
rect 63688 49010 63722 49066
rect 63688 48790 63722 48852
rect 63226 48756 63722 48790
rect 68216 49382 68712 49416
rect 68216 49106 68250 49382
rect 68678 49320 68712 49382
rect 68678 49106 68712 49162
rect 68216 49066 68712 49106
rect 68216 48790 68250 49066
rect 68678 49010 68712 49066
rect 68678 48790 68712 48852
rect 68216 48756 68712 48790
rect 73206 49382 73702 49416
rect 73206 49106 73240 49382
rect 73668 49320 73702 49382
rect 73668 49106 73702 49162
rect 73206 49066 73702 49106
rect 73206 48790 73240 49066
rect 73668 49010 73702 49066
rect 73668 48790 73702 48852
rect 73206 48756 73702 48790
rect 78196 49382 78692 49416
rect 78196 49106 78230 49382
rect 78658 49320 78692 49382
rect 78658 49106 78692 49162
rect 78196 49066 78692 49106
rect 78196 48790 78230 49066
rect 78658 49010 78692 49066
rect 78658 48790 78692 48852
rect 78196 48756 78692 48790
rect 3346 47672 3842 47706
rect 3346 47396 3380 47672
rect 3808 47610 3842 47672
rect 3808 47396 3842 47452
rect 3346 47356 3842 47396
rect 3346 47080 3380 47356
rect 3808 47300 3842 47356
rect 3808 47080 3842 47142
rect 3346 47046 3842 47080
rect 8336 47672 8832 47706
rect 8336 47396 8370 47672
rect 8798 47610 8832 47672
rect 8798 47396 8832 47452
rect 8336 47356 8832 47396
rect 8336 47080 8370 47356
rect 8798 47300 8832 47356
rect 8798 47080 8832 47142
rect 8336 47046 8832 47080
rect 13326 47672 13822 47706
rect 13326 47396 13360 47672
rect 13788 47610 13822 47672
rect 13788 47396 13822 47452
rect 13326 47356 13822 47396
rect 13326 47080 13360 47356
rect 13788 47300 13822 47356
rect 13788 47080 13822 47142
rect 13326 47046 13822 47080
rect 18316 47672 18812 47706
rect 18316 47396 18350 47672
rect 18778 47610 18812 47672
rect 18778 47396 18812 47452
rect 18316 47356 18812 47396
rect 18316 47080 18350 47356
rect 18778 47300 18812 47356
rect 18778 47080 18812 47142
rect 18316 47046 18812 47080
rect 23306 47672 23802 47706
rect 23306 47396 23340 47672
rect 23768 47610 23802 47672
rect 23768 47396 23802 47452
rect 23306 47356 23802 47396
rect 23306 47080 23340 47356
rect 23768 47300 23802 47356
rect 23768 47080 23802 47142
rect 23306 47046 23802 47080
rect 28296 47672 28792 47706
rect 28296 47396 28330 47672
rect 28758 47610 28792 47672
rect 28758 47396 28792 47452
rect 28296 47356 28792 47396
rect 28296 47080 28330 47356
rect 28758 47300 28792 47356
rect 28758 47080 28792 47142
rect 28296 47046 28792 47080
rect 33286 47672 33782 47706
rect 33286 47396 33320 47672
rect 33748 47610 33782 47672
rect 33748 47396 33782 47452
rect 33286 47356 33782 47396
rect 33286 47080 33320 47356
rect 33748 47300 33782 47356
rect 33748 47080 33782 47142
rect 33286 47046 33782 47080
rect 38276 47672 38772 47706
rect 38276 47396 38310 47672
rect 38738 47610 38772 47672
rect 38738 47396 38772 47452
rect 38276 47356 38772 47396
rect 38276 47080 38310 47356
rect 38738 47300 38772 47356
rect 38738 47080 38772 47142
rect 38276 47046 38772 47080
rect 43266 47672 43762 47706
rect 43266 47396 43300 47672
rect 43728 47610 43762 47672
rect 43728 47396 43762 47452
rect 43266 47356 43762 47396
rect 43266 47080 43300 47356
rect 43728 47300 43762 47356
rect 43728 47080 43762 47142
rect 43266 47046 43762 47080
rect 48256 47672 48752 47706
rect 48256 47396 48290 47672
rect 48718 47610 48752 47672
rect 48718 47396 48752 47452
rect 48256 47356 48752 47396
rect 48256 47080 48290 47356
rect 48718 47300 48752 47356
rect 48718 47080 48752 47142
rect 48256 47046 48752 47080
rect 53246 47672 53742 47706
rect 53246 47396 53280 47672
rect 53708 47610 53742 47672
rect 53708 47396 53742 47452
rect 53246 47356 53742 47396
rect 53246 47080 53280 47356
rect 53708 47300 53742 47356
rect 53708 47080 53742 47142
rect 53246 47046 53742 47080
rect 58236 47672 58732 47706
rect 58236 47396 58270 47672
rect 58698 47610 58732 47672
rect 58698 47396 58732 47452
rect 58236 47356 58732 47396
rect 58236 47080 58270 47356
rect 58698 47300 58732 47356
rect 58698 47080 58732 47142
rect 58236 47046 58732 47080
rect 63226 47672 63722 47706
rect 63226 47396 63260 47672
rect 63688 47610 63722 47672
rect 63688 47396 63722 47452
rect 63226 47356 63722 47396
rect 63226 47080 63260 47356
rect 63688 47300 63722 47356
rect 63688 47080 63722 47142
rect 63226 47046 63722 47080
rect 68216 47672 68712 47706
rect 68216 47396 68250 47672
rect 68678 47610 68712 47672
rect 68678 47396 68712 47452
rect 68216 47356 68712 47396
rect 68216 47080 68250 47356
rect 68678 47300 68712 47356
rect 68678 47080 68712 47142
rect 68216 47046 68712 47080
rect 73206 47672 73702 47706
rect 73206 47396 73240 47672
rect 73668 47610 73702 47672
rect 73668 47396 73702 47452
rect 73206 47356 73702 47396
rect 73206 47080 73240 47356
rect 73668 47300 73702 47356
rect 73668 47080 73702 47142
rect 73206 47046 73702 47080
rect 78196 47672 78692 47706
rect 78196 47396 78230 47672
rect 78658 47610 78692 47672
rect 78658 47396 78692 47452
rect 78196 47356 78692 47396
rect 78196 47080 78230 47356
rect 78658 47300 78692 47356
rect 78658 47080 78692 47142
rect 78196 47046 78692 47080
rect 3346 45962 3842 45996
rect 3346 45686 3380 45962
rect 3808 45900 3842 45962
rect 3808 45686 3842 45742
rect 3346 45646 3842 45686
rect 3346 45370 3380 45646
rect 3808 45590 3842 45646
rect 3808 45370 3842 45432
rect 3346 45336 3842 45370
rect 8336 45962 8832 45996
rect 8336 45686 8370 45962
rect 8798 45900 8832 45962
rect 8798 45686 8832 45742
rect 8336 45646 8832 45686
rect 8336 45370 8370 45646
rect 8798 45590 8832 45646
rect 8798 45370 8832 45432
rect 8336 45336 8832 45370
rect 13326 45962 13822 45996
rect 13326 45686 13360 45962
rect 13788 45900 13822 45962
rect 13788 45686 13822 45742
rect 13326 45646 13822 45686
rect 13326 45370 13360 45646
rect 13788 45590 13822 45646
rect 13788 45370 13822 45432
rect 13326 45336 13822 45370
rect 18316 45962 18812 45996
rect 18316 45686 18350 45962
rect 18778 45900 18812 45962
rect 18778 45686 18812 45742
rect 18316 45646 18812 45686
rect 18316 45370 18350 45646
rect 18778 45590 18812 45646
rect 18778 45370 18812 45432
rect 18316 45336 18812 45370
rect 23306 45962 23802 45996
rect 23306 45686 23340 45962
rect 23768 45900 23802 45962
rect 23768 45686 23802 45742
rect 23306 45646 23802 45686
rect 23306 45370 23340 45646
rect 23768 45590 23802 45646
rect 23768 45370 23802 45432
rect 23306 45336 23802 45370
rect 28296 45962 28792 45996
rect 28296 45686 28330 45962
rect 28758 45900 28792 45962
rect 28758 45686 28792 45742
rect 28296 45646 28792 45686
rect 28296 45370 28330 45646
rect 28758 45590 28792 45646
rect 28758 45370 28792 45432
rect 28296 45336 28792 45370
rect 33286 45962 33782 45996
rect 33286 45686 33320 45962
rect 33748 45900 33782 45962
rect 33748 45686 33782 45742
rect 33286 45646 33782 45686
rect 33286 45370 33320 45646
rect 33748 45590 33782 45646
rect 33748 45370 33782 45432
rect 33286 45336 33782 45370
rect 38276 45962 38772 45996
rect 38276 45686 38310 45962
rect 38738 45900 38772 45962
rect 38738 45686 38772 45742
rect 38276 45646 38772 45686
rect 38276 45370 38310 45646
rect 38738 45590 38772 45646
rect 38738 45370 38772 45432
rect 38276 45336 38772 45370
rect 43266 45962 43762 45996
rect 43266 45686 43300 45962
rect 43728 45900 43762 45962
rect 43728 45686 43762 45742
rect 43266 45646 43762 45686
rect 43266 45370 43300 45646
rect 43728 45590 43762 45646
rect 43728 45370 43762 45432
rect 43266 45336 43762 45370
rect 48256 45962 48752 45996
rect 48256 45686 48290 45962
rect 48718 45900 48752 45962
rect 48718 45686 48752 45742
rect 48256 45646 48752 45686
rect 48256 45370 48290 45646
rect 48718 45590 48752 45646
rect 48718 45370 48752 45432
rect 48256 45336 48752 45370
rect 53246 45962 53742 45996
rect 53246 45686 53280 45962
rect 53708 45900 53742 45962
rect 53708 45686 53742 45742
rect 53246 45646 53742 45686
rect 53246 45370 53280 45646
rect 53708 45590 53742 45646
rect 53708 45370 53742 45432
rect 53246 45336 53742 45370
rect 58236 45962 58732 45996
rect 58236 45686 58270 45962
rect 58698 45900 58732 45962
rect 58698 45686 58732 45742
rect 58236 45646 58732 45686
rect 58236 45370 58270 45646
rect 58698 45590 58732 45646
rect 58698 45370 58732 45432
rect 58236 45336 58732 45370
rect 63226 45962 63722 45996
rect 63226 45686 63260 45962
rect 63688 45900 63722 45962
rect 63688 45686 63722 45742
rect 63226 45646 63722 45686
rect 63226 45370 63260 45646
rect 63688 45590 63722 45646
rect 63688 45370 63722 45432
rect 63226 45336 63722 45370
rect 68216 45962 68712 45996
rect 68216 45686 68250 45962
rect 68678 45900 68712 45962
rect 68678 45686 68712 45742
rect 68216 45646 68712 45686
rect 68216 45370 68250 45646
rect 68678 45590 68712 45646
rect 68678 45370 68712 45432
rect 68216 45336 68712 45370
rect 73206 45962 73702 45996
rect 73206 45686 73240 45962
rect 73668 45900 73702 45962
rect 73668 45686 73702 45742
rect 73206 45646 73702 45686
rect 73206 45370 73240 45646
rect 73668 45590 73702 45646
rect 73668 45370 73702 45432
rect 73206 45336 73702 45370
rect 78196 45962 78692 45996
rect 78196 45686 78230 45962
rect 78658 45900 78692 45962
rect 78658 45686 78692 45742
rect 78196 45646 78692 45686
rect 78196 45370 78230 45646
rect 78658 45590 78692 45646
rect 78658 45370 78692 45432
rect 78196 45336 78692 45370
rect 3346 44252 3842 44286
rect 3346 43976 3380 44252
rect 3808 44190 3842 44252
rect 3808 43976 3842 44032
rect 3346 43936 3842 43976
rect 3346 43660 3380 43936
rect 3808 43880 3842 43936
rect 3808 43660 3842 43722
rect 3346 43626 3842 43660
rect 8336 44252 8832 44286
rect 8336 43976 8370 44252
rect 8798 44190 8832 44252
rect 8798 43976 8832 44032
rect 8336 43936 8832 43976
rect 8336 43660 8370 43936
rect 8798 43880 8832 43936
rect 8798 43660 8832 43722
rect 8336 43626 8832 43660
rect 13326 44252 13822 44286
rect 13326 43976 13360 44252
rect 13788 44190 13822 44252
rect 13788 43976 13822 44032
rect 13326 43936 13822 43976
rect 13326 43660 13360 43936
rect 13788 43880 13822 43936
rect 13788 43660 13822 43722
rect 13326 43626 13822 43660
rect 18316 44252 18812 44286
rect 18316 43976 18350 44252
rect 18778 44190 18812 44252
rect 18778 43976 18812 44032
rect 18316 43936 18812 43976
rect 18316 43660 18350 43936
rect 18778 43880 18812 43936
rect 18778 43660 18812 43722
rect 18316 43626 18812 43660
rect 23306 44252 23802 44286
rect 23306 43976 23340 44252
rect 23768 44190 23802 44252
rect 23768 43976 23802 44032
rect 23306 43936 23802 43976
rect 23306 43660 23340 43936
rect 23768 43880 23802 43936
rect 23768 43660 23802 43722
rect 23306 43626 23802 43660
rect 28296 44252 28792 44286
rect 28296 43976 28330 44252
rect 28758 44190 28792 44252
rect 28758 43976 28792 44032
rect 28296 43936 28792 43976
rect 28296 43660 28330 43936
rect 28758 43880 28792 43936
rect 28758 43660 28792 43722
rect 28296 43626 28792 43660
rect 33286 44252 33782 44286
rect 33286 43976 33320 44252
rect 33748 44190 33782 44252
rect 33748 43976 33782 44032
rect 33286 43936 33782 43976
rect 33286 43660 33320 43936
rect 33748 43880 33782 43936
rect 33748 43660 33782 43722
rect 33286 43626 33782 43660
rect 38276 44252 38772 44286
rect 38276 43976 38310 44252
rect 38738 44190 38772 44252
rect 38738 43976 38772 44032
rect 38276 43936 38772 43976
rect 38276 43660 38310 43936
rect 38738 43880 38772 43936
rect 38738 43660 38772 43722
rect 38276 43626 38772 43660
rect 43266 44252 43762 44286
rect 43266 43976 43300 44252
rect 43728 44190 43762 44252
rect 43728 43976 43762 44032
rect 43266 43936 43762 43976
rect 43266 43660 43300 43936
rect 43728 43880 43762 43936
rect 43728 43660 43762 43722
rect 43266 43626 43762 43660
rect 48256 44252 48752 44286
rect 48256 43976 48290 44252
rect 48718 44190 48752 44252
rect 48718 43976 48752 44032
rect 48256 43936 48752 43976
rect 48256 43660 48290 43936
rect 48718 43880 48752 43936
rect 48718 43660 48752 43722
rect 48256 43626 48752 43660
rect 53246 44252 53742 44286
rect 53246 43976 53280 44252
rect 53708 44190 53742 44252
rect 53708 43976 53742 44032
rect 53246 43936 53742 43976
rect 53246 43660 53280 43936
rect 53708 43880 53742 43936
rect 53708 43660 53742 43722
rect 53246 43626 53742 43660
rect 58236 44252 58732 44286
rect 58236 43976 58270 44252
rect 58698 44190 58732 44252
rect 58698 43976 58732 44032
rect 58236 43936 58732 43976
rect 58236 43660 58270 43936
rect 58698 43880 58732 43936
rect 58698 43660 58732 43722
rect 58236 43626 58732 43660
rect 63226 44252 63722 44286
rect 63226 43976 63260 44252
rect 63688 44190 63722 44252
rect 63688 43976 63722 44032
rect 63226 43936 63722 43976
rect 63226 43660 63260 43936
rect 63688 43880 63722 43936
rect 63688 43660 63722 43722
rect 63226 43626 63722 43660
rect 68216 44252 68712 44286
rect 68216 43976 68250 44252
rect 68678 44190 68712 44252
rect 68678 43976 68712 44032
rect 68216 43936 68712 43976
rect 68216 43660 68250 43936
rect 68678 43880 68712 43936
rect 68678 43660 68712 43722
rect 68216 43626 68712 43660
rect 73206 44252 73702 44286
rect 73206 43976 73240 44252
rect 73668 44190 73702 44252
rect 73668 43976 73702 44032
rect 73206 43936 73702 43976
rect 73206 43660 73240 43936
rect 73668 43880 73702 43936
rect 73668 43660 73702 43722
rect 73206 43626 73702 43660
rect 78196 44252 78692 44286
rect 78196 43976 78230 44252
rect 78658 44190 78692 44252
rect 78658 43976 78692 44032
rect 78196 43936 78692 43976
rect 78196 43660 78230 43936
rect 78658 43880 78692 43936
rect 78658 43660 78692 43722
rect 78196 43626 78692 43660
rect 3346 42542 3842 42576
rect 3346 42266 3380 42542
rect 3808 42480 3842 42542
rect 3808 42266 3842 42322
rect 3346 42226 3842 42266
rect 3346 41950 3380 42226
rect 3808 42170 3842 42226
rect 3808 41950 3842 42012
rect 3346 41916 3842 41950
rect 8336 42542 8832 42576
rect 8336 42266 8370 42542
rect 8798 42480 8832 42542
rect 8798 42266 8832 42322
rect 8336 42226 8832 42266
rect 8336 41950 8370 42226
rect 8798 42170 8832 42226
rect 8798 41950 8832 42012
rect 8336 41916 8832 41950
rect 13326 42542 13822 42576
rect 13326 42266 13360 42542
rect 13788 42480 13822 42542
rect 13788 42266 13822 42322
rect 13326 42226 13822 42266
rect 13326 41950 13360 42226
rect 13788 42170 13822 42226
rect 13788 41950 13822 42012
rect 13326 41916 13822 41950
rect 18316 42542 18812 42576
rect 18316 42266 18350 42542
rect 18778 42480 18812 42542
rect 18778 42266 18812 42322
rect 18316 42226 18812 42266
rect 18316 41950 18350 42226
rect 18778 42170 18812 42226
rect 18778 41950 18812 42012
rect 18316 41916 18812 41950
rect 23306 42542 23802 42576
rect 23306 42266 23340 42542
rect 23768 42480 23802 42542
rect 23768 42266 23802 42322
rect 23306 42226 23802 42266
rect 23306 41950 23340 42226
rect 23768 42170 23802 42226
rect 23768 41950 23802 42012
rect 23306 41916 23802 41950
rect 28296 42542 28792 42576
rect 28296 42266 28330 42542
rect 28758 42480 28792 42542
rect 28758 42266 28792 42322
rect 28296 42226 28792 42266
rect 28296 41950 28330 42226
rect 28758 42170 28792 42226
rect 28758 41950 28792 42012
rect 28296 41916 28792 41950
rect 33286 42542 33782 42576
rect 33286 42266 33320 42542
rect 33748 42480 33782 42542
rect 33748 42266 33782 42322
rect 33286 42226 33782 42266
rect 33286 41950 33320 42226
rect 33748 42170 33782 42226
rect 33748 41950 33782 42012
rect 33286 41916 33782 41950
rect 38276 42542 38772 42576
rect 38276 42266 38310 42542
rect 38738 42480 38772 42542
rect 38738 42266 38772 42322
rect 38276 42226 38772 42266
rect 38276 41950 38310 42226
rect 38738 42170 38772 42226
rect 38738 41950 38772 42012
rect 38276 41916 38772 41950
rect 43266 42542 43762 42576
rect 43266 42266 43300 42542
rect 43728 42480 43762 42542
rect 43728 42266 43762 42322
rect 43266 42226 43762 42266
rect 43266 41950 43300 42226
rect 43728 42170 43762 42226
rect 43728 41950 43762 42012
rect 43266 41916 43762 41950
rect 48256 42542 48752 42576
rect 48256 42266 48290 42542
rect 48718 42480 48752 42542
rect 48718 42266 48752 42322
rect 48256 42226 48752 42266
rect 48256 41950 48290 42226
rect 48718 42170 48752 42226
rect 48718 41950 48752 42012
rect 48256 41916 48752 41950
rect 53246 42542 53742 42576
rect 53246 42266 53280 42542
rect 53708 42480 53742 42542
rect 53708 42266 53742 42322
rect 53246 42226 53742 42266
rect 53246 41950 53280 42226
rect 53708 42170 53742 42226
rect 53708 41950 53742 42012
rect 53246 41916 53742 41950
rect 58236 42542 58732 42576
rect 58236 42266 58270 42542
rect 58698 42480 58732 42542
rect 58698 42266 58732 42322
rect 58236 42226 58732 42266
rect 58236 41950 58270 42226
rect 58698 42170 58732 42226
rect 58698 41950 58732 42012
rect 58236 41916 58732 41950
rect 63226 42542 63722 42576
rect 63226 42266 63260 42542
rect 63688 42480 63722 42542
rect 63688 42266 63722 42322
rect 63226 42226 63722 42266
rect 63226 41950 63260 42226
rect 63688 42170 63722 42226
rect 63688 41950 63722 42012
rect 63226 41916 63722 41950
rect 68216 42542 68712 42576
rect 68216 42266 68250 42542
rect 68678 42480 68712 42542
rect 68678 42266 68712 42322
rect 68216 42226 68712 42266
rect 68216 41950 68250 42226
rect 68678 42170 68712 42226
rect 68678 41950 68712 42012
rect 68216 41916 68712 41950
rect 73206 42542 73702 42576
rect 73206 42266 73240 42542
rect 73668 42480 73702 42542
rect 73668 42266 73702 42322
rect 73206 42226 73702 42266
rect 73206 41950 73240 42226
rect 73668 42170 73702 42226
rect 73668 41950 73702 42012
rect 73206 41916 73702 41950
rect 78196 42542 78692 42576
rect 78196 42266 78230 42542
rect 78658 42480 78692 42542
rect 78658 42266 78692 42322
rect 78196 42226 78692 42266
rect 78196 41950 78230 42226
rect 78658 42170 78692 42226
rect 78658 41950 78692 42012
rect 78196 41916 78692 41950
rect 3346 40832 3842 40866
rect 3346 40556 3380 40832
rect 3808 40770 3842 40832
rect 3808 40556 3842 40612
rect 3346 40516 3842 40556
rect 3346 40240 3380 40516
rect 3808 40460 3842 40516
rect 3808 40240 3842 40302
rect 3346 40206 3842 40240
rect 8336 40832 8832 40866
rect 8336 40556 8370 40832
rect 8798 40770 8832 40832
rect 8798 40556 8832 40612
rect 8336 40516 8832 40556
rect 8336 40240 8370 40516
rect 8798 40460 8832 40516
rect 8798 40240 8832 40302
rect 8336 40206 8832 40240
rect 13326 40832 13822 40866
rect 13326 40556 13360 40832
rect 13788 40770 13822 40832
rect 13788 40556 13822 40612
rect 13326 40516 13822 40556
rect 13326 40240 13360 40516
rect 13788 40460 13822 40516
rect 13788 40240 13822 40302
rect 13326 40206 13822 40240
rect 18316 40832 18812 40866
rect 18316 40556 18350 40832
rect 18778 40770 18812 40832
rect 18778 40556 18812 40612
rect 18316 40516 18812 40556
rect 18316 40240 18350 40516
rect 18778 40460 18812 40516
rect 18778 40240 18812 40302
rect 18316 40206 18812 40240
rect 23306 40832 23802 40866
rect 23306 40556 23340 40832
rect 23768 40770 23802 40832
rect 23768 40556 23802 40612
rect 23306 40516 23802 40556
rect 23306 40240 23340 40516
rect 23768 40460 23802 40516
rect 23768 40240 23802 40302
rect 23306 40206 23802 40240
rect 28296 40832 28792 40866
rect 28296 40556 28330 40832
rect 28758 40770 28792 40832
rect 28758 40556 28792 40612
rect 28296 40516 28792 40556
rect 28296 40240 28330 40516
rect 28758 40460 28792 40516
rect 28758 40240 28792 40302
rect 28296 40206 28792 40240
rect 33286 40832 33782 40866
rect 33286 40556 33320 40832
rect 33748 40770 33782 40832
rect 33748 40556 33782 40612
rect 33286 40516 33782 40556
rect 33286 40240 33320 40516
rect 33748 40460 33782 40516
rect 33748 40240 33782 40302
rect 33286 40206 33782 40240
rect 38276 40832 38772 40866
rect 38276 40556 38310 40832
rect 38738 40770 38772 40832
rect 38738 40556 38772 40612
rect 38276 40516 38772 40556
rect 38276 40240 38310 40516
rect 38738 40460 38772 40516
rect 38738 40240 38772 40302
rect 38276 40206 38772 40240
rect 43266 40832 43762 40866
rect 43266 40556 43300 40832
rect 43728 40770 43762 40832
rect 43728 40556 43762 40612
rect 43266 40516 43762 40556
rect 43266 40240 43300 40516
rect 43728 40460 43762 40516
rect 43728 40240 43762 40302
rect 43266 40206 43762 40240
rect 48256 40832 48752 40866
rect 48256 40556 48290 40832
rect 48718 40770 48752 40832
rect 48718 40556 48752 40612
rect 48256 40516 48752 40556
rect 48256 40240 48290 40516
rect 48718 40460 48752 40516
rect 48718 40240 48752 40302
rect 48256 40206 48752 40240
rect 53246 40832 53742 40866
rect 53246 40556 53280 40832
rect 53708 40770 53742 40832
rect 53708 40556 53742 40612
rect 53246 40516 53742 40556
rect 53246 40240 53280 40516
rect 53708 40460 53742 40516
rect 53708 40240 53742 40302
rect 53246 40206 53742 40240
rect 58236 40832 58732 40866
rect 58236 40556 58270 40832
rect 58698 40770 58732 40832
rect 58698 40556 58732 40612
rect 58236 40516 58732 40556
rect 58236 40240 58270 40516
rect 58698 40460 58732 40516
rect 58698 40240 58732 40302
rect 58236 40206 58732 40240
rect 63226 40832 63722 40866
rect 63226 40556 63260 40832
rect 63688 40770 63722 40832
rect 63688 40556 63722 40612
rect 63226 40516 63722 40556
rect 63226 40240 63260 40516
rect 63688 40460 63722 40516
rect 63688 40240 63722 40302
rect 63226 40206 63722 40240
rect 68216 40832 68712 40866
rect 68216 40556 68250 40832
rect 68678 40770 68712 40832
rect 68678 40556 68712 40612
rect 68216 40516 68712 40556
rect 68216 40240 68250 40516
rect 68678 40460 68712 40516
rect 68678 40240 68712 40302
rect 68216 40206 68712 40240
rect 73206 40832 73702 40866
rect 73206 40556 73240 40832
rect 73668 40770 73702 40832
rect 73668 40556 73702 40612
rect 73206 40516 73702 40556
rect 73206 40240 73240 40516
rect 73668 40460 73702 40516
rect 73668 40240 73702 40302
rect 73206 40206 73702 40240
rect 78196 40832 78692 40866
rect 78196 40556 78230 40832
rect 78658 40770 78692 40832
rect 78658 40556 78692 40612
rect 78196 40516 78692 40556
rect 78196 40240 78230 40516
rect 78658 40460 78692 40516
rect 78658 40240 78692 40302
rect 78196 40206 78692 40240
<< psubdiffcont >>
rect 2786 66262 2820 66420
rect 2786 65952 2820 66110
rect 7776 66262 7810 66420
rect 7776 65952 7810 66110
rect 12766 66262 12800 66420
rect 12766 65952 12800 66110
rect 17756 66262 17790 66420
rect 17756 65952 17790 66110
rect 22746 66262 22780 66420
rect 22746 65952 22780 66110
rect 27736 66262 27770 66420
rect 27736 65952 27770 66110
rect 32726 66262 32760 66420
rect 32726 65952 32760 66110
rect 37716 66262 37750 66420
rect 37716 65952 37750 66110
rect 42706 66262 42740 66420
rect 42706 65952 42740 66110
rect 47696 66262 47730 66420
rect 47696 65952 47730 66110
rect 52686 66262 52720 66420
rect 52686 65952 52720 66110
rect 57676 66262 57710 66420
rect 57676 65952 57710 66110
rect 62666 66262 62700 66420
rect 62666 65952 62700 66110
rect 67656 66262 67690 66420
rect 67656 65952 67690 66110
rect 72646 66262 72680 66420
rect 72646 65952 72680 66110
rect 77636 66262 77670 66420
rect 77636 65952 77670 66110
rect 2786 64552 2820 64710
rect 2786 64242 2820 64400
rect 7776 64552 7810 64710
rect 7776 64242 7810 64400
rect 12766 64552 12800 64710
rect 12766 64242 12800 64400
rect 17756 64552 17790 64710
rect 17756 64242 17790 64400
rect 22746 64552 22780 64710
rect 22746 64242 22780 64400
rect 27736 64552 27770 64710
rect 27736 64242 27770 64400
rect 32726 64552 32760 64710
rect 32726 64242 32760 64400
rect 37716 64552 37750 64710
rect 37716 64242 37750 64400
rect 42706 64552 42740 64710
rect 42706 64242 42740 64400
rect 47696 64552 47730 64710
rect 47696 64242 47730 64400
rect 52686 64552 52720 64710
rect 52686 64242 52720 64400
rect 57676 64552 57710 64710
rect 57676 64242 57710 64400
rect 62666 64552 62700 64710
rect 62666 64242 62700 64400
rect 67656 64552 67690 64710
rect 67656 64242 67690 64400
rect 72646 64552 72680 64710
rect 72646 64242 72680 64400
rect 77636 64552 77670 64710
rect 77636 64242 77670 64400
rect 2786 62842 2820 63000
rect 2786 62532 2820 62690
rect 7776 62842 7810 63000
rect 7776 62532 7810 62690
rect 12766 62842 12800 63000
rect 12766 62532 12800 62690
rect 17756 62842 17790 63000
rect 17756 62532 17790 62690
rect 22746 62842 22780 63000
rect 22746 62532 22780 62690
rect 27736 62842 27770 63000
rect 27736 62532 27770 62690
rect 32726 62842 32760 63000
rect 32726 62532 32760 62690
rect 37716 62842 37750 63000
rect 37716 62532 37750 62690
rect 42706 62842 42740 63000
rect 42706 62532 42740 62690
rect 47696 62842 47730 63000
rect 47696 62532 47730 62690
rect 52686 62842 52720 63000
rect 52686 62532 52720 62690
rect 57676 62842 57710 63000
rect 57676 62532 57710 62690
rect 62666 62842 62700 63000
rect 62666 62532 62700 62690
rect 67656 62842 67690 63000
rect 67656 62532 67690 62690
rect 72646 62842 72680 63000
rect 72646 62532 72680 62690
rect 77636 62842 77670 63000
rect 77636 62532 77670 62690
rect 2786 61132 2820 61290
rect 2786 60822 2820 60980
rect 7776 61132 7810 61290
rect 7776 60822 7810 60980
rect 12766 61132 12800 61290
rect 12766 60822 12800 60980
rect 17756 61132 17790 61290
rect 17756 60822 17790 60980
rect 22746 61132 22780 61290
rect 22746 60822 22780 60980
rect 27736 61132 27770 61290
rect 27736 60822 27770 60980
rect 32726 61132 32760 61290
rect 32726 60822 32760 60980
rect 37716 61132 37750 61290
rect 37716 60822 37750 60980
rect 42706 61132 42740 61290
rect 42706 60822 42740 60980
rect 47696 61132 47730 61290
rect 47696 60822 47730 60980
rect 52686 61132 52720 61290
rect 52686 60822 52720 60980
rect 57676 61132 57710 61290
rect 57676 60822 57710 60980
rect 62666 61132 62700 61290
rect 62666 60822 62700 60980
rect 67656 61132 67690 61290
rect 67656 60822 67690 60980
rect 72646 61132 72680 61290
rect 72646 60822 72680 60980
rect 77636 61132 77670 61290
rect 77636 60822 77670 60980
rect 2786 59422 2820 59580
rect 2786 59112 2820 59270
rect 7776 59422 7810 59580
rect 7776 59112 7810 59270
rect 12766 59422 12800 59580
rect 12766 59112 12800 59270
rect 17756 59422 17790 59580
rect 17756 59112 17790 59270
rect 22746 59422 22780 59580
rect 22746 59112 22780 59270
rect 27736 59422 27770 59580
rect 27736 59112 27770 59270
rect 32726 59422 32760 59580
rect 32726 59112 32760 59270
rect 37716 59422 37750 59580
rect 37716 59112 37750 59270
rect 42706 59422 42740 59580
rect 42706 59112 42740 59270
rect 47696 59422 47730 59580
rect 47696 59112 47730 59270
rect 52686 59422 52720 59580
rect 52686 59112 52720 59270
rect 57676 59422 57710 59580
rect 57676 59112 57710 59270
rect 62666 59422 62700 59580
rect 62666 59112 62700 59270
rect 67656 59422 67690 59580
rect 67656 59112 67690 59270
rect 72646 59422 72680 59580
rect 72646 59112 72680 59270
rect 77636 59422 77670 59580
rect 77636 59112 77670 59270
rect 2786 57712 2820 57870
rect 2786 57402 2820 57560
rect 7776 57712 7810 57870
rect 7776 57402 7810 57560
rect 12766 57712 12800 57870
rect 12766 57402 12800 57560
rect 17756 57712 17790 57870
rect 17756 57402 17790 57560
rect 22746 57712 22780 57870
rect 22746 57402 22780 57560
rect 27736 57712 27770 57870
rect 27736 57402 27770 57560
rect 32726 57712 32760 57870
rect 32726 57402 32760 57560
rect 37716 57712 37750 57870
rect 37716 57402 37750 57560
rect 42706 57712 42740 57870
rect 42706 57402 42740 57560
rect 47696 57712 47730 57870
rect 47696 57402 47730 57560
rect 52686 57712 52720 57870
rect 52686 57402 52720 57560
rect 57676 57712 57710 57870
rect 57676 57402 57710 57560
rect 62666 57712 62700 57870
rect 62666 57402 62700 57560
rect 67656 57712 67690 57870
rect 67656 57402 67690 57560
rect 72646 57712 72680 57870
rect 72646 57402 72680 57560
rect 77636 57712 77670 57870
rect 77636 57402 77670 57560
rect 2786 56002 2820 56160
rect 2786 55692 2820 55850
rect 7776 56002 7810 56160
rect 7776 55692 7810 55850
rect 12766 56002 12800 56160
rect 12766 55692 12800 55850
rect 17756 56002 17790 56160
rect 17756 55692 17790 55850
rect 22746 56002 22780 56160
rect 22746 55692 22780 55850
rect 27736 56002 27770 56160
rect 27736 55692 27770 55850
rect 32726 56002 32760 56160
rect 32726 55692 32760 55850
rect 37716 56002 37750 56160
rect 37716 55692 37750 55850
rect 42706 56002 42740 56160
rect 42706 55692 42740 55850
rect 47696 56002 47730 56160
rect 47696 55692 47730 55850
rect 52686 56002 52720 56160
rect 52686 55692 52720 55850
rect 57676 56002 57710 56160
rect 57676 55692 57710 55850
rect 62666 56002 62700 56160
rect 62666 55692 62700 55850
rect 67656 56002 67690 56160
rect 67656 55692 67690 55850
rect 72646 56002 72680 56160
rect 72646 55692 72680 55850
rect 77636 56002 77670 56160
rect 77636 55692 77670 55850
rect 2786 54292 2820 54450
rect 2786 53982 2820 54140
rect 7776 54292 7810 54450
rect 7776 53982 7810 54140
rect 12766 54292 12800 54450
rect 12766 53982 12800 54140
rect 17756 54292 17790 54450
rect 17756 53982 17790 54140
rect 22746 54292 22780 54450
rect 22746 53982 22780 54140
rect 27736 54292 27770 54450
rect 27736 53982 27770 54140
rect 32726 54292 32760 54450
rect 32726 53982 32760 54140
rect 37716 54292 37750 54450
rect 37716 53982 37750 54140
rect 42706 54292 42740 54450
rect 42706 53982 42740 54140
rect 47696 54292 47730 54450
rect 47696 53982 47730 54140
rect 52686 54292 52720 54450
rect 52686 53982 52720 54140
rect 57676 54292 57710 54450
rect 57676 53982 57710 54140
rect 62666 54292 62700 54450
rect 62666 53982 62700 54140
rect 67656 54292 67690 54450
rect 67656 53982 67690 54140
rect 72646 54292 72680 54450
rect 72646 53982 72680 54140
rect 77636 54292 77670 54450
rect 77636 53982 77670 54140
rect 2786 52582 2820 52740
rect 2786 52272 2820 52430
rect 7776 52582 7810 52740
rect 7776 52272 7810 52430
rect 12766 52582 12800 52740
rect 12766 52272 12800 52430
rect 17756 52582 17790 52740
rect 17756 52272 17790 52430
rect 22746 52582 22780 52740
rect 22746 52272 22780 52430
rect 27736 52582 27770 52740
rect 27736 52272 27770 52430
rect 32726 52582 32760 52740
rect 32726 52272 32760 52430
rect 37716 52582 37750 52740
rect 37716 52272 37750 52430
rect 42706 52582 42740 52740
rect 42706 52272 42740 52430
rect 47696 52582 47730 52740
rect 47696 52272 47730 52430
rect 52686 52582 52720 52740
rect 52686 52272 52720 52430
rect 57676 52582 57710 52740
rect 57676 52272 57710 52430
rect 62666 52582 62700 52740
rect 62666 52272 62700 52430
rect 67656 52582 67690 52740
rect 67656 52272 67690 52430
rect 72646 52582 72680 52740
rect 72646 52272 72680 52430
rect 77636 52582 77670 52740
rect 77636 52272 77670 52430
rect 2786 50872 2820 51030
rect 2786 50562 2820 50720
rect 7776 50872 7810 51030
rect 7776 50562 7810 50720
rect 12766 50872 12800 51030
rect 12766 50562 12800 50720
rect 17756 50872 17790 51030
rect 17756 50562 17790 50720
rect 22746 50872 22780 51030
rect 22746 50562 22780 50720
rect 27736 50872 27770 51030
rect 27736 50562 27770 50720
rect 32726 50872 32760 51030
rect 32726 50562 32760 50720
rect 37716 50872 37750 51030
rect 37716 50562 37750 50720
rect 42706 50872 42740 51030
rect 42706 50562 42740 50720
rect 47696 50872 47730 51030
rect 47696 50562 47730 50720
rect 52686 50872 52720 51030
rect 52686 50562 52720 50720
rect 57676 50872 57710 51030
rect 57676 50562 57710 50720
rect 62666 50872 62700 51030
rect 62666 50562 62700 50720
rect 67656 50872 67690 51030
rect 67656 50562 67690 50720
rect 72646 50872 72680 51030
rect 72646 50562 72680 50720
rect 77636 50872 77670 51030
rect 77636 50562 77670 50720
rect 2786 49162 2820 49320
rect 2786 48852 2820 49010
rect 7776 49162 7810 49320
rect 7776 48852 7810 49010
rect 12766 49162 12800 49320
rect 12766 48852 12800 49010
rect 17756 49162 17790 49320
rect 17756 48852 17790 49010
rect 22746 49162 22780 49320
rect 22746 48852 22780 49010
rect 27736 49162 27770 49320
rect 27736 48852 27770 49010
rect 32726 49162 32760 49320
rect 32726 48852 32760 49010
rect 37716 49162 37750 49320
rect 37716 48852 37750 49010
rect 42706 49162 42740 49320
rect 42706 48852 42740 49010
rect 47696 49162 47730 49320
rect 47696 48852 47730 49010
rect 52686 49162 52720 49320
rect 52686 48852 52720 49010
rect 57676 49162 57710 49320
rect 57676 48852 57710 49010
rect 62666 49162 62700 49320
rect 62666 48852 62700 49010
rect 67656 49162 67690 49320
rect 67656 48852 67690 49010
rect 72646 49162 72680 49320
rect 72646 48852 72680 49010
rect 77636 49162 77670 49320
rect 77636 48852 77670 49010
rect 2786 47452 2820 47610
rect 2786 47142 2820 47300
rect 7776 47452 7810 47610
rect 7776 47142 7810 47300
rect 12766 47452 12800 47610
rect 12766 47142 12800 47300
rect 17756 47452 17790 47610
rect 17756 47142 17790 47300
rect 22746 47452 22780 47610
rect 22746 47142 22780 47300
rect 27736 47452 27770 47610
rect 27736 47142 27770 47300
rect 32726 47452 32760 47610
rect 32726 47142 32760 47300
rect 37716 47452 37750 47610
rect 37716 47142 37750 47300
rect 42706 47452 42740 47610
rect 42706 47142 42740 47300
rect 47696 47452 47730 47610
rect 47696 47142 47730 47300
rect 52686 47452 52720 47610
rect 52686 47142 52720 47300
rect 57676 47452 57710 47610
rect 57676 47142 57710 47300
rect 62666 47452 62700 47610
rect 62666 47142 62700 47300
rect 67656 47452 67690 47610
rect 67656 47142 67690 47300
rect 72646 47452 72680 47610
rect 72646 47142 72680 47300
rect 77636 47452 77670 47610
rect 77636 47142 77670 47300
rect 2786 45742 2820 45900
rect 2786 45432 2820 45590
rect 7776 45742 7810 45900
rect 7776 45432 7810 45590
rect 12766 45742 12800 45900
rect 12766 45432 12800 45590
rect 17756 45742 17790 45900
rect 17756 45432 17790 45590
rect 22746 45742 22780 45900
rect 22746 45432 22780 45590
rect 27736 45742 27770 45900
rect 27736 45432 27770 45590
rect 32726 45742 32760 45900
rect 32726 45432 32760 45590
rect 37716 45742 37750 45900
rect 37716 45432 37750 45590
rect 42706 45742 42740 45900
rect 42706 45432 42740 45590
rect 47696 45742 47730 45900
rect 47696 45432 47730 45590
rect 52686 45742 52720 45900
rect 52686 45432 52720 45590
rect 57676 45742 57710 45900
rect 57676 45432 57710 45590
rect 62666 45742 62700 45900
rect 62666 45432 62700 45590
rect 67656 45742 67690 45900
rect 67656 45432 67690 45590
rect 72646 45742 72680 45900
rect 72646 45432 72680 45590
rect 77636 45742 77670 45900
rect 77636 45432 77670 45590
rect 2786 44032 2820 44190
rect 2786 43722 2820 43880
rect 7776 44032 7810 44190
rect 7776 43722 7810 43880
rect 12766 44032 12800 44190
rect 12766 43722 12800 43880
rect 17756 44032 17790 44190
rect 17756 43722 17790 43880
rect 22746 44032 22780 44190
rect 22746 43722 22780 43880
rect 27736 44032 27770 44190
rect 27736 43722 27770 43880
rect 32726 44032 32760 44190
rect 32726 43722 32760 43880
rect 37716 44032 37750 44190
rect 37716 43722 37750 43880
rect 42706 44032 42740 44190
rect 42706 43722 42740 43880
rect 47696 44032 47730 44190
rect 47696 43722 47730 43880
rect 52686 44032 52720 44190
rect 52686 43722 52720 43880
rect 57676 44032 57710 44190
rect 57676 43722 57710 43880
rect 62666 44032 62700 44190
rect 62666 43722 62700 43880
rect 67656 44032 67690 44190
rect 67656 43722 67690 43880
rect 72646 44032 72680 44190
rect 72646 43722 72680 43880
rect 77636 44032 77670 44190
rect 77636 43722 77670 43880
rect 2786 42322 2820 42480
rect 2786 42012 2820 42170
rect 7776 42322 7810 42480
rect 7776 42012 7810 42170
rect 12766 42322 12800 42480
rect 12766 42012 12800 42170
rect 17756 42322 17790 42480
rect 17756 42012 17790 42170
rect 22746 42322 22780 42480
rect 22746 42012 22780 42170
rect 27736 42322 27770 42480
rect 27736 42012 27770 42170
rect 32726 42322 32760 42480
rect 32726 42012 32760 42170
rect 37716 42322 37750 42480
rect 37716 42012 37750 42170
rect 42706 42322 42740 42480
rect 42706 42012 42740 42170
rect 47696 42322 47730 42480
rect 47696 42012 47730 42170
rect 52686 42322 52720 42480
rect 52686 42012 52720 42170
rect 57676 42322 57710 42480
rect 57676 42012 57710 42170
rect 62666 42322 62700 42480
rect 62666 42012 62700 42170
rect 67656 42322 67690 42480
rect 67656 42012 67690 42170
rect 72646 42322 72680 42480
rect 72646 42012 72680 42170
rect 77636 42322 77670 42480
rect 77636 42012 77670 42170
rect 2786 40612 2820 40770
rect 2786 40302 2820 40460
rect 7776 40612 7810 40770
rect 7776 40302 7810 40460
rect 12766 40612 12800 40770
rect 12766 40302 12800 40460
rect 17756 40612 17790 40770
rect 17756 40302 17790 40460
rect 22746 40612 22780 40770
rect 22746 40302 22780 40460
rect 27736 40612 27770 40770
rect 27736 40302 27770 40460
rect 32726 40612 32760 40770
rect 32726 40302 32760 40460
rect 37716 40612 37750 40770
rect 37716 40302 37750 40460
rect 42706 40612 42740 40770
rect 42706 40302 42740 40460
rect 47696 40612 47730 40770
rect 47696 40302 47730 40460
rect 52686 40612 52720 40770
rect 52686 40302 52720 40460
rect 57676 40612 57710 40770
rect 57676 40302 57710 40460
rect 62666 40612 62700 40770
rect 62666 40302 62700 40460
rect 67656 40612 67690 40770
rect 67656 40302 67690 40460
rect 72646 40612 72680 40770
rect 72646 40302 72680 40460
rect 77636 40612 77670 40770
rect 77636 40302 77670 40460
<< nsubdiffcont >>
rect 3808 66262 3842 66420
rect 3808 65952 3842 66110
rect 8798 66262 8832 66420
rect 8798 65952 8832 66110
rect 13788 66262 13822 66420
rect 13788 65952 13822 66110
rect 18778 66262 18812 66420
rect 18778 65952 18812 66110
rect 23768 66262 23802 66420
rect 23768 65952 23802 66110
rect 28758 66262 28792 66420
rect 28758 65952 28792 66110
rect 33748 66262 33782 66420
rect 33748 65952 33782 66110
rect 38738 66262 38772 66420
rect 38738 65952 38772 66110
rect 43728 66262 43762 66420
rect 43728 65952 43762 66110
rect 48718 66262 48752 66420
rect 48718 65952 48752 66110
rect 53708 66262 53742 66420
rect 53708 65952 53742 66110
rect 58698 66262 58732 66420
rect 58698 65952 58732 66110
rect 63688 66262 63722 66420
rect 63688 65952 63722 66110
rect 68678 66262 68712 66420
rect 68678 65952 68712 66110
rect 73668 66262 73702 66420
rect 73668 65952 73702 66110
rect 78658 66262 78692 66420
rect 78658 65952 78692 66110
rect 3808 64552 3842 64710
rect 3808 64242 3842 64400
rect 8798 64552 8832 64710
rect 8798 64242 8832 64400
rect 13788 64552 13822 64710
rect 13788 64242 13822 64400
rect 18778 64552 18812 64710
rect 18778 64242 18812 64400
rect 23768 64552 23802 64710
rect 23768 64242 23802 64400
rect 28758 64552 28792 64710
rect 28758 64242 28792 64400
rect 33748 64552 33782 64710
rect 33748 64242 33782 64400
rect 38738 64552 38772 64710
rect 38738 64242 38772 64400
rect 43728 64552 43762 64710
rect 43728 64242 43762 64400
rect 48718 64552 48752 64710
rect 48718 64242 48752 64400
rect 53708 64552 53742 64710
rect 53708 64242 53742 64400
rect 58698 64552 58732 64710
rect 58698 64242 58732 64400
rect 63688 64552 63722 64710
rect 63688 64242 63722 64400
rect 68678 64552 68712 64710
rect 68678 64242 68712 64400
rect 73668 64552 73702 64710
rect 73668 64242 73702 64400
rect 78658 64552 78692 64710
rect 78658 64242 78692 64400
rect 3808 62842 3842 63000
rect 3808 62532 3842 62690
rect 8798 62842 8832 63000
rect 8798 62532 8832 62690
rect 13788 62842 13822 63000
rect 13788 62532 13822 62690
rect 18778 62842 18812 63000
rect 18778 62532 18812 62690
rect 23768 62842 23802 63000
rect 23768 62532 23802 62690
rect 28758 62842 28792 63000
rect 28758 62532 28792 62690
rect 33748 62842 33782 63000
rect 33748 62532 33782 62690
rect 38738 62842 38772 63000
rect 38738 62532 38772 62690
rect 43728 62842 43762 63000
rect 43728 62532 43762 62690
rect 48718 62842 48752 63000
rect 48718 62532 48752 62690
rect 53708 62842 53742 63000
rect 53708 62532 53742 62690
rect 58698 62842 58732 63000
rect 58698 62532 58732 62690
rect 63688 62842 63722 63000
rect 63688 62532 63722 62690
rect 68678 62842 68712 63000
rect 68678 62532 68712 62690
rect 73668 62842 73702 63000
rect 73668 62532 73702 62690
rect 78658 62842 78692 63000
rect 78658 62532 78692 62690
rect 3808 61132 3842 61290
rect 3808 60822 3842 60980
rect 8798 61132 8832 61290
rect 8798 60822 8832 60980
rect 13788 61132 13822 61290
rect 13788 60822 13822 60980
rect 18778 61132 18812 61290
rect 18778 60822 18812 60980
rect 23768 61132 23802 61290
rect 23768 60822 23802 60980
rect 28758 61132 28792 61290
rect 28758 60822 28792 60980
rect 33748 61132 33782 61290
rect 33748 60822 33782 60980
rect 38738 61132 38772 61290
rect 38738 60822 38772 60980
rect 43728 61132 43762 61290
rect 43728 60822 43762 60980
rect 48718 61132 48752 61290
rect 48718 60822 48752 60980
rect 53708 61132 53742 61290
rect 53708 60822 53742 60980
rect 58698 61132 58732 61290
rect 58698 60822 58732 60980
rect 63688 61132 63722 61290
rect 63688 60822 63722 60980
rect 68678 61132 68712 61290
rect 68678 60822 68712 60980
rect 73668 61132 73702 61290
rect 73668 60822 73702 60980
rect 78658 61132 78692 61290
rect 78658 60822 78692 60980
rect 3808 59422 3842 59580
rect 3808 59112 3842 59270
rect 8798 59422 8832 59580
rect 8798 59112 8832 59270
rect 13788 59422 13822 59580
rect 13788 59112 13822 59270
rect 18778 59422 18812 59580
rect 18778 59112 18812 59270
rect 23768 59422 23802 59580
rect 23768 59112 23802 59270
rect 28758 59422 28792 59580
rect 28758 59112 28792 59270
rect 33748 59422 33782 59580
rect 33748 59112 33782 59270
rect 38738 59422 38772 59580
rect 38738 59112 38772 59270
rect 43728 59422 43762 59580
rect 43728 59112 43762 59270
rect 48718 59422 48752 59580
rect 48718 59112 48752 59270
rect 53708 59422 53742 59580
rect 53708 59112 53742 59270
rect 58698 59422 58732 59580
rect 58698 59112 58732 59270
rect 63688 59422 63722 59580
rect 63688 59112 63722 59270
rect 68678 59422 68712 59580
rect 68678 59112 68712 59270
rect 73668 59422 73702 59580
rect 73668 59112 73702 59270
rect 78658 59422 78692 59580
rect 78658 59112 78692 59270
rect 3808 57712 3842 57870
rect 3808 57402 3842 57560
rect 8798 57712 8832 57870
rect 8798 57402 8832 57560
rect 13788 57712 13822 57870
rect 13788 57402 13822 57560
rect 18778 57712 18812 57870
rect 18778 57402 18812 57560
rect 23768 57712 23802 57870
rect 23768 57402 23802 57560
rect 28758 57712 28792 57870
rect 28758 57402 28792 57560
rect 33748 57712 33782 57870
rect 33748 57402 33782 57560
rect 38738 57712 38772 57870
rect 38738 57402 38772 57560
rect 43728 57712 43762 57870
rect 43728 57402 43762 57560
rect 48718 57712 48752 57870
rect 48718 57402 48752 57560
rect 53708 57712 53742 57870
rect 53708 57402 53742 57560
rect 58698 57712 58732 57870
rect 58698 57402 58732 57560
rect 63688 57712 63722 57870
rect 63688 57402 63722 57560
rect 68678 57712 68712 57870
rect 68678 57402 68712 57560
rect 73668 57712 73702 57870
rect 73668 57402 73702 57560
rect 78658 57712 78692 57870
rect 78658 57402 78692 57560
rect 3808 56002 3842 56160
rect 3808 55692 3842 55850
rect 8798 56002 8832 56160
rect 8798 55692 8832 55850
rect 13788 56002 13822 56160
rect 13788 55692 13822 55850
rect 18778 56002 18812 56160
rect 18778 55692 18812 55850
rect 23768 56002 23802 56160
rect 23768 55692 23802 55850
rect 28758 56002 28792 56160
rect 28758 55692 28792 55850
rect 33748 56002 33782 56160
rect 33748 55692 33782 55850
rect 38738 56002 38772 56160
rect 38738 55692 38772 55850
rect 43728 56002 43762 56160
rect 43728 55692 43762 55850
rect 48718 56002 48752 56160
rect 48718 55692 48752 55850
rect 53708 56002 53742 56160
rect 53708 55692 53742 55850
rect 58698 56002 58732 56160
rect 58698 55692 58732 55850
rect 63688 56002 63722 56160
rect 63688 55692 63722 55850
rect 68678 56002 68712 56160
rect 68678 55692 68712 55850
rect 73668 56002 73702 56160
rect 73668 55692 73702 55850
rect 78658 56002 78692 56160
rect 78658 55692 78692 55850
rect 3808 54292 3842 54450
rect 3808 53982 3842 54140
rect 8798 54292 8832 54450
rect 8798 53982 8832 54140
rect 13788 54292 13822 54450
rect 13788 53982 13822 54140
rect 18778 54292 18812 54450
rect 18778 53982 18812 54140
rect 23768 54292 23802 54450
rect 23768 53982 23802 54140
rect 28758 54292 28792 54450
rect 28758 53982 28792 54140
rect 33748 54292 33782 54450
rect 33748 53982 33782 54140
rect 38738 54292 38772 54450
rect 38738 53982 38772 54140
rect 43728 54292 43762 54450
rect 43728 53982 43762 54140
rect 48718 54292 48752 54450
rect 48718 53982 48752 54140
rect 53708 54292 53742 54450
rect 53708 53982 53742 54140
rect 58698 54292 58732 54450
rect 58698 53982 58732 54140
rect 63688 54292 63722 54450
rect 63688 53982 63722 54140
rect 68678 54292 68712 54450
rect 68678 53982 68712 54140
rect 73668 54292 73702 54450
rect 73668 53982 73702 54140
rect 78658 54292 78692 54450
rect 78658 53982 78692 54140
rect 3808 52582 3842 52740
rect 3808 52272 3842 52430
rect 8798 52582 8832 52740
rect 8798 52272 8832 52430
rect 13788 52582 13822 52740
rect 13788 52272 13822 52430
rect 18778 52582 18812 52740
rect 18778 52272 18812 52430
rect 23768 52582 23802 52740
rect 23768 52272 23802 52430
rect 28758 52582 28792 52740
rect 28758 52272 28792 52430
rect 33748 52582 33782 52740
rect 33748 52272 33782 52430
rect 38738 52582 38772 52740
rect 38738 52272 38772 52430
rect 43728 52582 43762 52740
rect 43728 52272 43762 52430
rect 48718 52582 48752 52740
rect 48718 52272 48752 52430
rect 53708 52582 53742 52740
rect 53708 52272 53742 52430
rect 58698 52582 58732 52740
rect 58698 52272 58732 52430
rect 63688 52582 63722 52740
rect 63688 52272 63722 52430
rect 68678 52582 68712 52740
rect 68678 52272 68712 52430
rect 73668 52582 73702 52740
rect 73668 52272 73702 52430
rect 78658 52582 78692 52740
rect 78658 52272 78692 52430
rect 3808 50872 3842 51030
rect 3808 50562 3842 50720
rect 8798 50872 8832 51030
rect 8798 50562 8832 50720
rect 13788 50872 13822 51030
rect 13788 50562 13822 50720
rect 18778 50872 18812 51030
rect 18778 50562 18812 50720
rect 23768 50872 23802 51030
rect 23768 50562 23802 50720
rect 28758 50872 28792 51030
rect 28758 50562 28792 50720
rect 33748 50872 33782 51030
rect 33748 50562 33782 50720
rect 38738 50872 38772 51030
rect 38738 50562 38772 50720
rect 43728 50872 43762 51030
rect 43728 50562 43762 50720
rect 48718 50872 48752 51030
rect 48718 50562 48752 50720
rect 53708 50872 53742 51030
rect 53708 50562 53742 50720
rect 58698 50872 58732 51030
rect 58698 50562 58732 50720
rect 63688 50872 63722 51030
rect 63688 50562 63722 50720
rect 68678 50872 68712 51030
rect 68678 50562 68712 50720
rect 73668 50872 73702 51030
rect 73668 50562 73702 50720
rect 78658 50872 78692 51030
rect 78658 50562 78692 50720
rect 3808 49162 3842 49320
rect 3808 48852 3842 49010
rect 8798 49162 8832 49320
rect 8798 48852 8832 49010
rect 13788 49162 13822 49320
rect 13788 48852 13822 49010
rect 18778 49162 18812 49320
rect 18778 48852 18812 49010
rect 23768 49162 23802 49320
rect 23768 48852 23802 49010
rect 28758 49162 28792 49320
rect 28758 48852 28792 49010
rect 33748 49162 33782 49320
rect 33748 48852 33782 49010
rect 38738 49162 38772 49320
rect 38738 48852 38772 49010
rect 43728 49162 43762 49320
rect 43728 48852 43762 49010
rect 48718 49162 48752 49320
rect 48718 48852 48752 49010
rect 53708 49162 53742 49320
rect 53708 48852 53742 49010
rect 58698 49162 58732 49320
rect 58698 48852 58732 49010
rect 63688 49162 63722 49320
rect 63688 48852 63722 49010
rect 68678 49162 68712 49320
rect 68678 48852 68712 49010
rect 73668 49162 73702 49320
rect 73668 48852 73702 49010
rect 78658 49162 78692 49320
rect 78658 48852 78692 49010
rect 3808 47452 3842 47610
rect 3808 47142 3842 47300
rect 8798 47452 8832 47610
rect 8798 47142 8832 47300
rect 13788 47452 13822 47610
rect 13788 47142 13822 47300
rect 18778 47452 18812 47610
rect 18778 47142 18812 47300
rect 23768 47452 23802 47610
rect 23768 47142 23802 47300
rect 28758 47452 28792 47610
rect 28758 47142 28792 47300
rect 33748 47452 33782 47610
rect 33748 47142 33782 47300
rect 38738 47452 38772 47610
rect 38738 47142 38772 47300
rect 43728 47452 43762 47610
rect 43728 47142 43762 47300
rect 48718 47452 48752 47610
rect 48718 47142 48752 47300
rect 53708 47452 53742 47610
rect 53708 47142 53742 47300
rect 58698 47452 58732 47610
rect 58698 47142 58732 47300
rect 63688 47452 63722 47610
rect 63688 47142 63722 47300
rect 68678 47452 68712 47610
rect 68678 47142 68712 47300
rect 73668 47452 73702 47610
rect 73668 47142 73702 47300
rect 78658 47452 78692 47610
rect 78658 47142 78692 47300
rect 3808 45742 3842 45900
rect 3808 45432 3842 45590
rect 8798 45742 8832 45900
rect 8798 45432 8832 45590
rect 13788 45742 13822 45900
rect 13788 45432 13822 45590
rect 18778 45742 18812 45900
rect 18778 45432 18812 45590
rect 23768 45742 23802 45900
rect 23768 45432 23802 45590
rect 28758 45742 28792 45900
rect 28758 45432 28792 45590
rect 33748 45742 33782 45900
rect 33748 45432 33782 45590
rect 38738 45742 38772 45900
rect 38738 45432 38772 45590
rect 43728 45742 43762 45900
rect 43728 45432 43762 45590
rect 48718 45742 48752 45900
rect 48718 45432 48752 45590
rect 53708 45742 53742 45900
rect 53708 45432 53742 45590
rect 58698 45742 58732 45900
rect 58698 45432 58732 45590
rect 63688 45742 63722 45900
rect 63688 45432 63722 45590
rect 68678 45742 68712 45900
rect 68678 45432 68712 45590
rect 73668 45742 73702 45900
rect 73668 45432 73702 45590
rect 78658 45742 78692 45900
rect 78658 45432 78692 45590
rect 3808 44032 3842 44190
rect 3808 43722 3842 43880
rect 8798 44032 8832 44190
rect 8798 43722 8832 43880
rect 13788 44032 13822 44190
rect 13788 43722 13822 43880
rect 18778 44032 18812 44190
rect 18778 43722 18812 43880
rect 23768 44032 23802 44190
rect 23768 43722 23802 43880
rect 28758 44032 28792 44190
rect 28758 43722 28792 43880
rect 33748 44032 33782 44190
rect 33748 43722 33782 43880
rect 38738 44032 38772 44190
rect 38738 43722 38772 43880
rect 43728 44032 43762 44190
rect 43728 43722 43762 43880
rect 48718 44032 48752 44190
rect 48718 43722 48752 43880
rect 53708 44032 53742 44190
rect 53708 43722 53742 43880
rect 58698 44032 58732 44190
rect 58698 43722 58732 43880
rect 63688 44032 63722 44190
rect 63688 43722 63722 43880
rect 68678 44032 68712 44190
rect 68678 43722 68712 43880
rect 73668 44032 73702 44190
rect 73668 43722 73702 43880
rect 78658 44032 78692 44190
rect 78658 43722 78692 43880
rect 3808 42322 3842 42480
rect 3808 42012 3842 42170
rect 8798 42322 8832 42480
rect 8798 42012 8832 42170
rect 13788 42322 13822 42480
rect 13788 42012 13822 42170
rect 18778 42322 18812 42480
rect 18778 42012 18812 42170
rect 23768 42322 23802 42480
rect 23768 42012 23802 42170
rect 28758 42322 28792 42480
rect 28758 42012 28792 42170
rect 33748 42322 33782 42480
rect 33748 42012 33782 42170
rect 38738 42322 38772 42480
rect 38738 42012 38772 42170
rect 43728 42322 43762 42480
rect 43728 42012 43762 42170
rect 48718 42322 48752 42480
rect 48718 42012 48752 42170
rect 53708 42322 53742 42480
rect 53708 42012 53742 42170
rect 58698 42322 58732 42480
rect 58698 42012 58732 42170
rect 63688 42322 63722 42480
rect 63688 42012 63722 42170
rect 68678 42322 68712 42480
rect 68678 42012 68712 42170
rect 73668 42322 73702 42480
rect 73668 42012 73702 42170
rect 78658 42322 78692 42480
rect 78658 42012 78692 42170
rect 3808 40612 3842 40770
rect 3808 40302 3842 40460
rect 8798 40612 8832 40770
rect 8798 40302 8832 40460
rect 13788 40612 13822 40770
rect 13788 40302 13822 40460
rect 18778 40612 18812 40770
rect 18778 40302 18812 40460
rect 23768 40612 23802 40770
rect 23768 40302 23802 40460
rect 28758 40612 28792 40770
rect 28758 40302 28792 40460
rect 33748 40612 33782 40770
rect 33748 40302 33782 40460
rect 38738 40612 38772 40770
rect 38738 40302 38772 40460
rect 43728 40612 43762 40770
rect 43728 40302 43762 40460
rect 48718 40612 48752 40770
rect 48718 40302 48752 40460
rect 53708 40612 53742 40770
rect 53708 40302 53742 40460
rect 58698 40612 58732 40770
rect 58698 40302 58732 40460
rect 63688 40612 63722 40770
rect 63688 40302 63722 40460
rect 68678 40612 68712 40770
rect 68678 40302 68712 40460
rect 73668 40612 73702 40770
rect 73668 40302 73702 40460
rect 78658 40612 78692 40770
rect 78658 40302 78692 40460
<< poly >>
rect 2872 66358 2938 66374
rect 2872 66324 2888 66358
rect 2922 66356 2938 66358
rect 2922 66326 2960 66356
rect 3160 66326 3186 66356
rect 2922 66324 2938 66326
rect 2872 66308 2938 66324
rect 2872 66048 2938 66064
rect 2872 66014 2888 66048
rect 2922 66046 2938 66048
rect 2922 66016 2960 66046
rect 3160 66016 3186 66046
rect 2922 66014 2938 66016
rect 2872 65998 2938 66014
rect 3689 66358 3755 66374
rect 3689 66356 3705 66358
rect 3432 66326 3458 66356
rect 3658 66326 3705 66356
rect 3689 66324 3705 66326
rect 3739 66324 3755 66358
rect 3689 66308 3755 66324
rect 3689 66048 3755 66064
rect 3689 66046 3705 66048
rect 3432 66016 3458 66046
rect 3658 66016 3705 66046
rect 3689 66014 3705 66016
rect 3739 66014 3755 66048
rect 3689 65998 3755 66014
rect 7862 66358 7928 66374
rect 7862 66324 7878 66358
rect 7912 66356 7928 66358
rect 7912 66326 7950 66356
rect 8150 66326 8176 66356
rect 7912 66324 7928 66326
rect 7862 66308 7928 66324
rect 7862 66048 7928 66064
rect 7862 66014 7878 66048
rect 7912 66046 7928 66048
rect 7912 66016 7950 66046
rect 8150 66016 8176 66046
rect 7912 66014 7928 66016
rect 7862 65998 7928 66014
rect 8679 66358 8745 66374
rect 8679 66356 8695 66358
rect 8422 66326 8448 66356
rect 8648 66326 8695 66356
rect 8679 66324 8695 66326
rect 8729 66324 8745 66358
rect 8679 66308 8745 66324
rect 8679 66048 8745 66064
rect 8679 66046 8695 66048
rect 8422 66016 8448 66046
rect 8648 66016 8695 66046
rect 8679 66014 8695 66016
rect 8729 66014 8745 66048
rect 8679 65998 8745 66014
rect 12852 66358 12918 66374
rect 12852 66324 12868 66358
rect 12902 66356 12918 66358
rect 12902 66326 12940 66356
rect 13140 66326 13166 66356
rect 12902 66324 12918 66326
rect 12852 66308 12918 66324
rect 12852 66048 12918 66064
rect 12852 66014 12868 66048
rect 12902 66046 12918 66048
rect 12902 66016 12940 66046
rect 13140 66016 13166 66046
rect 12902 66014 12918 66016
rect 12852 65998 12918 66014
rect 13669 66358 13735 66374
rect 13669 66356 13685 66358
rect 13412 66326 13438 66356
rect 13638 66326 13685 66356
rect 13669 66324 13685 66326
rect 13719 66324 13735 66358
rect 13669 66308 13735 66324
rect 13669 66048 13735 66064
rect 13669 66046 13685 66048
rect 13412 66016 13438 66046
rect 13638 66016 13685 66046
rect 13669 66014 13685 66016
rect 13719 66014 13735 66048
rect 13669 65998 13735 66014
rect 17842 66358 17908 66374
rect 17842 66324 17858 66358
rect 17892 66356 17908 66358
rect 17892 66326 17930 66356
rect 18130 66326 18156 66356
rect 17892 66324 17908 66326
rect 17842 66308 17908 66324
rect 17842 66048 17908 66064
rect 17842 66014 17858 66048
rect 17892 66046 17908 66048
rect 17892 66016 17930 66046
rect 18130 66016 18156 66046
rect 17892 66014 17908 66016
rect 17842 65998 17908 66014
rect 18659 66358 18725 66374
rect 18659 66356 18675 66358
rect 18402 66326 18428 66356
rect 18628 66326 18675 66356
rect 18659 66324 18675 66326
rect 18709 66324 18725 66358
rect 18659 66308 18725 66324
rect 18659 66048 18725 66064
rect 18659 66046 18675 66048
rect 18402 66016 18428 66046
rect 18628 66016 18675 66046
rect 18659 66014 18675 66016
rect 18709 66014 18725 66048
rect 18659 65998 18725 66014
rect 22832 66358 22898 66374
rect 22832 66324 22848 66358
rect 22882 66356 22898 66358
rect 22882 66326 22920 66356
rect 23120 66326 23146 66356
rect 22882 66324 22898 66326
rect 22832 66308 22898 66324
rect 22832 66048 22898 66064
rect 22832 66014 22848 66048
rect 22882 66046 22898 66048
rect 22882 66016 22920 66046
rect 23120 66016 23146 66046
rect 22882 66014 22898 66016
rect 22832 65998 22898 66014
rect 23649 66358 23715 66374
rect 23649 66356 23665 66358
rect 23392 66326 23418 66356
rect 23618 66326 23665 66356
rect 23649 66324 23665 66326
rect 23699 66324 23715 66358
rect 23649 66308 23715 66324
rect 23649 66048 23715 66064
rect 23649 66046 23665 66048
rect 23392 66016 23418 66046
rect 23618 66016 23665 66046
rect 23649 66014 23665 66016
rect 23699 66014 23715 66048
rect 23649 65998 23715 66014
rect 27822 66358 27888 66374
rect 27822 66324 27838 66358
rect 27872 66356 27888 66358
rect 27872 66326 27910 66356
rect 28110 66326 28136 66356
rect 27872 66324 27888 66326
rect 27822 66308 27888 66324
rect 27822 66048 27888 66064
rect 27822 66014 27838 66048
rect 27872 66046 27888 66048
rect 27872 66016 27910 66046
rect 28110 66016 28136 66046
rect 27872 66014 27888 66016
rect 27822 65998 27888 66014
rect 28639 66358 28705 66374
rect 28639 66356 28655 66358
rect 28382 66326 28408 66356
rect 28608 66326 28655 66356
rect 28639 66324 28655 66326
rect 28689 66324 28705 66358
rect 28639 66308 28705 66324
rect 28639 66048 28705 66064
rect 28639 66046 28655 66048
rect 28382 66016 28408 66046
rect 28608 66016 28655 66046
rect 28639 66014 28655 66016
rect 28689 66014 28705 66048
rect 28639 65998 28705 66014
rect 32812 66358 32878 66374
rect 32812 66324 32828 66358
rect 32862 66356 32878 66358
rect 32862 66326 32900 66356
rect 33100 66326 33126 66356
rect 32862 66324 32878 66326
rect 32812 66308 32878 66324
rect 32812 66048 32878 66064
rect 32812 66014 32828 66048
rect 32862 66046 32878 66048
rect 32862 66016 32900 66046
rect 33100 66016 33126 66046
rect 32862 66014 32878 66016
rect 32812 65998 32878 66014
rect 33629 66358 33695 66374
rect 33629 66356 33645 66358
rect 33372 66326 33398 66356
rect 33598 66326 33645 66356
rect 33629 66324 33645 66326
rect 33679 66324 33695 66358
rect 33629 66308 33695 66324
rect 33629 66048 33695 66064
rect 33629 66046 33645 66048
rect 33372 66016 33398 66046
rect 33598 66016 33645 66046
rect 33629 66014 33645 66016
rect 33679 66014 33695 66048
rect 33629 65998 33695 66014
rect 37802 66358 37868 66374
rect 37802 66324 37818 66358
rect 37852 66356 37868 66358
rect 37852 66326 37890 66356
rect 38090 66326 38116 66356
rect 37852 66324 37868 66326
rect 37802 66308 37868 66324
rect 37802 66048 37868 66064
rect 37802 66014 37818 66048
rect 37852 66046 37868 66048
rect 37852 66016 37890 66046
rect 38090 66016 38116 66046
rect 37852 66014 37868 66016
rect 37802 65998 37868 66014
rect 38619 66358 38685 66374
rect 38619 66356 38635 66358
rect 38362 66326 38388 66356
rect 38588 66326 38635 66356
rect 38619 66324 38635 66326
rect 38669 66324 38685 66358
rect 38619 66308 38685 66324
rect 38619 66048 38685 66064
rect 38619 66046 38635 66048
rect 38362 66016 38388 66046
rect 38588 66016 38635 66046
rect 38619 66014 38635 66016
rect 38669 66014 38685 66048
rect 38619 65998 38685 66014
rect 42792 66358 42858 66374
rect 42792 66324 42808 66358
rect 42842 66356 42858 66358
rect 42842 66326 42880 66356
rect 43080 66326 43106 66356
rect 42842 66324 42858 66326
rect 42792 66308 42858 66324
rect 42792 66048 42858 66064
rect 42792 66014 42808 66048
rect 42842 66046 42858 66048
rect 42842 66016 42880 66046
rect 43080 66016 43106 66046
rect 42842 66014 42858 66016
rect 42792 65998 42858 66014
rect 43609 66358 43675 66374
rect 43609 66356 43625 66358
rect 43352 66326 43378 66356
rect 43578 66326 43625 66356
rect 43609 66324 43625 66326
rect 43659 66324 43675 66358
rect 43609 66308 43675 66324
rect 43609 66048 43675 66064
rect 43609 66046 43625 66048
rect 43352 66016 43378 66046
rect 43578 66016 43625 66046
rect 43609 66014 43625 66016
rect 43659 66014 43675 66048
rect 43609 65998 43675 66014
rect 47782 66358 47848 66374
rect 47782 66324 47798 66358
rect 47832 66356 47848 66358
rect 47832 66326 47870 66356
rect 48070 66326 48096 66356
rect 47832 66324 47848 66326
rect 47782 66308 47848 66324
rect 47782 66048 47848 66064
rect 47782 66014 47798 66048
rect 47832 66046 47848 66048
rect 47832 66016 47870 66046
rect 48070 66016 48096 66046
rect 47832 66014 47848 66016
rect 47782 65998 47848 66014
rect 48599 66358 48665 66374
rect 48599 66356 48615 66358
rect 48342 66326 48368 66356
rect 48568 66326 48615 66356
rect 48599 66324 48615 66326
rect 48649 66324 48665 66358
rect 48599 66308 48665 66324
rect 48599 66048 48665 66064
rect 48599 66046 48615 66048
rect 48342 66016 48368 66046
rect 48568 66016 48615 66046
rect 48599 66014 48615 66016
rect 48649 66014 48665 66048
rect 48599 65998 48665 66014
rect 52772 66358 52838 66374
rect 52772 66324 52788 66358
rect 52822 66356 52838 66358
rect 52822 66326 52860 66356
rect 53060 66326 53086 66356
rect 52822 66324 52838 66326
rect 52772 66308 52838 66324
rect 52772 66048 52838 66064
rect 52772 66014 52788 66048
rect 52822 66046 52838 66048
rect 52822 66016 52860 66046
rect 53060 66016 53086 66046
rect 52822 66014 52838 66016
rect 52772 65998 52838 66014
rect 53589 66358 53655 66374
rect 53589 66356 53605 66358
rect 53332 66326 53358 66356
rect 53558 66326 53605 66356
rect 53589 66324 53605 66326
rect 53639 66324 53655 66358
rect 53589 66308 53655 66324
rect 53589 66048 53655 66064
rect 53589 66046 53605 66048
rect 53332 66016 53358 66046
rect 53558 66016 53605 66046
rect 53589 66014 53605 66016
rect 53639 66014 53655 66048
rect 53589 65998 53655 66014
rect 57762 66358 57828 66374
rect 57762 66324 57778 66358
rect 57812 66356 57828 66358
rect 57812 66326 57850 66356
rect 58050 66326 58076 66356
rect 57812 66324 57828 66326
rect 57762 66308 57828 66324
rect 57762 66048 57828 66064
rect 57762 66014 57778 66048
rect 57812 66046 57828 66048
rect 57812 66016 57850 66046
rect 58050 66016 58076 66046
rect 57812 66014 57828 66016
rect 57762 65998 57828 66014
rect 58579 66358 58645 66374
rect 58579 66356 58595 66358
rect 58322 66326 58348 66356
rect 58548 66326 58595 66356
rect 58579 66324 58595 66326
rect 58629 66324 58645 66358
rect 58579 66308 58645 66324
rect 58579 66048 58645 66064
rect 58579 66046 58595 66048
rect 58322 66016 58348 66046
rect 58548 66016 58595 66046
rect 58579 66014 58595 66016
rect 58629 66014 58645 66048
rect 58579 65998 58645 66014
rect 62752 66358 62818 66374
rect 62752 66324 62768 66358
rect 62802 66356 62818 66358
rect 62802 66326 62840 66356
rect 63040 66326 63066 66356
rect 62802 66324 62818 66326
rect 62752 66308 62818 66324
rect 62752 66048 62818 66064
rect 62752 66014 62768 66048
rect 62802 66046 62818 66048
rect 62802 66016 62840 66046
rect 63040 66016 63066 66046
rect 62802 66014 62818 66016
rect 62752 65998 62818 66014
rect 63569 66358 63635 66374
rect 63569 66356 63585 66358
rect 63312 66326 63338 66356
rect 63538 66326 63585 66356
rect 63569 66324 63585 66326
rect 63619 66324 63635 66358
rect 63569 66308 63635 66324
rect 63569 66048 63635 66064
rect 63569 66046 63585 66048
rect 63312 66016 63338 66046
rect 63538 66016 63585 66046
rect 63569 66014 63585 66016
rect 63619 66014 63635 66048
rect 63569 65998 63635 66014
rect 67742 66358 67808 66374
rect 67742 66324 67758 66358
rect 67792 66356 67808 66358
rect 67792 66326 67830 66356
rect 68030 66326 68056 66356
rect 67792 66324 67808 66326
rect 67742 66308 67808 66324
rect 67742 66048 67808 66064
rect 67742 66014 67758 66048
rect 67792 66046 67808 66048
rect 67792 66016 67830 66046
rect 68030 66016 68056 66046
rect 67792 66014 67808 66016
rect 67742 65998 67808 66014
rect 68559 66358 68625 66374
rect 68559 66356 68575 66358
rect 68302 66326 68328 66356
rect 68528 66326 68575 66356
rect 68559 66324 68575 66326
rect 68609 66324 68625 66358
rect 68559 66308 68625 66324
rect 68559 66048 68625 66064
rect 68559 66046 68575 66048
rect 68302 66016 68328 66046
rect 68528 66016 68575 66046
rect 68559 66014 68575 66016
rect 68609 66014 68625 66048
rect 68559 65998 68625 66014
rect 72732 66358 72798 66374
rect 72732 66324 72748 66358
rect 72782 66356 72798 66358
rect 72782 66326 72820 66356
rect 73020 66326 73046 66356
rect 72782 66324 72798 66326
rect 72732 66308 72798 66324
rect 72732 66048 72798 66064
rect 72732 66014 72748 66048
rect 72782 66046 72798 66048
rect 72782 66016 72820 66046
rect 73020 66016 73046 66046
rect 72782 66014 72798 66016
rect 72732 65998 72798 66014
rect 73549 66358 73615 66374
rect 73549 66356 73565 66358
rect 73292 66326 73318 66356
rect 73518 66326 73565 66356
rect 73549 66324 73565 66326
rect 73599 66324 73615 66358
rect 73549 66308 73615 66324
rect 73549 66048 73615 66064
rect 73549 66046 73565 66048
rect 73292 66016 73318 66046
rect 73518 66016 73565 66046
rect 73549 66014 73565 66016
rect 73599 66014 73615 66048
rect 73549 65998 73615 66014
rect 77722 66358 77788 66374
rect 77722 66324 77738 66358
rect 77772 66356 77788 66358
rect 77772 66326 77810 66356
rect 78010 66326 78036 66356
rect 77772 66324 77788 66326
rect 77722 66308 77788 66324
rect 77722 66048 77788 66064
rect 77722 66014 77738 66048
rect 77772 66046 77788 66048
rect 77772 66016 77810 66046
rect 78010 66016 78036 66046
rect 77772 66014 77788 66016
rect 77722 65998 77788 66014
rect 78539 66358 78605 66374
rect 78539 66356 78555 66358
rect 78282 66326 78308 66356
rect 78508 66326 78555 66356
rect 78539 66324 78555 66326
rect 78589 66324 78605 66358
rect 78539 66308 78605 66324
rect 78539 66048 78605 66064
rect 78539 66046 78555 66048
rect 78282 66016 78308 66046
rect 78508 66016 78555 66046
rect 78539 66014 78555 66016
rect 78589 66014 78605 66048
rect 78539 65998 78605 66014
rect 2872 64648 2938 64664
rect 2872 64614 2888 64648
rect 2922 64646 2938 64648
rect 2922 64616 2960 64646
rect 3160 64616 3186 64646
rect 2922 64614 2938 64616
rect 2872 64598 2938 64614
rect 2872 64338 2938 64354
rect 2872 64304 2888 64338
rect 2922 64336 2938 64338
rect 2922 64306 2960 64336
rect 3160 64306 3186 64336
rect 2922 64304 2938 64306
rect 2872 64288 2938 64304
rect 3689 64648 3755 64664
rect 3689 64646 3705 64648
rect 3432 64616 3458 64646
rect 3658 64616 3705 64646
rect 3689 64614 3705 64616
rect 3739 64614 3755 64648
rect 3689 64598 3755 64614
rect 3689 64338 3755 64354
rect 3689 64336 3705 64338
rect 3432 64306 3458 64336
rect 3658 64306 3705 64336
rect 3689 64304 3705 64306
rect 3739 64304 3755 64338
rect 3689 64288 3755 64304
rect 7862 64648 7928 64664
rect 7862 64614 7878 64648
rect 7912 64646 7928 64648
rect 7912 64616 7950 64646
rect 8150 64616 8176 64646
rect 7912 64614 7928 64616
rect 7862 64598 7928 64614
rect 7862 64338 7928 64354
rect 7862 64304 7878 64338
rect 7912 64336 7928 64338
rect 7912 64306 7950 64336
rect 8150 64306 8176 64336
rect 7912 64304 7928 64306
rect 7862 64288 7928 64304
rect 8679 64648 8745 64664
rect 8679 64646 8695 64648
rect 8422 64616 8448 64646
rect 8648 64616 8695 64646
rect 8679 64614 8695 64616
rect 8729 64614 8745 64648
rect 8679 64598 8745 64614
rect 8679 64338 8745 64354
rect 8679 64336 8695 64338
rect 8422 64306 8448 64336
rect 8648 64306 8695 64336
rect 8679 64304 8695 64306
rect 8729 64304 8745 64338
rect 8679 64288 8745 64304
rect 12852 64648 12918 64664
rect 12852 64614 12868 64648
rect 12902 64646 12918 64648
rect 12902 64616 12940 64646
rect 13140 64616 13166 64646
rect 12902 64614 12918 64616
rect 12852 64598 12918 64614
rect 12852 64338 12918 64354
rect 12852 64304 12868 64338
rect 12902 64336 12918 64338
rect 12902 64306 12940 64336
rect 13140 64306 13166 64336
rect 12902 64304 12918 64306
rect 12852 64288 12918 64304
rect 13669 64648 13735 64664
rect 13669 64646 13685 64648
rect 13412 64616 13438 64646
rect 13638 64616 13685 64646
rect 13669 64614 13685 64616
rect 13719 64614 13735 64648
rect 13669 64598 13735 64614
rect 13669 64338 13735 64354
rect 13669 64336 13685 64338
rect 13412 64306 13438 64336
rect 13638 64306 13685 64336
rect 13669 64304 13685 64306
rect 13719 64304 13735 64338
rect 13669 64288 13735 64304
rect 17842 64648 17908 64664
rect 17842 64614 17858 64648
rect 17892 64646 17908 64648
rect 17892 64616 17930 64646
rect 18130 64616 18156 64646
rect 17892 64614 17908 64616
rect 17842 64598 17908 64614
rect 17842 64338 17908 64354
rect 17842 64304 17858 64338
rect 17892 64336 17908 64338
rect 17892 64306 17930 64336
rect 18130 64306 18156 64336
rect 17892 64304 17908 64306
rect 17842 64288 17908 64304
rect 18659 64648 18725 64664
rect 18659 64646 18675 64648
rect 18402 64616 18428 64646
rect 18628 64616 18675 64646
rect 18659 64614 18675 64616
rect 18709 64614 18725 64648
rect 18659 64598 18725 64614
rect 18659 64338 18725 64354
rect 18659 64336 18675 64338
rect 18402 64306 18428 64336
rect 18628 64306 18675 64336
rect 18659 64304 18675 64306
rect 18709 64304 18725 64338
rect 18659 64288 18725 64304
rect 22832 64648 22898 64664
rect 22832 64614 22848 64648
rect 22882 64646 22898 64648
rect 22882 64616 22920 64646
rect 23120 64616 23146 64646
rect 22882 64614 22898 64616
rect 22832 64598 22898 64614
rect 22832 64338 22898 64354
rect 22832 64304 22848 64338
rect 22882 64336 22898 64338
rect 22882 64306 22920 64336
rect 23120 64306 23146 64336
rect 22882 64304 22898 64306
rect 22832 64288 22898 64304
rect 23649 64648 23715 64664
rect 23649 64646 23665 64648
rect 23392 64616 23418 64646
rect 23618 64616 23665 64646
rect 23649 64614 23665 64616
rect 23699 64614 23715 64648
rect 23649 64598 23715 64614
rect 23649 64338 23715 64354
rect 23649 64336 23665 64338
rect 23392 64306 23418 64336
rect 23618 64306 23665 64336
rect 23649 64304 23665 64306
rect 23699 64304 23715 64338
rect 23649 64288 23715 64304
rect 27822 64648 27888 64664
rect 27822 64614 27838 64648
rect 27872 64646 27888 64648
rect 27872 64616 27910 64646
rect 28110 64616 28136 64646
rect 27872 64614 27888 64616
rect 27822 64598 27888 64614
rect 27822 64338 27888 64354
rect 27822 64304 27838 64338
rect 27872 64336 27888 64338
rect 27872 64306 27910 64336
rect 28110 64306 28136 64336
rect 27872 64304 27888 64306
rect 27822 64288 27888 64304
rect 28639 64648 28705 64664
rect 28639 64646 28655 64648
rect 28382 64616 28408 64646
rect 28608 64616 28655 64646
rect 28639 64614 28655 64616
rect 28689 64614 28705 64648
rect 28639 64598 28705 64614
rect 28639 64338 28705 64354
rect 28639 64336 28655 64338
rect 28382 64306 28408 64336
rect 28608 64306 28655 64336
rect 28639 64304 28655 64306
rect 28689 64304 28705 64338
rect 28639 64288 28705 64304
rect 32812 64648 32878 64664
rect 32812 64614 32828 64648
rect 32862 64646 32878 64648
rect 32862 64616 32900 64646
rect 33100 64616 33126 64646
rect 32862 64614 32878 64616
rect 32812 64598 32878 64614
rect 32812 64338 32878 64354
rect 32812 64304 32828 64338
rect 32862 64336 32878 64338
rect 32862 64306 32900 64336
rect 33100 64306 33126 64336
rect 32862 64304 32878 64306
rect 32812 64288 32878 64304
rect 33629 64648 33695 64664
rect 33629 64646 33645 64648
rect 33372 64616 33398 64646
rect 33598 64616 33645 64646
rect 33629 64614 33645 64616
rect 33679 64614 33695 64648
rect 33629 64598 33695 64614
rect 33629 64338 33695 64354
rect 33629 64336 33645 64338
rect 33372 64306 33398 64336
rect 33598 64306 33645 64336
rect 33629 64304 33645 64306
rect 33679 64304 33695 64338
rect 33629 64288 33695 64304
rect 37802 64648 37868 64664
rect 37802 64614 37818 64648
rect 37852 64646 37868 64648
rect 37852 64616 37890 64646
rect 38090 64616 38116 64646
rect 37852 64614 37868 64616
rect 37802 64598 37868 64614
rect 37802 64338 37868 64354
rect 37802 64304 37818 64338
rect 37852 64336 37868 64338
rect 37852 64306 37890 64336
rect 38090 64306 38116 64336
rect 37852 64304 37868 64306
rect 37802 64288 37868 64304
rect 38619 64648 38685 64664
rect 38619 64646 38635 64648
rect 38362 64616 38388 64646
rect 38588 64616 38635 64646
rect 38619 64614 38635 64616
rect 38669 64614 38685 64648
rect 38619 64598 38685 64614
rect 38619 64338 38685 64354
rect 38619 64336 38635 64338
rect 38362 64306 38388 64336
rect 38588 64306 38635 64336
rect 38619 64304 38635 64306
rect 38669 64304 38685 64338
rect 38619 64288 38685 64304
rect 42792 64648 42858 64664
rect 42792 64614 42808 64648
rect 42842 64646 42858 64648
rect 42842 64616 42880 64646
rect 43080 64616 43106 64646
rect 42842 64614 42858 64616
rect 42792 64598 42858 64614
rect 42792 64338 42858 64354
rect 42792 64304 42808 64338
rect 42842 64336 42858 64338
rect 42842 64306 42880 64336
rect 43080 64306 43106 64336
rect 42842 64304 42858 64306
rect 42792 64288 42858 64304
rect 43609 64648 43675 64664
rect 43609 64646 43625 64648
rect 43352 64616 43378 64646
rect 43578 64616 43625 64646
rect 43609 64614 43625 64616
rect 43659 64614 43675 64648
rect 43609 64598 43675 64614
rect 43609 64338 43675 64354
rect 43609 64336 43625 64338
rect 43352 64306 43378 64336
rect 43578 64306 43625 64336
rect 43609 64304 43625 64306
rect 43659 64304 43675 64338
rect 43609 64288 43675 64304
rect 47782 64648 47848 64664
rect 47782 64614 47798 64648
rect 47832 64646 47848 64648
rect 47832 64616 47870 64646
rect 48070 64616 48096 64646
rect 47832 64614 47848 64616
rect 47782 64598 47848 64614
rect 47782 64338 47848 64354
rect 47782 64304 47798 64338
rect 47832 64336 47848 64338
rect 47832 64306 47870 64336
rect 48070 64306 48096 64336
rect 47832 64304 47848 64306
rect 47782 64288 47848 64304
rect 48599 64648 48665 64664
rect 48599 64646 48615 64648
rect 48342 64616 48368 64646
rect 48568 64616 48615 64646
rect 48599 64614 48615 64616
rect 48649 64614 48665 64648
rect 48599 64598 48665 64614
rect 48599 64338 48665 64354
rect 48599 64336 48615 64338
rect 48342 64306 48368 64336
rect 48568 64306 48615 64336
rect 48599 64304 48615 64306
rect 48649 64304 48665 64338
rect 48599 64288 48665 64304
rect 52772 64648 52838 64664
rect 52772 64614 52788 64648
rect 52822 64646 52838 64648
rect 52822 64616 52860 64646
rect 53060 64616 53086 64646
rect 52822 64614 52838 64616
rect 52772 64598 52838 64614
rect 52772 64338 52838 64354
rect 52772 64304 52788 64338
rect 52822 64336 52838 64338
rect 52822 64306 52860 64336
rect 53060 64306 53086 64336
rect 52822 64304 52838 64306
rect 52772 64288 52838 64304
rect 53589 64648 53655 64664
rect 53589 64646 53605 64648
rect 53332 64616 53358 64646
rect 53558 64616 53605 64646
rect 53589 64614 53605 64616
rect 53639 64614 53655 64648
rect 53589 64598 53655 64614
rect 53589 64338 53655 64354
rect 53589 64336 53605 64338
rect 53332 64306 53358 64336
rect 53558 64306 53605 64336
rect 53589 64304 53605 64306
rect 53639 64304 53655 64338
rect 53589 64288 53655 64304
rect 57762 64648 57828 64664
rect 57762 64614 57778 64648
rect 57812 64646 57828 64648
rect 57812 64616 57850 64646
rect 58050 64616 58076 64646
rect 57812 64614 57828 64616
rect 57762 64598 57828 64614
rect 57762 64338 57828 64354
rect 57762 64304 57778 64338
rect 57812 64336 57828 64338
rect 57812 64306 57850 64336
rect 58050 64306 58076 64336
rect 57812 64304 57828 64306
rect 57762 64288 57828 64304
rect 58579 64648 58645 64664
rect 58579 64646 58595 64648
rect 58322 64616 58348 64646
rect 58548 64616 58595 64646
rect 58579 64614 58595 64616
rect 58629 64614 58645 64648
rect 58579 64598 58645 64614
rect 58579 64338 58645 64354
rect 58579 64336 58595 64338
rect 58322 64306 58348 64336
rect 58548 64306 58595 64336
rect 58579 64304 58595 64306
rect 58629 64304 58645 64338
rect 58579 64288 58645 64304
rect 62752 64648 62818 64664
rect 62752 64614 62768 64648
rect 62802 64646 62818 64648
rect 62802 64616 62840 64646
rect 63040 64616 63066 64646
rect 62802 64614 62818 64616
rect 62752 64598 62818 64614
rect 62752 64338 62818 64354
rect 62752 64304 62768 64338
rect 62802 64336 62818 64338
rect 62802 64306 62840 64336
rect 63040 64306 63066 64336
rect 62802 64304 62818 64306
rect 62752 64288 62818 64304
rect 63569 64648 63635 64664
rect 63569 64646 63585 64648
rect 63312 64616 63338 64646
rect 63538 64616 63585 64646
rect 63569 64614 63585 64616
rect 63619 64614 63635 64648
rect 63569 64598 63635 64614
rect 63569 64338 63635 64354
rect 63569 64336 63585 64338
rect 63312 64306 63338 64336
rect 63538 64306 63585 64336
rect 63569 64304 63585 64306
rect 63619 64304 63635 64338
rect 63569 64288 63635 64304
rect 67742 64648 67808 64664
rect 67742 64614 67758 64648
rect 67792 64646 67808 64648
rect 67792 64616 67830 64646
rect 68030 64616 68056 64646
rect 67792 64614 67808 64616
rect 67742 64598 67808 64614
rect 67742 64338 67808 64354
rect 67742 64304 67758 64338
rect 67792 64336 67808 64338
rect 67792 64306 67830 64336
rect 68030 64306 68056 64336
rect 67792 64304 67808 64306
rect 67742 64288 67808 64304
rect 68559 64648 68625 64664
rect 68559 64646 68575 64648
rect 68302 64616 68328 64646
rect 68528 64616 68575 64646
rect 68559 64614 68575 64616
rect 68609 64614 68625 64648
rect 68559 64598 68625 64614
rect 68559 64338 68625 64354
rect 68559 64336 68575 64338
rect 68302 64306 68328 64336
rect 68528 64306 68575 64336
rect 68559 64304 68575 64306
rect 68609 64304 68625 64338
rect 68559 64288 68625 64304
rect 72732 64648 72798 64664
rect 72732 64614 72748 64648
rect 72782 64646 72798 64648
rect 72782 64616 72820 64646
rect 73020 64616 73046 64646
rect 72782 64614 72798 64616
rect 72732 64598 72798 64614
rect 72732 64338 72798 64354
rect 72732 64304 72748 64338
rect 72782 64336 72798 64338
rect 72782 64306 72820 64336
rect 73020 64306 73046 64336
rect 72782 64304 72798 64306
rect 72732 64288 72798 64304
rect 73549 64648 73615 64664
rect 73549 64646 73565 64648
rect 73292 64616 73318 64646
rect 73518 64616 73565 64646
rect 73549 64614 73565 64616
rect 73599 64614 73615 64648
rect 73549 64598 73615 64614
rect 73549 64338 73615 64354
rect 73549 64336 73565 64338
rect 73292 64306 73318 64336
rect 73518 64306 73565 64336
rect 73549 64304 73565 64306
rect 73599 64304 73615 64338
rect 73549 64288 73615 64304
rect 77722 64648 77788 64664
rect 77722 64614 77738 64648
rect 77772 64646 77788 64648
rect 77772 64616 77810 64646
rect 78010 64616 78036 64646
rect 77772 64614 77788 64616
rect 77722 64598 77788 64614
rect 77722 64338 77788 64354
rect 77722 64304 77738 64338
rect 77772 64336 77788 64338
rect 77772 64306 77810 64336
rect 78010 64306 78036 64336
rect 77772 64304 77788 64306
rect 77722 64288 77788 64304
rect 78539 64648 78605 64664
rect 78539 64646 78555 64648
rect 78282 64616 78308 64646
rect 78508 64616 78555 64646
rect 78539 64614 78555 64616
rect 78589 64614 78605 64648
rect 78539 64598 78605 64614
rect 78539 64338 78605 64354
rect 78539 64336 78555 64338
rect 78282 64306 78308 64336
rect 78508 64306 78555 64336
rect 78539 64304 78555 64306
rect 78589 64304 78605 64338
rect 78539 64288 78605 64304
rect 2872 62938 2938 62954
rect 2872 62904 2888 62938
rect 2922 62936 2938 62938
rect 2922 62906 2960 62936
rect 3160 62906 3186 62936
rect 2922 62904 2938 62906
rect 2872 62888 2938 62904
rect 2872 62628 2938 62644
rect 2872 62594 2888 62628
rect 2922 62626 2938 62628
rect 2922 62596 2960 62626
rect 3160 62596 3186 62626
rect 2922 62594 2938 62596
rect 2872 62578 2938 62594
rect 3689 62938 3755 62954
rect 3689 62936 3705 62938
rect 3432 62906 3458 62936
rect 3658 62906 3705 62936
rect 3689 62904 3705 62906
rect 3739 62904 3755 62938
rect 3689 62888 3755 62904
rect 3689 62628 3755 62644
rect 3689 62626 3705 62628
rect 3432 62596 3458 62626
rect 3658 62596 3705 62626
rect 3689 62594 3705 62596
rect 3739 62594 3755 62628
rect 3689 62578 3755 62594
rect 7862 62938 7928 62954
rect 7862 62904 7878 62938
rect 7912 62936 7928 62938
rect 7912 62906 7950 62936
rect 8150 62906 8176 62936
rect 7912 62904 7928 62906
rect 7862 62888 7928 62904
rect 7862 62628 7928 62644
rect 7862 62594 7878 62628
rect 7912 62626 7928 62628
rect 7912 62596 7950 62626
rect 8150 62596 8176 62626
rect 7912 62594 7928 62596
rect 7862 62578 7928 62594
rect 8679 62938 8745 62954
rect 8679 62936 8695 62938
rect 8422 62906 8448 62936
rect 8648 62906 8695 62936
rect 8679 62904 8695 62906
rect 8729 62904 8745 62938
rect 8679 62888 8745 62904
rect 8679 62628 8745 62644
rect 8679 62626 8695 62628
rect 8422 62596 8448 62626
rect 8648 62596 8695 62626
rect 8679 62594 8695 62596
rect 8729 62594 8745 62628
rect 8679 62578 8745 62594
rect 12852 62938 12918 62954
rect 12852 62904 12868 62938
rect 12902 62936 12918 62938
rect 12902 62906 12940 62936
rect 13140 62906 13166 62936
rect 12902 62904 12918 62906
rect 12852 62888 12918 62904
rect 12852 62628 12918 62644
rect 12852 62594 12868 62628
rect 12902 62626 12918 62628
rect 12902 62596 12940 62626
rect 13140 62596 13166 62626
rect 12902 62594 12918 62596
rect 12852 62578 12918 62594
rect 13669 62938 13735 62954
rect 13669 62936 13685 62938
rect 13412 62906 13438 62936
rect 13638 62906 13685 62936
rect 13669 62904 13685 62906
rect 13719 62904 13735 62938
rect 13669 62888 13735 62904
rect 13669 62628 13735 62644
rect 13669 62626 13685 62628
rect 13412 62596 13438 62626
rect 13638 62596 13685 62626
rect 13669 62594 13685 62596
rect 13719 62594 13735 62628
rect 13669 62578 13735 62594
rect 17842 62938 17908 62954
rect 17842 62904 17858 62938
rect 17892 62936 17908 62938
rect 17892 62906 17930 62936
rect 18130 62906 18156 62936
rect 17892 62904 17908 62906
rect 17842 62888 17908 62904
rect 17842 62628 17908 62644
rect 17842 62594 17858 62628
rect 17892 62626 17908 62628
rect 17892 62596 17930 62626
rect 18130 62596 18156 62626
rect 17892 62594 17908 62596
rect 17842 62578 17908 62594
rect 18659 62938 18725 62954
rect 18659 62936 18675 62938
rect 18402 62906 18428 62936
rect 18628 62906 18675 62936
rect 18659 62904 18675 62906
rect 18709 62904 18725 62938
rect 18659 62888 18725 62904
rect 18659 62628 18725 62644
rect 18659 62626 18675 62628
rect 18402 62596 18428 62626
rect 18628 62596 18675 62626
rect 18659 62594 18675 62596
rect 18709 62594 18725 62628
rect 18659 62578 18725 62594
rect 22832 62938 22898 62954
rect 22832 62904 22848 62938
rect 22882 62936 22898 62938
rect 22882 62906 22920 62936
rect 23120 62906 23146 62936
rect 22882 62904 22898 62906
rect 22832 62888 22898 62904
rect 22832 62628 22898 62644
rect 22832 62594 22848 62628
rect 22882 62626 22898 62628
rect 22882 62596 22920 62626
rect 23120 62596 23146 62626
rect 22882 62594 22898 62596
rect 22832 62578 22898 62594
rect 23649 62938 23715 62954
rect 23649 62936 23665 62938
rect 23392 62906 23418 62936
rect 23618 62906 23665 62936
rect 23649 62904 23665 62906
rect 23699 62904 23715 62938
rect 23649 62888 23715 62904
rect 23649 62628 23715 62644
rect 23649 62626 23665 62628
rect 23392 62596 23418 62626
rect 23618 62596 23665 62626
rect 23649 62594 23665 62596
rect 23699 62594 23715 62628
rect 23649 62578 23715 62594
rect 27822 62938 27888 62954
rect 27822 62904 27838 62938
rect 27872 62936 27888 62938
rect 27872 62906 27910 62936
rect 28110 62906 28136 62936
rect 27872 62904 27888 62906
rect 27822 62888 27888 62904
rect 27822 62628 27888 62644
rect 27822 62594 27838 62628
rect 27872 62626 27888 62628
rect 27872 62596 27910 62626
rect 28110 62596 28136 62626
rect 27872 62594 27888 62596
rect 27822 62578 27888 62594
rect 28639 62938 28705 62954
rect 28639 62936 28655 62938
rect 28382 62906 28408 62936
rect 28608 62906 28655 62936
rect 28639 62904 28655 62906
rect 28689 62904 28705 62938
rect 28639 62888 28705 62904
rect 28639 62628 28705 62644
rect 28639 62626 28655 62628
rect 28382 62596 28408 62626
rect 28608 62596 28655 62626
rect 28639 62594 28655 62596
rect 28689 62594 28705 62628
rect 28639 62578 28705 62594
rect 32812 62938 32878 62954
rect 32812 62904 32828 62938
rect 32862 62936 32878 62938
rect 32862 62906 32900 62936
rect 33100 62906 33126 62936
rect 32862 62904 32878 62906
rect 32812 62888 32878 62904
rect 32812 62628 32878 62644
rect 32812 62594 32828 62628
rect 32862 62626 32878 62628
rect 32862 62596 32900 62626
rect 33100 62596 33126 62626
rect 32862 62594 32878 62596
rect 32812 62578 32878 62594
rect 33629 62938 33695 62954
rect 33629 62936 33645 62938
rect 33372 62906 33398 62936
rect 33598 62906 33645 62936
rect 33629 62904 33645 62906
rect 33679 62904 33695 62938
rect 33629 62888 33695 62904
rect 33629 62628 33695 62644
rect 33629 62626 33645 62628
rect 33372 62596 33398 62626
rect 33598 62596 33645 62626
rect 33629 62594 33645 62596
rect 33679 62594 33695 62628
rect 33629 62578 33695 62594
rect 37802 62938 37868 62954
rect 37802 62904 37818 62938
rect 37852 62936 37868 62938
rect 37852 62906 37890 62936
rect 38090 62906 38116 62936
rect 37852 62904 37868 62906
rect 37802 62888 37868 62904
rect 37802 62628 37868 62644
rect 37802 62594 37818 62628
rect 37852 62626 37868 62628
rect 37852 62596 37890 62626
rect 38090 62596 38116 62626
rect 37852 62594 37868 62596
rect 37802 62578 37868 62594
rect 38619 62938 38685 62954
rect 38619 62936 38635 62938
rect 38362 62906 38388 62936
rect 38588 62906 38635 62936
rect 38619 62904 38635 62906
rect 38669 62904 38685 62938
rect 38619 62888 38685 62904
rect 38619 62628 38685 62644
rect 38619 62626 38635 62628
rect 38362 62596 38388 62626
rect 38588 62596 38635 62626
rect 38619 62594 38635 62596
rect 38669 62594 38685 62628
rect 38619 62578 38685 62594
rect 42792 62938 42858 62954
rect 42792 62904 42808 62938
rect 42842 62936 42858 62938
rect 42842 62906 42880 62936
rect 43080 62906 43106 62936
rect 42842 62904 42858 62906
rect 42792 62888 42858 62904
rect 42792 62628 42858 62644
rect 42792 62594 42808 62628
rect 42842 62626 42858 62628
rect 42842 62596 42880 62626
rect 43080 62596 43106 62626
rect 42842 62594 42858 62596
rect 42792 62578 42858 62594
rect 43609 62938 43675 62954
rect 43609 62936 43625 62938
rect 43352 62906 43378 62936
rect 43578 62906 43625 62936
rect 43609 62904 43625 62906
rect 43659 62904 43675 62938
rect 43609 62888 43675 62904
rect 43609 62628 43675 62644
rect 43609 62626 43625 62628
rect 43352 62596 43378 62626
rect 43578 62596 43625 62626
rect 43609 62594 43625 62596
rect 43659 62594 43675 62628
rect 43609 62578 43675 62594
rect 47782 62938 47848 62954
rect 47782 62904 47798 62938
rect 47832 62936 47848 62938
rect 47832 62906 47870 62936
rect 48070 62906 48096 62936
rect 47832 62904 47848 62906
rect 47782 62888 47848 62904
rect 47782 62628 47848 62644
rect 47782 62594 47798 62628
rect 47832 62626 47848 62628
rect 47832 62596 47870 62626
rect 48070 62596 48096 62626
rect 47832 62594 47848 62596
rect 47782 62578 47848 62594
rect 48599 62938 48665 62954
rect 48599 62936 48615 62938
rect 48342 62906 48368 62936
rect 48568 62906 48615 62936
rect 48599 62904 48615 62906
rect 48649 62904 48665 62938
rect 48599 62888 48665 62904
rect 48599 62628 48665 62644
rect 48599 62626 48615 62628
rect 48342 62596 48368 62626
rect 48568 62596 48615 62626
rect 48599 62594 48615 62596
rect 48649 62594 48665 62628
rect 48599 62578 48665 62594
rect 52772 62938 52838 62954
rect 52772 62904 52788 62938
rect 52822 62936 52838 62938
rect 52822 62906 52860 62936
rect 53060 62906 53086 62936
rect 52822 62904 52838 62906
rect 52772 62888 52838 62904
rect 52772 62628 52838 62644
rect 52772 62594 52788 62628
rect 52822 62626 52838 62628
rect 52822 62596 52860 62626
rect 53060 62596 53086 62626
rect 52822 62594 52838 62596
rect 52772 62578 52838 62594
rect 53589 62938 53655 62954
rect 53589 62936 53605 62938
rect 53332 62906 53358 62936
rect 53558 62906 53605 62936
rect 53589 62904 53605 62906
rect 53639 62904 53655 62938
rect 53589 62888 53655 62904
rect 53589 62628 53655 62644
rect 53589 62626 53605 62628
rect 53332 62596 53358 62626
rect 53558 62596 53605 62626
rect 53589 62594 53605 62596
rect 53639 62594 53655 62628
rect 53589 62578 53655 62594
rect 57762 62938 57828 62954
rect 57762 62904 57778 62938
rect 57812 62936 57828 62938
rect 57812 62906 57850 62936
rect 58050 62906 58076 62936
rect 57812 62904 57828 62906
rect 57762 62888 57828 62904
rect 57762 62628 57828 62644
rect 57762 62594 57778 62628
rect 57812 62626 57828 62628
rect 57812 62596 57850 62626
rect 58050 62596 58076 62626
rect 57812 62594 57828 62596
rect 57762 62578 57828 62594
rect 58579 62938 58645 62954
rect 58579 62936 58595 62938
rect 58322 62906 58348 62936
rect 58548 62906 58595 62936
rect 58579 62904 58595 62906
rect 58629 62904 58645 62938
rect 58579 62888 58645 62904
rect 58579 62628 58645 62644
rect 58579 62626 58595 62628
rect 58322 62596 58348 62626
rect 58548 62596 58595 62626
rect 58579 62594 58595 62596
rect 58629 62594 58645 62628
rect 58579 62578 58645 62594
rect 62752 62938 62818 62954
rect 62752 62904 62768 62938
rect 62802 62936 62818 62938
rect 62802 62906 62840 62936
rect 63040 62906 63066 62936
rect 62802 62904 62818 62906
rect 62752 62888 62818 62904
rect 62752 62628 62818 62644
rect 62752 62594 62768 62628
rect 62802 62626 62818 62628
rect 62802 62596 62840 62626
rect 63040 62596 63066 62626
rect 62802 62594 62818 62596
rect 62752 62578 62818 62594
rect 63569 62938 63635 62954
rect 63569 62936 63585 62938
rect 63312 62906 63338 62936
rect 63538 62906 63585 62936
rect 63569 62904 63585 62906
rect 63619 62904 63635 62938
rect 63569 62888 63635 62904
rect 63569 62628 63635 62644
rect 63569 62626 63585 62628
rect 63312 62596 63338 62626
rect 63538 62596 63585 62626
rect 63569 62594 63585 62596
rect 63619 62594 63635 62628
rect 63569 62578 63635 62594
rect 67742 62938 67808 62954
rect 67742 62904 67758 62938
rect 67792 62936 67808 62938
rect 67792 62906 67830 62936
rect 68030 62906 68056 62936
rect 67792 62904 67808 62906
rect 67742 62888 67808 62904
rect 67742 62628 67808 62644
rect 67742 62594 67758 62628
rect 67792 62626 67808 62628
rect 67792 62596 67830 62626
rect 68030 62596 68056 62626
rect 67792 62594 67808 62596
rect 67742 62578 67808 62594
rect 68559 62938 68625 62954
rect 68559 62936 68575 62938
rect 68302 62906 68328 62936
rect 68528 62906 68575 62936
rect 68559 62904 68575 62906
rect 68609 62904 68625 62938
rect 68559 62888 68625 62904
rect 68559 62628 68625 62644
rect 68559 62626 68575 62628
rect 68302 62596 68328 62626
rect 68528 62596 68575 62626
rect 68559 62594 68575 62596
rect 68609 62594 68625 62628
rect 68559 62578 68625 62594
rect 72732 62938 72798 62954
rect 72732 62904 72748 62938
rect 72782 62936 72798 62938
rect 72782 62906 72820 62936
rect 73020 62906 73046 62936
rect 72782 62904 72798 62906
rect 72732 62888 72798 62904
rect 72732 62628 72798 62644
rect 72732 62594 72748 62628
rect 72782 62626 72798 62628
rect 72782 62596 72820 62626
rect 73020 62596 73046 62626
rect 72782 62594 72798 62596
rect 72732 62578 72798 62594
rect 73549 62938 73615 62954
rect 73549 62936 73565 62938
rect 73292 62906 73318 62936
rect 73518 62906 73565 62936
rect 73549 62904 73565 62906
rect 73599 62904 73615 62938
rect 73549 62888 73615 62904
rect 73549 62628 73615 62644
rect 73549 62626 73565 62628
rect 73292 62596 73318 62626
rect 73518 62596 73565 62626
rect 73549 62594 73565 62596
rect 73599 62594 73615 62628
rect 73549 62578 73615 62594
rect 77722 62938 77788 62954
rect 77722 62904 77738 62938
rect 77772 62936 77788 62938
rect 77772 62906 77810 62936
rect 78010 62906 78036 62936
rect 77772 62904 77788 62906
rect 77722 62888 77788 62904
rect 77722 62628 77788 62644
rect 77722 62594 77738 62628
rect 77772 62626 77788 62628
rect 77772 62596 77810 62626
rect 78010 62596 78036 62626
rect 77772 62594 77788 62596
rect 77722 62578 77788 62594
rect 78539 62938 78605 62954
rect 78539 62936 78555 62938
rect 78282 62906 78308 62936
rect 78508 62906 78555 62936
rect 78539 62904 78555 62906
rect 78589 62904 78605 62938
rect 78539 62888 78605 62904
rect 78539 62628 78605 62644
rect 78539 62626 78555 62628
rect 78282 62596 78308 62626
rect 78508 62596 78555 62626
rect 78539 62594 78555 62596
rect 78589 62594 78605 62628
rect 78539 62578 78605 62594
rect 2872 61228 2938 61244
rect 2872 61194 2888 61228
rect 2922 61226 2938 61228
rect 2922 61196 2960 61226
rect 3160 61196 3186 61226
rect 2922 61194 2938 61196
rect 2872 61178 2938 61194
rect 2872 60918 2938 60934
rect 2872 60884 2888 60918
rect 2922 60916 2938 60918
rect 2922 60886 2960 60916
rect 3160 60886 3186 60916
rect 2922 60884 2938 60886
rect 2872 60868 2938 60884
rect 3689 61228 3755 61244
rect 3689 61226 3705 61228
rect 3432 61196 3458 61226
rect 3658 61196 3705 61226
rect 3689 61194 3705 61196
rect 3739 61194 3755 61228
rect 3689 61178 3755 61194
rect 3689 60918 3755 60934
rect 3689 60916 3705 60918
rect 3432 60886 3458 60916
rect 3658 60886 3705 60916
rect 3689 60884 3705 60886
rect 3739 60884 3755 60918
rect 3689 60868 3755 60884
rect 7862 61228 7928 61244
rect 7862 61194 7878 61228
rect 7912 61226 7928 61228
rect 7912 61196 7950 61226
rect 8150 61196 8176 61226
rect 7912 61194 7928 61196
rect 7862 61178 7928 61194
rect 7862 60918 7928 60934
rect 7862 60884 7878 60918
rect 7912 60916 7928 60918
rect 7912 60886 7950 60916
rect 8150 60886 8176 60916
rect 7912 60884 7928 60886
rect 7862 60868 7928 60884
rect 8679 61228 8745 61244
rect 8679 61226 8695 61228
rect 8422 61196 8448 61226
rect 8648 61196 8695 61226
rect 8679 61194 8695 61196
rect 8729 61194 8745 61228
rect 8679 61178 8745 61194
rect 8679 60918 8745 60934
rect 8679 60916 8695 60918
rect 8422 60886 8448 60916
rect 8648 60886 8695 60916
rect 8679 60884 8695 60886
rect 8729 60884 8745 60918
rect 8679 60868 8745 60884
rect 12852 61228 12918 61244
rect 12852 61194 12868 61228
rect 12902 61226 12918 61228
rect 12902 61196 12940 61226
rect 13140 61196 13166 61226
rect 12902 61194 12918 61196
rect 12852 61178 12918 61194
rect 12852 60918 12918 60934
rect 12852 60884 12868 60918
rect 12902 60916 12918 60918
rect 12902 60886 12940 60916
rect 13140 60886 13166 60916
rect 12902 60884 12918 60886
rect 12852 60868 12918 60884
rect 13669 61228 13735 61244
rect 13669 61226 13685 61228
rect 13412 61196 13438 61226
rect 13638 61196 13685 61226
rect 13669 61194 13685 61196
rect 13719 61194 13735 61228
rect 13669 61178 13735 61194
rect 13669 60918 13735 60934
rect 13669 60916 13685 60918
rect 13412 60886 13438 60916
rect 13638 60886 13685 60916
rect 13669 60884 13685 60886
rect 13719 60884 13735 60918
rect 13669 60868 13735 60884
rect 17842 61228 17908 61244
rect 17842 61194 17858 61228
rect 17892 61226 17908 61228
rect 17892 61196 17930 61226
rect 18130 61196 18156 61226
rect 17892 61194 17908 61196
rect 17842 61178 17908 61194
rect 17842 60918 17908 60934
rect 17842 60884 17858 60918
rect 17892 60916 17908 60918
rect 17892 60886 17930 60916
rect 18130 60886 18156 60916
rect 17892 60884 17908 60886
rect 17842 60868 17908 60884
rect 18659 61228 18725 61244
rect 18659 61226 18675 61228
rect 18402 61196 18428 61226
rect 18628 61196 18675 61226
rect 18659 61194 18675 61196
rect 18709 61194 18725 61228
rect 18659 61178 18725 61194
rect 18659 60918 18725 60934
rect 18659 60916 18675 60918
rect 18402 60886 18428 60916
rect 18628 60886 18675 60916
rect 18659 60884 18675 60886
rect 18709 60884 18725 60918
rect 18659 60868 18725 60884
rect 22832 61228 22898 61244
rect 22832 61194 22848 61228
rect 22882 61226 22898 61228
rect 22882 61196 22920 61226
rect 23120 61196 23146 61226
rect 22882 61194 22898 61196
rect 22832 61178 22898 61194
rect 22832 60918 22898 60934
rect 22832 60884 22848 60918
rect 22882 60916 22898 60918
rect 22882 60886 22920 60916
rect 23120 60886 23146 60916
rect 22882 60884 22898 60886
rect 22832 60868 22898 60884
rect 23649 61228 23715 61244
rect 23649 61226 23665 61228
rect 23392 61196 23418 61226
rect 23618 61196 23665 61226
rect 23649 61194 23665 61196
rect 23699 61194 23715 61228
rect 23649 61178 23715 61194
rect 23649 60918 23715 60934
rect 23649 60916 23665 60918
rect 23392 60886 23418 60916
rect 23618 60886 23665 60916
rect 23649 60884 23665 60886
rect 23699 60884 23715 60918
rect 23649 60868 23715 60884
rect 27822 61228 27888 61244
rect 27822 61194 27838 61228
rect 27872 61226 27888 61228
rect 27872 61196 27910 61226
rect 28110 61196 28136 61226
rect 27872 61194 27888 61196
rect 27822 61178 27888 61194
rect 27822 60918 27888 60934
rect 27822 60884 27838 60918
rect 27872 60916 27888 60918
rect 27872 60886 27910 60916
rect 28110 60886 28136 60916
rect 27872 60884 27888 60886
rect 27822 60868 27888 60884
rect 28639 61228 28705 61244
rect 28639 61226 28655 61228
rect 28382 61196 28408 61226
rect 28608 61196 28655 61226
rect 28639 61194 28655 61196
rect 28689 61194 28705 61228
rect 28639 61178 28705 61194
rect 28639 60918 28705 60934
rect 28639 60916 28655 60918
rect 28382 60886 28408 60916
rect 28608 60886 28655 60916
rect 28639 60884 28655 60886
rect 28689 60884 28705 60918
rect 28639 60868 28705 60884
rect 32812 61228 32878 61244
rect 32812 61194 32828 61228
rect 32862 61226 32878 61228
rect 32862 61196 32900 61226
rect 33100 61196 33126 61226
rect 32862 61194 32878 61196
rect 32812 61178 32878 61194
rect 32812 60918 32878 60934
rect 32812 60884 32828 60918
rect 32862 60916 32878 60918
rect 32862 60886 32900 60916
rect 33100 60886 33126 60916
rect 32862 60884 32878 60886
rect 32812 60868 32878 60884
rect 33629 61228 33695 61244
rect 33629 61226 33645 61228
rect 33372 61196 33398 61226
rect 33598 61196 33645 61226
rect 33629 61194 33645 61196
rect 33679 61194 33695 61228
rect 33629 61178 33695 61194
rect 33629 60918 33695 60934
rect 33629 60916 33645 60918
rect 33372 60886 33398 60916
rect 33598 60886 33645 60916
rect 33629 60884 33645 60886
rect 33679 60884 33695 60918
rect 33629 60868 33695 60884
rect 37802 61228 37868 61244
rect 37802 61194 37818 61228
rect 37852 61226 37868 61228
rect 37852 61196 37890 61226
rect 38090 61196 38116 61226
rect 37852 61194 37868 61196
rect 37802 61178 37868 61194
rect 37802 60918 37868 60934
rect 37802 60884 37818 60918
rect 37852 60916 37868 60918
rect 37852 60886 37890 60916
rect 38090 60886 38116 60916
rect 37852 60884 37868 60886
rect 37802 60868 37868 60884
rect 38619 61228 38685 61244
rect 38619 61226 38635 61228
rect 38362 61196 38388 61226
rect 38588 61196 38635 61226
rect 38619 61194 38635 61196
rect 38669 61194 38685 61228
rect 38619 61178 38685 61194
rect 38619 60918 38685 60934
rect 38619 60916 38635 60918
rect 38362 60886 38388 60916
rect 38588 60886 38635 60916
rect 38619 60884 38635 60886
rect 38669 60884 38685 60918
rect 38619 60868 38685 60884
rect 42792 61228 42858 61244
rect 42792 61194 42808 61228
rect 42842 61226 42858 61228
rect 42842 61196 42880 61226
rect 43080 61196 43106 61226
rect 42842 61194 42858 61196
rect 42792 61178 42858 61194
rect 42792 60918 42858 60934
rect 42792 60884 42808 60918
rect 42842 60916 42858 60918
rect 42842 60886 42880 60916
rect 43080 60886 43106 60916
rect 42842 60884 42858 60886
rect 42792 60868 42858 60884
rect 43609 61228 43675 61244
rect 43609 61226 43625 61228
rect 43352 61196 43378 61226
rect 43578 61196 43625 61226
rect 43609 61194 43625 61196
rect 43659 61194 43675 61228
rect 43609 61178 43675 61194
rect 43609 60918 43675 60934
rect 43609 60916 43625 60918
rect 43352 60886 43378 60916
rect 43578 60886 43625 60916
rect 43609 60884 43625 60886
rect 43659 60884 43675 60918
rect 43609 60868 43675 60884
rect 47782 61228 47848 61244
rect 47782 61194 47798 61228
rect 47832 61226 47848 61228
rect 47832 61196 47870 61226
rect 48070 61196 48096 61226
rect 47832 61194 47848 61196
rect 47782 61178 47848 61194
rect 47782 60918 47848 60934
rect 47782 60884 47798 60918
rect 47832 60916 47848 60918
rect 47832 60886 47870 60916
rect 48070 60886 48096 60916
rect 47832 60884 47848 60886
rect 47782 60868 47848 60884
rect 48599 61228 48665 61244
rect 48599 61226 48615 61228
rect 48342 61196 48368 61226
rect 48568 61196 48615 61226
rect 48599 61194 48615 61196
rect 48649 61194 48665 61228
rect 48599 61178 48665 61194
rect 48599 60918 48665 60934
rect 48599 60916 48615 60918
rect 48342 60886 48368 60916
rect 48568 60886 48615 60916
rect 48599 60884 48615 60886
rect 48649 60884 48665 60918
rect 48599 60868 48665 60884
rect 52772 61228 52838 61244
rect 52772 61194 52788 61228
rect 52822 61226 52838 61228
rect 52822 61196 52860 61226
rect 53060 61196 53086 61226
rect 52822 61194 52838 61196
rect 52772 61178 52838 61194
rect 52772 60918 52838 60934
rect 52772 60884 52788 60918
rect 52822 60916 52838 60918
rect 52822 60886 52860 60916
rect 53060 60886 53086 60916
rect 52822 60884 52838 60886
rect 52772 60868 52838 60884
rect 53589 61228 53655 61244
rect 53589 61226 53605 61228
rect 53332 61196 53358 61226
rect 53558 61196 53605 61226
rect 53589 61194 53605 61196
rect 53639 61194 53655 61228
rect 53589 61178 53655 61194
rect 53589 60918 53655 60934
rect 53589 60916 53605 60918
rect 53332 60886 53358 60916
rect 53558 60886 53605 60916
rect 53589 60884 53605 60886
rect 53639 60884 53655 60918
rect 53589 60868 53655 60884
rect 57762 61228 57828 61244
rect 57762 61194 57778 61228
rect 57812 61226 57828 61228
rect 57812 61196 57850 61226
rect 58050 61196 58076 61226
rect 57812 61194 57828 61196
rect 57762 61178 57828 61194
rect 57762 60918 57828 60934
rect 57762 60884 57778 60918
rect 57812 60916 57828 60918
rect 57812 60886 57850 60916
rect 58050 60886 58076 60916
rect 57812 60884 57828 60886
rect 57762 60868 57828 60884
rect 58579 61228 58645 61244
rect 58579 61226 58595 61228
rect 58322 61196 58348 61226
rect 58548 61196 58595 61226
rect 58579 61194 58595 61196
rect 58629 61194 58645 61228
rect 58579 61178 58645 61194
rect 58579 60918 58645 60934
rect 58579 60916 58595 60918
rect 58322 60886 58348 60916
rect 58548 60886 58595 60916
rect 58579 60884 58595 60886
rect 58629 60884 58645 60918
rect 58579 60868 58645 60884
rect 62752 61228 62818 61244
rect 62752 61194 62768 61228
rect 62802 61226 62818 61228
rect 62802 61196 62840 61226
rect 63040 61196 63066 61226
rect 62802 61194 62818 61196
rect 62752 61178 62818 61194
rect 62752 60918 62818 60934
rect 62752 60884 62768 60918
rect 62802 60916 62818 60918
rect 62802 60886 62840 60916
rect 63040 60886 63066 60916
rect 62802 60884 62818 60886
rect 62752 60868 62818 60884
rect 63569 61228 63635 61244
rect 63569 61226 63585 61228
rect 63312 61196 63338 61226
rect 63538 61196 63585 61226
rect 63569 61194 63585 61196
rect 63619 61194 63635 61228
rect 63569 61178 63635 61194
rect 63569 60918 63635 60934
rect 63569 60916 63585 60918
rect 63312 60886 63338 60916
rect 63538 60886 63585 60916
rect 63569 60884 63585 60886
rect 63619 60884 63635 60918
rect 63569 60868 63635 60884
rect 67742 61228 67808 61244
rect 67742 61194 67758 61228
rect 67792 61226 67808 61228
rect 67792 61196 67830 61226
rect 68030 61196 68056 61226
rect 67792 61194 67808 61196
rect 67742 61178 67808 61194
rect 67742 60918 67808 60934
rect 67742 60884 67758 60918
rect 67792 60916 67808 60918
rect 67792 60886 67830 60916
rect 68030 60886 68056 60916
rect 67792 60884 67808 60886
rect 67742 60868 67808 60884
rect 68559 61228 68625 61244
rect 68559 61226 68575 61228
rect 68302 61196 68328 61226
rect 68528 61196 68575 61226
rect 68559 61194 68575 61196
rect 68609 61194 68625 61228
rect 68559 61178 68625 61194
rect 68559 60918 68625 60934
rect 68559 60916 68575 60918
rect 68302 60886 68328 60916
rect 68528 60886 68575 60916
rect 68559 60884 68575 60886
rect 68609 60884 68625 60918
rect 68559 60868 68625 60884
rect 72732 61228 72798 61244
rect 72732 61194 72748 61228
rect 72782 61226 72798 61228
rect 72782 61196 72820 61226
rect 73020 61196 73046 61226
rect 72782 61194 72798 61196
rect 72732 61178 72798 61194
rect 72732 60918 72798 60934
rect 72732 60884 72748 60918
rect 72782 60916 72798 60918
rect 72782 60886 72820 60916
rect 73020 60886 73046 60916
rect 72782 60884 72798 60886
rect 72732 60868 72798 60884
rect 73549 61228 73615 61244
rect 73549 61226 73565 61228
rect 73292 61196 73318 61226
rect 73518 61196 73565 61226
rect 73549 61194 73565 61196
rect 73599 61194 73615 61228
rect 73549 61178 73615 61194
rect 73549 60918 73615 60934
rect 73549 60916 73565 60918
rect 73292 60886 73318 60916
rect 73518 60886 73565 60916
rect 73549 60884 73565 60886
rect 73599 60884 73615 60918
rect 73549 60868 73615 60884
rect 77722 61228 77788 61244
rect 77722 61194 77738 61228
rect 77772 61226 77788 61228
rect 77772 61196 77810 61226
rect 78010 61196 78036 61226
rect 77772 61194 77788 61196
rect 77722 61178 77788 61194
rect 77722 60918 77788 60934
rect 77722 60884 77738 60918
rect 77772 60916 77788 60918
rect 77772 60886 77810 60916
rect 78010 60886 78036 60916
rect 77772 60884 77788 60886
rect 77722 60868 77788 60884
rect 78539 61228 78605 61244
rect 78539 61226 78555 61228
rect 78282 61196 78308 61226
rect 78508 61196 78555 61226
rect 78539 61194 78555 61196
rect 78589 61194 78605 61228
rect 78539 61178 78605 61194
rect 78539 60918 78605 60934
rect 78539 60916 78555 60918
rect 78282 60886 78308 60916
rect 78508 60886 78555 60916
rect 78539 60884 78555 60886
rect 78589 60884 78605 60918
rect 78539 60868 78605 60884
rect 2872 59518 2938 59534
rect 2872 59484 2888 59518
rect 2922 59516 2938 59518
rect 2922 59486 2960 59516
rect 3160 59486 3186 59516
rect 2922 59484 2938 59486
rect 2872 59468 2938 59484
rect 2872 59208 2938 59224
rect 2872 59174 2888 59208
rect 2922 59206 2938 59208
rect 2922 59176 2960 59206
rect 3160 59176 3186 59206
rect 2922 59174 2938 59176
rect 2872 59158 2938 59174
rect 3689 59518 3755 59534
rect 3689 59516 3705 59518
rect 3432 59486 3458 59516
rect 3658 59486 3705 59516
rect 3689 59484 3705 59486
rect 3739 59484 3755 59518
rect 3689 59468 3755 59484
rect 3689 59208 3755 59224
rect 3689 59206 3705 59208
rect 3432 59176 3458 59206
rect 3658 59176 3705 59206
rect 3689 59174 3705 59176
rect 3739 59174 3755 59208
rect 3689 59158 3755 59174
rect 7862 59518 7928 59534
rect 7862 59484 7878 59518
rect 7912 59516 7928 59518
rect 7912 59486 7950 59516
rect 8150 59486 8176 59516
rect 7912 59484 7928 59486
rect 7862 59468 7928 59484
rect 7862 59208 7928 59224
rect 7862 59174 7878 59208
rect 7912 59206 7928 59208
rect 7912 59176 7950 59206
rect 8150 59176 8176 59206
rect 7912 59174 7928 59176
rect 7862 59158 7928 59174
rect 8679 59518 8745 59534
rect 8679 59516 8695 59518
rect 8422 59486 8448 59516
rect 8648 59486 8695 59516
rect 8679 59484 8695 59486
rect 8729 59484 8745 59518
rect 8679 59468 8745 59484
rect 8679 59208 8745 59224
rect 8679 59206 8695 59208
rect 8422 59176 8448 59206
rect 8648 59176 8695 59206
rect 8679 59174 8695 59176
rect 8729 59174 8745 59208
rect 8679 59158 8745 59174
rect 12852 59518 12918 59534
rect 12852 59484 12868 59518
rect 12902 59516 12918 59518
rect 12902 59486 12940 59516
rect 13140 59486 13166 59516
rect 12902 59484 12918 59486
rect 12852 59468 12918 59484
rect 12852 59208 12918 59224
rect 12852 59174 12868 59208
rect 12902 59206 12918 59208
rect 12902 59176 12940 59206
rect 13140 59176 13166 59206
rect 12902 59174 12918 59176
rect 12852 59158 12918 59174
rect 13669 59518 13735 59534
rect 13669 59516 13685 59518
rect 13412 59486 13438 59516
rect 13638 59486 13685 59516
rect 13669 59484 13685 59486
rect 13719 59484 13735 59518
rect 13669 59468 13735 59484
rect 13669 59208 13735 59224
rect 13669 59206 13685 59208
rect 13412 59176 13438 59206
rect 13638 59176 13685 59206
rect 13669 59174 13685 59176
rect 13719 59174 13735 59208
rect 13669 59158 13735 59174
rect 17842 59518 17908 59534
rect 17842 59484 17858 59518
rect 17892 59516 17908 59518
rect 17892 59486 17930 59516
rect 18130 59486 18156 59516
rect 17892 59484 17908 59486
rect 17842 59468 17908 59484
rect 17842 59208 17908 59224
rect 17842 59174 17858 59208
rect 17892 59206 17908 59208
rect 17892 59176 17930 59206
rect 18130 59176 18156 59206
rect 17892 59174 17908 59176
rect 17842 59158 17908 59174
rect 18659 59518 18725 59534
rect 18659 59516 18675 59518
rect 18402 59486 18428 59516
rect 18628 59486 18675 59516
rect 18659 59484 18675 59486
rect 18709 59484 18725 59518
rect 18659 59468 18725 59484
rect 18659 59208 18725 59224
rect 18659 59206 18675 59208
rect 18402 59176 18428 59206
rect 18628 59176 18675 59206
rect 18659 59174 18675 59176
rect 18709 59174 18725 59208
rect 18659 59158 18725 59174
rect 22832 59518 22898 59534
rect 22832 59484 22848 59518
rect 22882 59516 22898 59518
rect 22882 59486 22920 59516
rect 23120 59486 23146 59516
rect 22882 59484 22898 59486
rect 22832 59468 22898 59484
rect 22832 59208 22898 59224
rect 22832 59174 22848 59208
rect 22882 59206 22898 59208
rect 22882 59176 22920 59206
rect 23120 59176 23146 59206
rect 22882 59174 22898 59176
rect 22832 59158 22898 59174
rect 23649 59518 23715 59534
rect 23649 59516 23665 59518
rect 23392 59486 23418 59516
rect 23618 59486 23665 59516
rect 23649 59484 23665 59486
rect 23699 59484 23715 59518
rect 23649 59468 23715 59484
rect 23649 59208 23715 59224
rect 23649 59206 23665 59208
rect 23392 59176 23418 59206
rect 23618 59176 23665 59206
rect 23649 59174 23665 59176
rect 23699 59174 23715 59208
rect 23649 59158 23715 59174
rect 27822 59518 27888 59534
rect 27822 59484 27838 59518
rect 27872 59516 27888 59518
rect 27872 59486 27910 59516
rect 28110 59486 28136 59516
rect 27872 59484 27888 59486
rect 27822 59468 27888 59484
rect 27822 59208 27888 59224
rect 27822 59174 27838 59208
rect 27872 59206 27888 59208
rect 27872 59176 27910 59206
rect 28110 59176 28136 59206
rect 27872 59174 27888 59176
rect 27822 59158 27888 59174
rect 28639 59518 28705 59534
rect 28639 59516 28655 59518
rect 28382 59486 28408 59516
rect 28608 59486 28655 59516
rect 28639 59484 28655 59486
rect 28689 59484 28705 59518
rect 28639 59468 28705 59484
rect 28639 59208 28705 59224
rect 28639 59206 28655 59208
rect 28382 59176 28408 59206
rect 28608 59176 28655 59206
rect 28639 59174 28655 59176
rect 28689 59174 28705 59208
rect 28639 59158 28705 59174
rect 32812 59518 32878 59534
rect 32812 59484 32828 59518
rect 32862 59516 32878 59518
rect 32862 59486 32900 59516
rect 33100 59486 33126 59516
rect 32862 59484 32878 59486
rect 32812 59468 32878 59484
rect 32812 59208 32878 59224
rect 32812 59174 32828 59208
rect 32862 59206 32878 59208
rect 32862 59176 32900 59206
rect 33100 59176 33126 59206
rect 32862 59174 32878 59176
rect 32812 59158 32878 59174
rect 33629 59518 33695 59534
rect 33629 59516 33645 59518
rect 33372 59486 33398 59516
rect 33598 59486 33645 59516
rect 33629 59484 33645 59486
rect 33679 59484 33695 59518
rect 33629 59468 33695 59484
rect 33629 59208 33695 59224
rect 33629 59206 33645 59208
rect 33372 59176 33398 59206
rect 33598 59176 33645 59206
rect 33629 59174 33645 59176
rect 33679 59174 33695 59208
rect 33629 59158 33695 59174
rect 37802 59518 37868 59534
rect 37802 59484 37818 59518
rect 37852 59516 37868 59518
rect 37852 59486 37890 59516
rect 38090 59486 38116 59516
rect 37852 59484 37868 59486
rect 37802 59468 37868 59484
rect 37802 59208 37868 59224
rect 37802 59174 37818 59208
rect 37852 59206 37868 59208
rect 37852 59176 37890 59206
rect 38090 59176 38116 59206
rect 37852 59174 37868 59176
rect 37802 59158 37868 59174
rect 38619 59518 38685 59534
rect 38619 59516 38635 59518
rect 38362 59486 38388 59516
rect 38588 59486 38635 59516
rect 38619 59484 38635 59486
rect 38669 59484 38685 59518
rect 38619 59468 38685 59484
rect 38619 59208 38685 59224
rect 38619 59206 38635 59208
rect 38362 59176 38388 59206
rect 38588 59176 38635 59206
rect 38619 59174 38635 59176
rect 38669 59174 38685 59208
rect 38619 59158 38685 59174
rect 42792 59518 42858 59534
rect 42792 59484 42808 59518
rect 42842 59516 42858 59518
rect 42842 59486 42880 59516
rect 43080 59486 43106 59516
rect 42842 59484 42858 59486
rect 42792 59468 42858 59484
rect 42792 59208 42858 59224
rect 42792 59174 42808 59208
rect 42842 59206 42858 59208
rect 42842 59176 42880 59206
rect 43080 59176 43106 59206
rect 42842 59174 42858 59176
rect 42792 59158 42858 59174
rect 43609 59518 43675 59534
rect 43609 59516 43625 59518
rect 43352 59486 43378 59516
rect 43578 59486 43625 59516
rect 43609 59484 43625 59486
rect 43659 59484 43675 59518
rect 43609 59468 43675 59484
rect 43609 59208 43675 59224
rect 43609 59206 43625 59208
rect 43352 59176 43378 59206
rect 43578 59176 43625 59206
rect 43609 59174 43625 59176
rect 43659 59174 43675 59208
rect 43609 59158 43675 59174
rect 47782 59518 47848 59534
rect 47782 59484 47798 59518
rect 47832 59516 47848 59518
rect 47832 59486 47870 59516
rect 48070 59486 48096 59516
rect 47832 59484 47848 59486
rect 47782 59468 47848 59484
rect 47782 59208 47848 59224
rect 47782 59174 47798 59208
rect 47832 59206 47848 59208
rect 47832 59176 47870 59206
rect 48070 59176 48096 59206
rect 47832 59174 47848 59176
rect 47782 59158 47848 59174
rect 48599 59518 48665 59534
rect 48599 59516 48615 59518
rect 48342 59486 48368 59516
rect 48568 59486 48615 59516
rect 48599 59484 48615 59486
rect 48649 59484 48665 59518
rect 48599 59468 48665 59484
rect 48599 59208 48665 59224
rect 48599 59206 48615 59208
rect 48342 59176 48368 59206
rect 48568 59176 48615 59206
rect 48599 59174 48615 59176
rect 48649 59174 48665 59208
rect 48599 59158 48665 59174
rect 52772 59518 52838 59534
rect 52772 59484 52788 59518
rect 52822 59516 52838 59518
rect 52822 59486 52860 59516
rect 53060 59486 53086 59516
rect 52822 59484 52838 59486
rect 52772 59468 52838 59484
rect 52772 59208 52838 59224
rect 52772 59174 52788 59208
rect 52822 59206 52838 59208
rect 52822 59176 52860 59206
rect 53060 59176 53086 59206
rect 52822 59174 52838 59176
rect 52772 59158 52838 59174
rect 53589 59518 53655 59534
rect 53589 59516 53605 59518
rect 53332 59486 53358 59516
rect 53558 59486 53605 59516
rect 53589 59484 53605 59486
rect 53639 59484 53655 59518
rect 53589 59468 53655 59484
rect 53589 59208 53655 59224
rect 53589 59206 53605 59208
rect 53332 59176 53358 59206
rect 53558 59176 53605 59206
rect 53589 59174 53605 59176
rect 53639 59174 53655 59208
rect 53589 59158 53655 59174
rect 57762 59518 57828 59534
rect 57762 59484 57778 59518
rect 57812 59516 57828 59518
rect 57812 59486 57850 59516
rect 58050 59486 58076 59516
rect 57812 59484 57828 59486
rect 57762 59468 57828 59484
rect 57762 59208 57828 59224
rect 57762 59174 57778 59208
rect 57812 59206 57828 59208
rect 57812 59176 57850 59206
rect 58050 59176 58076 59206
rect 57812 59174 57828 59176
rect 57762 59158 57828 59174
rect 58579 59518 58645 59534
rect 58579 59516 58595 59518
rect 58322 59486 58348 59516
rect 58548 59486 58595 59516
rect 58579 59484 58595 59486
rect 58629 59484 58645 59518
rect 58579 59468 58645 59484
rect 58579 59208 58645 59224
rect 58579 59206 58595 59208
rect 58322 59176 58348 59206
rect 58548 59176 58595 59206
rect 58579 59174 58595 59176
rect 58629 59174 58645 59208
rect 58579 59158 58645 59174
rect 62752 59518 62818 59534
rect 62752 59484 62768 59518
rect 62802 59516 62818 59518
rect 62802 59486 62840 59516
rect 63040 59486 63066 59516
rect 62802 59484 62818 59486
rect 62752 59468 62818 59484
rect 62752 59208 62818 59224
rect 62752 59174 62768 59208
rect 62802 59206 62818 59208
rect 62802 59176 62840 59206
rect 63040 59176 63066 59206
rect 62802 59174 62818 59176
rect 62752 59158 62818 59174
rect 63569 59518 63635 59534
rect 63569 59516 63585 59518
rect 63312 59486 63338 59516
rect 63538 59486 63585 59516
rect 63569 59484 63585 59486
rect 63619 59484 63635 59518
rect 63569 59468 63635 59484
rect 63569 59208 63635 59224
rect 63569 59206 63585 59208
rect 63312 59176 63338 59206
rect 63538 59176 63585 59206
rect 63569 59174 63585 59176
rect 63619 59174 63635 59208
rect 63569 59158 63635 59174
rect 67742 59518 67808 59534
rect 67742 59484 67758 59518
rect 67792 59516 67808 59518
rect 67792 59486 67830 59516
rect 68030 59486 68056 59516
rect 67792 59484 67808 59486
rect 67742 59468 67808 59484
rect 67742 59208 67808 59224
rect 67742 59174 67758 59208
rect 67792 59206 67808 59208
rect 67792 59176 67830 59206
rect 68030 59176 68056 59206
rect 67792 59174 67808 59176
rect 67742 59158 67808 59174
rect 68559 59518 68625 59534
rect 68559 59516 68575 59518
rect 68302 59486 68328 59516
rect 68528 59486 68575 59516
rect 68559 59484 68575 59486
rect 68609 59484 68625 59518
rect 68559 59468 68625 59484
rect 68559 59208 68625 59224
rect 68559 59206 68575 59208
rect 68302 59176 68328 59206
rect 68528 59176 68575 59206
rect 68559 59174 68575 59176
rect 68609 59174 68625 59208
rect 68559 59158 68625 59174
rect 72732 59518 72798 59534
rect 72732 59484 72748 59518
rect 72782 59516 72798 59518
rect 72782 59486 72820 59516
rect 73020 59486 73046 59516
rect 72782 59484 72798 59486
rect 72732 59468 72798 59484
rect 72732 59208 72798 59224
rect 72732 59174 72748 59208
rect 72782 59206 72798 59208
rect 72782 59176 72820 59206
rect 73020 59176 73046 59206
rect 72782 59174 72798 59176
rect 72732 59158 72798 59174
rect 73549 59518 73615 59534
rect 73549 59516 73565 59518
rect 73292 59486 73318 59516
rect 73518 59486 73565 59516
rect 73549 59484 73565 59486
rect 73599 59484 73615 59518
rect 73549 59468 73615 59484
rect 73549 59208 73615 59224
rect 73549 59206 73565 59208
rect 73292 59176 73318 59206
rect 73518 59176 73565 59206
rect 73549 59174 73565 59176
rect 73599 59174 73615 59208
rect 73549 59158 73615 59174
rect 77722 59518 77788 59534
rect 77722 59484 77738 59518
rect 77772 59516 77788 59518
rect 77772 59486 77810 59516
rect 78010 59486 78036 59516
rect 77772 59484 77788 59486
rect 77722 59468 77788 59484
rect 77722 59208 77788 59224
rect 77722 59174 77738 59208
rect 77772 59206 77788 59208
rect 77772 59176 77810 59206
rect 78010 59176 78036 59206
rect 77772 59174 77788 59176
rect 77722 59158 77788 59174
rect 78539 59518 78605 59534
rect 78539 59516 78555 59518
rect 78282 59486 78308 59516
rect 78508 59486 78555 59516
rect 78539 59484 78555 59486
rect 78589 59484 78605 59518
rect 78539 59468 78605 59484
rect 78539 59208 78605 59224
rect 78539 59206 78555 59208
rect 78282 59176 78308 59206
rect 78508 59176 78555 59206
rect 78539 59174 78555 59176
rect 78589 59174 78605 59208
rect 78539 59158 78605 59174
rect 2872 57808 2938 57824
rect 2872 57774 2888 57808
rect 2922 57806 2938 57808
rect 2922 57776 2960 57806
rect 3160 57776 3186 57806
rect 2922 57774 2938 57776
rect 2872 57758 2938 57774
rect 2872 57498 2938 57514
rect 2872 57464 2888 57498
rect 2922 57496 2938 57498
rect 2922 57466 2960 57496
rect 3160 57466 3186 57496
rect 2922 57464 2938 57466
rect 2872 57448 2938 57464
rect 3689 57808 3755 57824
rect 3689 57806 3705 57808
rect 3432 57776 3458 57806
rect 3658 57776 3705 57806
rect 3689 57774 3705 57776
rect 3739 57774 3755 57808
rect 3689 57758 3755 57774
rect 3689 57498 3755 57514
rect 3689 57496 3705 57498
rect 3432 57466 3458 57496
rect 3658 57466 3705 57496
rect 3689 57464 3705 57466
rect 3739 57464 3755 57498
rect 3689 57448 3755 57464
rect 7862 57808 7928 57824
rect 7862 57774 7878 57808
rect 7912 57806 7928 57808
rect 7912 57776 7950 57806
rect 8150 57776 8176 57806
rect 7912 57774 7928 57776
rect 7862 57758 7928 57774
rect 7862 57498 7928 57514
rect 7862 57464 7878 57498
rect 7912 57496 7928 57498
rect 7912 57466 7950 57496
rect 8150 57466 8176 57496
rect 7912 57464 7928 57466
rect 7862 57448 7928 57464
rect 8679 57808 8745 57824
rect 8679 57806 8695 57808
rect 8422 57776 8448 57806
rect 8648 57776 8695 57806
rect 8679 57774 8695 57776
rect 8729 57774 8745 57808
rect 8679 57758 8745 57774
rect 8679 57498 8745 57514
rect 8679 57496 8695 57498
rect 8422 57466 8448 57496
rect 8648 57466 8695 57496
rect 8679 57464 8695 57466
rect 8729 57464 8745 57498
rect 8679 57448 8745 57464
rect 12852 57808 12918 57824
rect 12852 57774 12868 57808
rect 12902 57806 12918 57808
rect 12902 57776 12940 57806
rect 13140 57776 13166 57806
rect 12902 57774 12918 57776
rect 12852 57758 12918 57774
rect 12852 57498 12918 57514
rect 12852 57464 12868 57498
rect 12902 57496 12918 57498
rect 12902 57466 12940 57496
rect 13140 57466 13166 57496
rect 12902 57464 12918 57466
rect 12852 57448 12918 57464
rect 13669 57808 13735 57824
rect 13669 57806 13685 57808
rect 13412 57776 13438 57806
rect 13638 57776 13685 57806
rect 13669 57774 13685 57776
rect 13719 57774 13735 57808
rect 13669 57758 13735 57774
rect 13669 57498 13735 57514
rect 13669 57496 13685 57498
rect 13412 57466 13438 57496
rect 13638 57466 13685 57496
rect 13669 57464 13685 57466
rect 13719 57464 13735 57498
rect 13669 57448 13735 57464
rect 17842 57808 17908 57824
rect 17842 57774 17858 57808
rect 17892 57806 17908 57808
rect 17892 57776 17930 57806
rect 18130 57776 18156 57806
rect 17892 57774 17908 57776
rect 17842 57758 17908 57774
rect 17842 57498 17908 57514
rect 17842 57464 17858 57498
rect 17892 57496 17908 57498
rect 17892 57466 17930 57496
rect 18130 57466 18156 57496
rect 17892 57464 17908 57466
rect 17842 57448 17908 57464
rect 18659 57808 18725 57824
rect 18659 57806 18675 57808
rect 18402 57776 18428 57806
rect 18628 57776 18675 57806
rect 18659 57774 18675 57776
rect 18709 57774 18725 57808
rect 18659 57758 18725 57774
rect 18659 57498 18725 57514
rect 18659 57496 18675 57498
rect 18402 57466 18428 57496
rect 18628 57466 18675 57496
rect 18659 57464 18675 57466
rect 18709 57464 18725 57498
rect 18659 57448 18725 57464
rect 22832 57808 22898 57824
rect 22832 57774 22848 57808
rect 22882 57806 22898 57808
rect 22882 57776 22920 57806
rect 23120 57776 23146 57806
rect 22882 57774 22898 57776
rect 22832 57758 22898 57774
rect 22832 57498 22898 57514
rect 22832 57464 22848 57498
rect 22882 57496 22898 57498
rect 22882 57466 22920 57496
rect 23120 57466 23146 57496
rect 22882 57464 22898 57466
rect 22832 57448 22898 57464
rect 23649 57808 23715 57824
rect 23649 57806 23665 57808
rect 23392 57776 23418 57806
rect 23618 57776 23665 57806
rect 23649 57774 23665 57776
rect 23699 57774 23715 57808
rect 23649 57758 23715 57774
rect 23649 57498 23715 57514
rect 23649 57496 23665 57498
rect 23392 57466 23418 57496
rect 23618 57466 23665 57496
rect 23649 57464 23665 57466
rect 23699 57464 23715 57498
rect 23649 57448 23715 57464
rect 27822 57808 27888 57824
rect 27822 57774 27838 57808
rect 27872 57806 27888 57808
rect 27872 57776 27910 57806
rect 28110 57776 28136 57806
rect 27872 57774 27888 57776
rect 27822 57758 27888 57774
rect 27822 57498 27888 57514
rect 27822 57464 27838 57498
rect 27872 57496 27888 57498
rect 27872 57466 27910 57496
rect 28110 57466 28136 57496
rect 27872 57464 27888 57466
rect 27822 57448 27888 57464
rect 28639 57808 28705 57824
rect 28639 57806 28655 57808
rect 28382 57776 28408 57806
rect 28608 57776 28655 57806
rect 28639 57774 28655 57776
rect 28689 57774 28705 57808
rect 28639 57758 28705 57774
rect 28639 57498 28705 57514
rect 28639 57496 28655 57498
rect 28382 57466 28408 57496
rect 28608 57466 28655 57496
rect 28639 57464 28655 57466
rect 28689 57464 28705 57498
rect 28639 57448 28705 57464
rect 32812 57808 32878 57824
rect 32812 57774 32828 57808
rect 32862 57806 32878 57808
rect 32862 57776 32900 57806
rect 33100 57776 33126 57806
rect 32862 57774 32878 57776
rect 32812 57758 32878 57774
rect 32812 57498 32878 57514
rect 32812 57464 32828 57498
rect 32862 57496 32878 57498
rect 32862 57466 32900 57496
rect 33100 57466 33126 57496
rect 32862 57464 32878 57466
rect 32812 57448 32878 57464
rect 33629 57808 33695 57824
rect 33629 57806 33645 57808
rect 33372 57776 33398 57806
rect 33598 57776 33645 57806
rect 33629 57774 33645 57776
rect 33679 57774 33695 57808
rect 33629 57758 33695 57774
rect 33629 57498 33695 57514
rect 33629 57496 33645 57498
rect 33372 57466 33398 57496
rect 33598 57466 33645 57496
rect 33629 57464 33645 57466
rect 33679 57464 33695 57498
rect 33629 57448 33695 57464
rect 37802 57808 37868 57824
rect 37802 57774 37818 57808
rect 37852 57806 37868 57808
rect 37852 57776 37890 57806
rect 38090 57776 38116 57806
rect 37852 57774 37868 57776
rect 37802 57758 37868 57774
rect 37802 57498 37868 57514
rect 37802 57464 37818 57498
rect 37852 57496 37868 57498
rect 37852 57466 37890 57496
rect 38090 57466 38116 57496
rect 37852 57464 37868 57466
rect 37802 57448 37868 57464
rect 38619 57808 38685 57824
rect 38619 57806 38635 57808
rect 38362 57776 38388 57806
rect 38588 57776 38635 57806
rect 38619 57774 38635 57776
rect 38669 57774 38685 57808
rect 38619 57758 38685 57774
rect 38619 57498 38685 57514
rect 38619 57496 38635 57498
rect 38362 57466 38388 57496
rect 38588 57466 38635 57496
rect 38619 57464 38635 57466
rect 38669 57464 38685 57498
rect 38619 57448 38685 57464
rect 42792 57808 42858 57824
rect 42792 57774 42808 57808
rect 42842 57806 42858 57808
rect 42842 57776 42880 57806
rect 43080 57776 43106 57806
rect 42842 57774 42858 57776
rect 42792 57758 42858 57774
rect 42792 57498 42858 57514
rect 42792 57464 42808 57498
rect 42842 57496 42858 57498
rect 42842 57466 42880 57496
rect 43080 57466 43106 57496
rect 42842 57464 42858 57466
rect 42792 57448 42858 57464
rect 43609 57808 43675 57824
rect 43609 57806 43625 57808
rect 43352 57776 43378 57806
rect 43578 57776 43625 57806
rect 43609 57774 43625 57776
rect 43659 57774 43675 57808
rect 43609 57758 43675 57774
rect 43609 57498 43675 57514
rect 43609 57496 43625 57498
rect 43352 57466 43378 57496
rect 43578 57466 43625 57496
rect 43609 57464 43625 57466
rect 43659 57464 43675 57498
rect 43609 57448 43675 57464
rect 47782 57808 47848 57824
rect 47782 57774 47798 57808
rect 47832 57806 47848 57808
rect 47832 57776 47870 57806
rect 48070 57776 48096 57806
rect 47832 57774 47848 57776
rect 47782 57758 47848 57774
rect 47782 57498 47848 57514
rect 47782 57464 47798 57498
rect 47832 57496 47848 57498
rect 47832 57466 47870 57496
rect 48070 57466 48096 57496
rect 47832 57464 47848 57466
rect 47782 57448 47848 57464
rect 48599 57808 48665 57824
rect 48599 57806 48615 57808
rect 48342 57776 48368 57806
rect 48568 57776 48615 57806
rect 48599 57774 48615 57776
rect 48649 57774 48665 57808
rect 48599 57758 48665 57774
rect 48599 57498 48665 57514
rect 48599 57496 48615 57498
rect 48342 57466 48368 57496
rect 48568 57466 48615 57496
rect 48599 57464 48615 57466
rect 48649 57464 48665 57498
rect 48599 57448 48665 57464
rect 52772 57808 52838 57824
rect 52772 57774 52788 57808
rect 52822 57806 52838 57808
rect 52822 57776 52860 57806
rect 53060 57776 53086 57806
rect 52822 57774 52838 57776
rect 52772 57758 52838 57774
rect 52772 57498 52838 57514
rect 52772 57464 52788 57498
rect 52822 57496 52838 57498
rect 52822 57466 52860 57496
rect 53060 57466 53086 57496
rect 52822 57464 52838 57466
rect 52772 57448 52838 57464
rect 53589 57808 53655 57824
rect 53589 57806 53605 57808
rect 53332 57776 53358 57806
rect 53558 57776 53605 57806
rect 53589 57774 53605 57776
rect 53639 57774 53655 57808
rect 53589 57758 53655 57774
rect 53589 57498 53655 57514
rect 53589 57496 53605 57498
rect 53332 57466 53358 57496
rect 53558 57466 53605 57496
rect 53589 57464 53605 57466
rect 53639 57464 53655 57498
rect 53589 57448 53655 57464
rect 57762 57808 57828 57824
rect 57762 57774 57778 57808
rect 57812 57806 57828 57808
rect 57812 57776 57850 57806
rect 58050 57776 58076 57806
rect 57812 57774 57828 57776
rect 57762 57758 57828 57774
rect 57762 57498 57828 57514
rect 57762 57464 57778 57498
rect 57812 57496 57828 57498
rect 57812 57466 57850 57496
rect 58050 57466 58076 57496
rect 57812 57464 57828 57466
rect 57762 57448 57828 57464
rect 58579 57808 58645 57824
rect 58579 57806 58595 57808
rect 58322 57776 58348 57806
rect 58548 57776 58595 57806
rect 58579 57774 58595 57776
rect 58629 57774 58645 57808
rect 58579 57758 58645 57774
rect 58579 57498 58645 57514
rect 58579 57496 58595 57498
rect 58322 57466 58348 57496
rect 58548 57466 58595 57496
rect 58579 57464 58595 57466
rect 58629 57464 58645 57498
rect 58579 57448 58645 57464
rect 62752 57808 62818 57824
rect 62752 57774 62768 57808
rect 62802 57806 62818 57808
rect 62802 57776 62840 57806
rect 63040 57776 63066 57806
rect 62802 57774 62818 57776
rect 62752 57758 62818 57774
rect 62752 57498 62818 57514
rect 62752 57464 62768 57498
rect 62802 57496 62818 57498
rect 62802 57466 62840 57496
rect 63040 57466 63066 57496
rect 62802 57464 62818 57466
rect 62752 57448 62818 57464
rect 63569 57808 63635 57824
rect 63569 57806 63585 57808
rect 63312 57776 63338 57806
rect 63538 57776 63585 57806
rect 63569 57774 63585 57776
rect 63619 57774 63635 57808
rect 63569 57758 63635 57774
rect 63569 57498 63635 57514
rect 63569 57496 63585 57498
rect 63312 57466 63338 57496
rect 63538 57466 63585 57496
rect 63569 57464 63585 57466
rect 63619 57464 63635 57498
rect 63569 57448 63635 57464
rect 67742 57808 67808 57824
rect 67742 57774 67758 57808
rect 67792 57806 67808 57808
rect 67792 57776 67830 57806
rect 68030 57776 68056 57806
rect 67792 57774 67808 57776
rect 67742 57758 67808 57774
rect 67742 57498 67808 57514
rect 67742 57464 67758 57498
rect 67792 57496 67808 57498
rect 67792 57466 67830 57496
rect 68030 57466 68056 57496
rect 67792 57464 67808 57466
rect 67742 57448 67808 57464
rect 68559 57808 68625 57824
rect 68559 57806 68575 57808
rect 68302 57776 68328 57806
rect 68528 57776 68575 57806
rect 68559 57774 68575 57776
rect 68609 57774 68625 57808
rect 68559 57758 68625 57774
rect 68559 57498 68625 57514
rect 68559 57496 68575 57498
rect 68302 57466 68328 57496
rect 68528 57466 68575 57496
rect 68559 57464 68575 57466
rect 68609 57464 68625 57498
rect 68559 57448 68625 57464
rect 72732 57808 72798 57824
rect 72732 57774 72748 57808
rect 72782 57806 72798 57808
rect 72782 57776 72820 57806
rect 73020 57776 73046 57806
rect 72782 57774 72798 57776
rect 72732 57758 72798 57774
rect 72732 57498 72798 57514
rect 72732 57464 72748 57498
rect 72782 57496 72798 57498
rect 72782 57466 72820 57496
rect 73020 57466 73046 57496
rect 72782 57464 72798 57466
rect 72732 57448 72798 57464
rect 73549 57808 73615 57824
rect 73549 57806 73565 57808
rect 73292 57776 73318 57806
rect 73518 57776 73565 57806
rect 73549 57774 73565 57776
rect 73599 57774 73615 57808
rect 73549 57758 73615 57774
rect 73549 57498 73615 57514
rect 73549 57496 73565 57498
rect 73292 57466 73318 57496
rect 73518 57466 73565 57496
rect 73549 57464 73565 57466
rect 73599 57464 73615 57498
rect 73549 57448 73615 57464
rect 77722 57808 77788 57824
rect 77722 57774 77738 57808
rect 77772 57806 77788 57808
rect 77772 57776 77810 57806
rect 78010 57776 78036 57806
rect 77772 57774 77788 57776
rect 77722 57758 77788 57774
rect 77722 57498 77788 57514
rect 77722 57464 77738 57498
rect 77772 57496 77788 57498
rect 77772 57466 77810 57496
rect 78010 57466 78036 57496
rect 77772 57464 77788 57466
rect 77722 57448 77788 57464
rect 78539 57808 78605 57824
rect 78539 57806 78555 57808
rect 78282 57776 78308 57806
rect 78508 57776 78555 57806
rect 78539 57774 78555 57776
rect 78589 57774 78605 57808
rect 78539 57758 78605 57774
rect 78539 57498 78605 57514
rect 78539 57496 78555 57498
rect 78282 57466 78308 57496
rect 78508 57466 78555 57496
rect 78539 57464 78555 57466
rect 78589 57464 78605 57498
rect 78539 57448 78605 57464
rect 2872 56098 2938 56114
rect 2872 56064 2888 56098
rect 2922 56096 2938 56098
rect 2922 56066 2960 56096
rect 3160 56066 3186 56096
rect 2922 56064 2938 56066
rect 2872 56048 2938 56064
rect 2872 55788 2938 55804
rect 2872 55754 2888 55788
rect 2922 55786 2938 55788
rect 2922 55756 2960 55786
rect 3160 55756 3186 55786
rect 2922 55754 2938 55756
rect 2872 55738 2938 55754
rect 3689 56098 3755 56114
rect 3689 56096 3705 56098
rect 3432 56066 3458 56096
rect 3658 56066 3705 56096
rect 3689 56064 3705 56066
rect 3739 56064 3755 56098
rect 3689 56048 3755 56064
rect 3689 55788 3755 55804
rect 3689 55786 3705 55788
rect 3432 55756 3458 55786
rect 3658 55756 3705 55786
rect 3689 55754 3705 55756
rect 3739 55754 3755 55788
rect 3689 55738 3755 55754
rect 7862 56098 7928 56114
rect 7862 56064 7878 56098
rect 7912 56096 7928 56098
rect 7912 56066 7950 56096
rect 8150 56066 8176 56096
rect 7912 56064 7928 56066
rect 7862 56048 7928 56064
rect 7862 55788 7928 55804
rect 7862 55754 7878 55788
rect 7912 55786 7928 55788
rect 7912 55756 7950 55786
rect 8150 55756 8176 55786
rect 7912 55754 7928 55756
rect 7862 55738 7928 55754
rect 8679 56098 8745 56114
rect 8679 56096 8695 56098
rect 8422 56066 8448 56096
rect 8648 56066 8695 56096
rect 8679 56064 8695 56066
rect 8729 56064 8745 56098
rect 8679 56048 8745 56064
rect 8679 55788 8745 55804
rect 8679 55786 8695 55788
rect 8422 55756 8448 55786
rect 8648 55756 8695 55786
rect 8679 55754 8695 55756
rect 8729 55754 8745 55788
rect 8679 55738 8745 55754
rect 12852 56098 12918 56114
rect 12852 56064 12868 56098
rect 12902 56096 12918 56098
rect 12902 56066 12940 56096
rect 13140 56066 13166 56096
rect 12902 56064 12918 56066
rect 12852 56048 12918 56064
rect 12852 55788 12918 55804
rect 12852 55754 12868 55788
rect 12902 55786 12918 55788
rect 12902 55756 12940 55786
rect 13140 55756 13166 55786
rect 12902 55754 12918 55756
rect 12852 55738 12918 55754
rect 13669 56098 13735 56114
rect 13669 56096 13685 56098
rect 13412 56066 13438 56096
rect 13638 56066 13685 56096
rect 13669 56064 13685 56066
rect 13719 56064 13735 56098
rect 13669 56048 13735 56064
rect 13669 55788 13735 55804
rect 13669 55786 13685 55788
rect 13412 55756 13438 55786
rect 13638 55756 13685 55786
rect 13669 55754 13685 55756
rect 13719 55754 13735 55788
rect 13669 55738 13735 55754
rect 17842 56098 17908 56114
rect 17842 56064 17858 56098
rect 17892 56096 17908 56098
rect 17892 56066 17930 56096
rect 18130 56066 18156 56096
rect 17892 56064 17908 56066
rect 17842 56048 17908 56064
rect 17842 55788 17908 55804
rect 17842 55754 17858 55788
rect 17892 55786 17908 55788
rect 17892 55756 17930 55786
rect 18130 55756 18156 55786
rect 17892 55754 17908 55756
rect 17842 55738 17908 55754
rect 18659 56098 18725 56114
rect 18659 56096 18675 56098
rect 18402 56066 18428 56096
rect 18628 56066 18675 56096
rect 18659 56064 18675 56066
rect 18709 56064 18725 56098
rect 18659 56048 18725 56064
rect 18659 55788 18725 55804
rect 18659 55786 18675 55788
rect 18402 55756 18428 55786
rect 18628 55756 18675 55786
rect 18659 55754 18675 55756
rect 18709 55754 18725 55788
rect 18659 55738 18725 55754
rect 22832 56098 22898 56114
rect 22832 56064 22848 56098
rect 22882 56096 22898 56098
rect 22882 56066 22920 56096
rect 23120 56066 23146 56096
rect 22882 56064 22898 56066
rect 22832 56048 22898 56064
rect 22832 55788 22898 55804
rect 22832 55754 22848 55788
rect 22882 55786 22898 55788
rect 22882 55756 22920 55786
rect 23120 55756 23146 55786
rect 22882 55754 22898 55756
rect 22832 55738 22898 55754
rect 23649 56098 23715 56114
rect 23649 56096 23665 56098
rect 23392 56066 23418 56096
rect 23618 56066 23665 56096
rect 23649 56064 23665 56066
rect 23699 56064 23715 56098
rect 23649 56048 23715 56064
rect 23649 55788 23715 55804
rect 23649 55786 23665 55788
rect 23392 55756 23418 55786
rect 23618 55756 23665 55786
rect 23649 55754 23665 55756
rect 23699 55754 23715 55788
rect 23649 55738 23715 55754
rect 27822 56098 27888 56114
rect 27822 56064 27838 56098
rect 27872 56096 27888 56098
rect 27872 56066 27910 56096
rect 28110 56066 28136 56096
rect 27872 56064 27888 56066
rect 27822 56048 27888 56064
rect 27822 55788 27888 55804
rect 27822 55754 27838 55788
rect 27872 55786 27888 55788
rect 27872 55756 27910 55786
rect 28110 55756 28136 55786
rect 27872 55754 27888 55756
rect 27822 55738 27888 55754
rect 28639 56098 28705 56114
rect 28639 56096 28655 56098
rect 28382 56066 28408 56096
rect 28608 56066 28655 56096
rect 28639 56064 28655 56066
rect 28689 56064 28705 56098
rect 28639 56048 28705 56064
rect 28639 55788 28705 55804
rect 28639 55786 28655 55788
rect 28382 55756 28408 55786
rect 28608 55756 28655 55786
rect 28639 55754 28655 55756
rect 28689 55754 28705 55788
rect 28639 55738 28705 55754
rect 32812 56098 32878 56114
rect 32812 56064 32828 56098
rect 32862 56096 32878 56098
rect 32862 56066 32900 56096
rect 33100 56066 33126 56096
rect 32862 56064 32878 56066
rect 32812 56048 32878 56064
rect 32812 55788 32878 55804
rect 32812 55754 32828 55788
rect 32862 55786 32878 55788
rect 32862 55756 32900 55786
rect 33100 55756 33126 55786
rect 32862 55754 32878 55756
rect 32812 55738 32878 55754
rect 33629 56098 33695 56114
rect 33629 56096 33645 56098
rect 33372 56066 33398 56096
rect 33598 56066 33645 56096
rect 33629 56064 33645 56066
rect 33679 56064 33695 56098
rect 33629 56048 33695 56064
rect 33629 55788 33695 55804
rect 33629 55786 33645 55788
rect 33372 55756 33398 55786
rect 33598 55756 33645 55786
rect 33629 55754 33645 55756
rect 33679 55754 33695 55788
rect 33629 55738 33695 55754
rect 37802 56098 37868 56114
rect 37802 56064 37818 56098
rect 37852 56096 37868 56098
rect 37852 56066 37890 56096
rect 38090 56066 38116 56096
rect 37852 56064 37868 56066
rect 37802 56048 37868 56064
rect 37802 55788 37868 55804
rect 37802 55754 37818 55788
rect 37852 55786 37868 55788
rect 37852 55756 37890 55786
rect 38090 55756 38116 55786
rect 37852 55754 37868 55756
rect 37802 55738 37868 55754
rect 38619 56098 38685 56114
rect 38619 56096 38635 56098
rect 38362 56066 38388 56096
rect 38588 56066 38635 56096
rect 38619 56064 38635 56066
rect 38669 56064 38685 56098
rect 38619 56048 38685 56064
rect 38619 55788 38685 55804
rect 38619 55786 38635 55788
rect 38362 55756 38388 55786
rect 38588 55756 38635 55786
rect 38619 55754 38635 55756
rect 38669 55754 38685 55788
rect 38619 55738 38685 55754
rect 42792 56098 42858 56114
rect 42792 56064 42808 56098
rect 42842 56096 42858 56098
rect 42842 56066 42880 56096
rect 43080 56066 43106 56096
rect 42842 56064 42858 56066
rect 42792 56048 42858 56064
rect 42792 55788 42858 55804
rect 42792 55754 42808 55788
rect 42842 55786 42858 55788
rect 42842 55756 42880 55786
rect 43080 55756 43106 55786
rect 42842 55754 42858 55756
rect 42792 55738 42858 55754
rect 43609 56098 43675 56114
rect 43609 56096 43625 56098
rect 43352 56066 43378 56096
rect 43578 56066 43625 56096
rect 43609 56064 43625 56066
rect 43659 56064 43675 56098
rect 43609 56048 43675 56064
rect 43609 55788 43675 55804
rect 43609 55786 43625 55788
rect 43352 55756 43378 55786
rect 43578 55756 43625 55786
rect 43609 55754 43625 55756
rect 43659 55754 43675 55788
rect 43609 55738 43675 55754
rect 47782 56098 47848 56114
rect 47782 56064 47798 56098
rect 47832 56096 47848 56098
rect 47832 56066 47870 56096
rect 48070 56066 48096 56096
rect 47832 56064 47848 56066
rect 47782 56048 47848 56064
rect 47782 55788 47848 55804
rect 47782 55754 47798 55788
rect 47832 55786 47848 55788
rect 47832 55756 47870 55786
rect 48070 55756 48096 55786
rect 47832 55754 47848 55756
rect 47782 55738 47848 55754
rect 48599 56098 48665 56114
rect 48599 56096 48615 56098
rect 48342 56066 48368 56096
rect 48568 56066 48615 56096
rect 48599 56064 48615 56066
rect 48649 56064 48665 56098
rect 48599 56048 48665 56064
rect 48599 55788 48665 55804
rect 48599 55786 48615 55788
rect 48342 55756 48368 55786
rect 48568 55756 48615 55786
rect 48599 55754 48615 55756
rect 48649 55754 48665 55788
rect 48599 55738 48665 55754
rect 52772 56098 52838 56114
rect 52772 56064 52788 56098
rect 52822 56096 52838 56098
rect 52822 56066 52860 56096
rect 53060 56066 53086 56096
rect 52822 56064 52838 56066
rect 52772 56048 52838 56064
rect 52772 55788 52838 55804
rect 52772 55754 52788 55788
rect 52822 55786 52838 55788
rect 52822 55756 52860 55786
rect 53060 55756 53086 55786
rect 52822 55754 52838 55756
rect 52772 55738 52838 55754
rect 53589 56098 53655 56114
rect 53589 56096 53605 56098
rect 53332 56066 53358 56096
rect 53558 56066 53605 56096
rect 53589 56064 53605 56066
rect 53639 56064 53655 56098
rect 53589 56048 53655 56064
rect 53589 55788 53655 55804
rect 53589 55786 53605 55788
rect 53332 55756 53358 55786
rect 53558 55756 53605 55786
rect 53589 55754 53605 55756
rect 53639 55754 53655 55788
rect 53589 55738 53655 55754
rect 57762 56098 57828 56114
rect 57762 56064 57778 56098
rect 57812 56096 57828 56098
rect 57812 56066 57850 56096
rect 58050 56066 58076 56096
rect 57812 56064 57828 56066
rect 57762 56048 57828 56064
rect 57762 55788 57828 55804
rect 57762 55754 57778 55788
rect 57812 55786 57828 55788
rect 57812 55756 57850 55786
rect 58050 55756 58076 55786
rect 57812 55754 57828 55756
rect 57762 55738 57828 55754
rect 58579 56098 58645 56114
rect 58579 56096 58595 56098
rect 58322 56066 58348 56096
rect 58548 56066 58595 56096
rect 58579 56064 58595 56066
rect 58629 56064 58645 56098
rect 58579 56048 58645 56064
rect 58579 55788 58645 55804
rect 58579 55786 58595 55788
rect 58322 55756 58348 55786
rect 58548 55756 58595 55786
rect 58579 55754 58595 55756
rect 58629 55754 58645 55788
rect 58579 55738 58645 55754
rect 62752 56098 62818 56114
rect 62752 56064 62768 56098
rect 62802 56096 62818 56098
rect 62802 56066 62840 56096
rect 63040 56066 63066 56096
rect 62802 56064 62818 56066
rect 62752 56048 62818 56064
rect 62752 55788 62818 55804
rect 62752 55754 62768 55788
rect 62802 55786 62818 55788
rect 62802 55756 62840 55786
rect 63040 55756 63066 55786
rect 62802 55754 62818 55756
rect 62752 55738 62818 55754
rect 63569 56098 63635 56114
rect 63569 56096 63585 56098
rect 63312 56066 63338 56096
rect 63538 56066 63585 56096
rect 63569 56064 63585 56066
rect 63619 56064 63635 56098
rect 63569 56048 63635 56064
rect 63569 55788 63635 55804
rect 63569 55786 63585 55788
rect 63312 55756 63338 55786
rect 63538 55756 63585 55786
rect 63569 55754 63585 55756
rect 63619 55754 63635 55788
rect 63569 55738 63635 55754
rect 67742 56098 67808 56114
rect 67742 56064 67758 56098
rect 67792 56096 67808 56098
rect 67792 56066 67830 56096
rect 68030 56066 68056 56096
rect 67792 56064 67808 56066
rect 67742 56048 67808 56064
rect 67742 55788 67808 55804
rect 67742 55754 67758 55788
rect 67792 55786 67808 55788
rect 67792 55756 67830 55786
rect 68030 55756 68056 55786
rect 67792 55754 67808 55756
rect 67742 55738 67808 55754
rect 68559 56098 68625 56114
rect 68559 56096 68575 56098
rect 68302 56066 68328 56096
rect 68528 56066 68575 56096
rect 68559 56064 68575 56066
rect 68609 56064 68625 56098
rect 68559 56048 68625 56064
rect 68559 55788 68625 55804
rect 68559 55786 68575 55788
rect 68302 55756 68328 55786
rect 68528 55756 68575 55786
rect 68559 55754 68575 55756
rect 68609 55754 68625 55788
rect 68559 55738 68625 55754
rect 72732 56098 72798 56114
rect 72732 56064 72748 56098
rect 72782 56096 72798 56098
rect 72782 56066 72820 56096
rect 73020 56066 73046 56096
rect 72782 56064 72798 56066
rect 72732 56048 72798 56064
rect 72732 55788 72798 55804
rect 72732 55754 72748 55788
rect 72782 55786 72798 55788
rect 72782 55756 72820 55786
rect 73020 55756 73046 55786
rect 72782 55754 72798 55756
rect 72732 55738 72798 55754
rect 73549 56098 73615 56114
rect 73549 56096 73565 56098
rect 73292 56066 73318 56096
rect 73518 56066 73565 56096
rect 73549 56064 73565 56066
rect 73599 56064 73615 56098
rect 73549 56048 73615 56064
rect 73549 55788 73615 55804
rect 73549 55786 73565 55788
rect 73292 55756 73318 55786
rect 73518 55756 73565 55786
rect 73549 55754 73565 55756
rect 73599 55754 73615 55788
rect 73549 55738 73615 55754
rect 77722 56098 77788 56114
rect 77722 56064 77738 56098
rect 77772 56096 77788 56098
rect 77772 56066 77810 56096
rect 78010 56066 78036 56096
rect 77772 56064 77788 56066
rect 77722 56048 77788 56064
rect 77722 55788 77788 55804
rect 77722 55754 77738 55788
rect 77772 55786 77788 55788
rect 77772 55756 77810 55786
rect 78010 55756 78036 55786
rect 77772 55754 77788 55756
rect 77722 55738 77788 55754
rect 78539 56098 78605 56114
rect 78539 56096 78555 56098
rect 78282 56066 78308 56096
rect 78508 56066 78555 56096
rect 78539 56064 78555 56066
rect 78589 56064 78605 56098
rect 78539 56048 78605 56064
rect 78539 55788 78605 55804
rect 78539 55786 78555 55788
rect 78282 55756 78308 55786
rect 78508 55756 78555 55786
rect 78539 55754 78555 55756
rect 78589 55754 78605 55788
rect 78539 55738 78605 55754
rect 2872 54388 2938 54404
rect 2872 54354 2888 54388
rect 2922 54386 2938 54388
rect 2922 54356 2960 54386
rect 3160 54356 3186 54386
rect 2922 54354 2938 54356
rect 2872 54338 2938 54354
rect 2872 54078 2938 54094
rect 2872 54044 2888 54078
rect 2922 54076 2938 54078
rect 2922 54046 2960 54076
rect 3160 54046 3186 54076
rect 2922 54044 2938 54046
rect 2872 54028 2938 54044
rect 3689 54388 3755 54404
rect 3689 54386 3705 54388
rect 3432 54356 3458 54386
rect 3658 54356 3705 54386
rect 3689 54354 3705 54356
rect 3739 54354 3755 54388
rect 3689 54338 3755 54354
rect 3689 54078 3755 54094
rect 3689 54076 3705 54078
rect 3432 54046 3458 54076
rect 3658 54046 3705 54076
rect 3689 54044 3705 54046
rect 3739 54044 3755 54078
rect 3689 54028 3755 54044
rect 7862 54388 7928 54404
rect 7862 54354 7878 54388
rect 7912 54386 7928 54388
rect 7912 54356 7950 54386
rect 8150 54356 8176 54386
rect 7912 54354 7928 54356
rect 7862 54338 7928 54354
rect 7862 54078 7928 54094
rect 7862 54044 7878 54078
rect 7912 54076 7928 54078
rect 7912 54046 7950 54076
rect 8150 54046 8176 54076
rect 7912 54044 7928 54046
rect 7862 54028 7928 54044
rect 8679 54388 8745 54404
rect 8679 54386 8695 54388
rect 8422 54356 8448 54386
rect 8648 54356 8695 54386
rect 8679 54354 8695 54356
rect 8729 54354 8745 54388
rect 8679 54338 8745 54354
rect 8679 54078 8745 54094
rect 8679 54076 8695 54078
rect 8422 54046 8448 54076
rect 8648 54046 8695 54076
rect 8679 54044 8695 54046
rect 8729 54044 8745 54078
rect 8679 54028 8745 54044
rect 12852 54388 12918 54404
rect 12852 54354 12868 54388
rect 12902 54386 12918 54388
rect 12902 54356 12940 54386
rect 13140 54356 13166 54386
rect 12902 54354 12918 54356
rect 12852 54338 12918 54354
rect 12852 54078 12918 54094
rect 12852 54044 12868 54078
rect 12902 54076 12918 54078
rect 12902 54046 12940 54076
rect 13140 54046 13166 54076
rect 12902 54044 12918 54046
rect 12852 54028 12918 54044
rect 13669 54388 13735 54404
rect 13669 54386 13685 54388
rect 13412 54356 13438 54386
rect 13638 54356 13685 54386
rect 13669 54354 13685 54356
rect 13719 54354 13735 54388
rect 13669 54338 13735 54354
rect 13669 54078 13735 54094
rect 13669 54076 13685 54078
rect 13412 54046 13438 54076
rect 13638 54046 13685 54076
rect 13669 54044 13685 54046
rect 13719 54044 13735 54078
rect 13669 54028 13735 54044
rect 17842 54388 17908 54404
rect 17842 54354 17858 54388
rect 17892 54386 17908 54388
rect 17892 54356 17930 54386
rect 18130 54356 18156 54386
rect 17892 54354 17908 54356
rect 17842 54338 17908 54354
rect 17842 54078 17908 54094
rect 17842 54044 17858 54078
rect 17892 54076 17908 54078
rect 17892 54046 17930 54076
rect 18130 54046 18156 54076
rect 17892 54044 17908 54046
rect 17842 54028 17908 54044
rect 18659 54388 18725 54404
rect 18659 54386 18675 54388
rect 18402 54356 18428 54386
rect 18628 54356 18675 54386
rect 18659 54354 18675 54356
rect 18709 54354 18725 54388
rect 18659 54338 18725 54354
rect 18659 54078 18725 54094
rect 18659 54076 18675 54078
rect 18402 54046 18428 54076
rect 18628 54046 18675 54076
rect 18659 54044 18675 54046
rect 18709 54044 18725 54078
rect 18659 54028 18725 54044
rect 22832 54388 22898 54404
rect 22832 54354 22848 54388
rect 22882 54386 22898 54388
rect 22882 54356 22920 54386
rect 23120 54356 23146 54386
rect 22882 54354 22898 54356
rect 22832 54338 22898 54354
rect 22832 54078 22898 54094
rect 22832 54044 22848 54078
rect 22882 54076 22898 54078
rect 22882 54046 22920 54076
rect 23120 54046 23146 54076
rect 22882 54044 22898 54046
rect 22832 54028 22898 54044
rect 23649 54388 23715 54404
rect 23649 54386 23665 54388
rect 23392 54356 23418 54386
rect 23618 54356 23665 54386
rect 23649 54354 23665 54356
rect 23699 54354 23715 54388
rect 23649 54338 23715 54354
rect 23649 54078 23715 54094
rect 23649 54076 23665 54078
rect 23392 54046 23418 54076
rect 23618 54046 23665 54076
rect 23649 54044 23665 54046
rect 23699 54044 23715 54078
rect 23649 54028 23715 54044
rect 27822 54388 27888 54404
rect 27822 54354 27838 54388
rect 27872 54386 27888 54388
rect 27872 54356 27910 54386
rect 28110 54356 28136 54386
rect 27872 54354 27888 54356
rect 27822 54338 27888 54354
rect 27822 54078 27888 54094
rect 27822 54044 27838 54078
rect 27872 54076 27888 54078
rect 27872 54046 27910 54076
rect 28110 54046 28136 54076
rect 27872 54044 27888 54046
rect 27822 54028 27888 54044
rect 28639 54388 28705 54404
rect 28639 54386 28655 54388
rect 28382 54356 28408 54386
rect 28608 54356 28655 54386
rect 28639 54354 28655 54356
rect 28689 54354 28705 54388
rect 28639 54338 28705 54354
rect 28639 54078 28705 54094
rect 28639 54076 28655 54078
rect 28382 54046 28408 54076
rect 28608 54046 28655 54076
rect 28639 54044 28655 54046
rect 28689 54044 28705 54078
rect 28639 54028 28705 54044
rect 32812 54388 32878 54404
rect 32812 54354 32828 54388
rect 32862 54386 32878 54388
rect 32862 54356 32900 54386
rect 33100 54356 33126 54386
rect 32862 54354 32878 54356
rect 32812 54338 32878 54354
rect 32812 54078 32878 54094
rect 32812 54044 32828 54078
rect 32862 54076 32878 54078
rect 32862 54046 32900 54076
rect 33100 54046 33126 54076
rect 32862 54044 32878 54046
rect 32812 54028 32878 54044
rect 33629 54388 33695 54404
rect 33629 54386 33645 54388
rect 33372 54356 33398 54386
rect 33598 54356 33645 54386
rect 33629 54354 33645 54356
rect 33679 54354 33695 54388
rect 33629 54338 33695 54354
rect 33629 54078 33695 54094
rect 33629 54076 33645 54078
rect 33372 54046 33398 54076
rect 33598 54046 33645 54076
rect 33629 54044 33645 54046
rect 33679 54044 33695 54078
rect 33629 54028 33695 54044
rect 37802 54388 37868 54404
rect 37802 54354 37818 54388
rect 37852 54386 37868 54388
rect 37852 54356 37890 54386
rect 38090 54356 38116 54386
rect 37852 54354 37868 54356
rect 37802 54338 37868 54354
rect 37802 54078 37868 54094
rect 37802 54044 37818 54078
rect 37852 54076 37868 54078
rect 37852 54046 37890 54076
rect 38090 54046 38116 54076
rect 37852 54044 37868 54046
rect 37802 54028 37868 54044
rect 38619 54388 38685 54404
rect 38619 54386 38635 54388
rect 38362 54356 38388 54386
rect 38588 54356 38635 54386
rect 38619 54354 38635 54356
rect 38669 54354 38685 54388
rect 38619 54338 38685 54354
rect 38619 54078 38685 54094
rect 38619 54076 38635 54078
rect 38362 54046 38388 54076
rect 38588 54046 38635 54076
rect 38619 54044 38635 54046
rect 38669 54044 38685 54078
rect 38619 54028 38685 54044
rect 42792 54388 42858 54404
rect 42792 54354 42808 54388
rect 42842 54386 42858 54388
rect 42842 54356 42880 54386
rect 43080 54356 43106 54386
rect 42842 54354 42858 54356
rect 42792 54338 42858 54354
rect 42792 54078 42858 54094
rect 42792 54044 42808 54078
rect 42842 54076 42858 54078
rect 42842 54046 42880 54076
rect 43080 54046 43106 54076
rect 42842 54044 42858 54046
rect 42792 54028 42858 54044
rect 43609 54388 43675 54404
rect 43609 54386 43625 54388
rect 43352 54356 43378 54386
rect 43578 54356 43625 54386
rect 43609 54354 43625 54356
rect 43659 54354 43675 54388
rect 43609 54338 43675 54354
rect 43609 54078 43675 54094
rect 43609 54076 43625 54078
rect 43352 54046 43378 54076
rect 43578 54046 43625 54076
rect 43609 54044 43625 54046
rect 43659 54044 43675 54078
rect 43609 54028 43675 54044
rect 47782 54388 47848 54404
rect 47782 54354 47798 54388
rect 47832 54386 47848 54388
rect 47832 54356 47870 54386
rect 48070 54356 48096 54386
rect 47832 54354 47848 54356
rect 47782 54338 47848 54354
rect 47782 54078 47848 54094
rect 47782 54044 47798 54078
rect 47832 54076 47848 54078
rect 47832 54046 47870 54076
rect 48070 54046 48096 54076
rect 47832 54044 47848 54046
rect 47782 54028 47848 54044
rect 48599 54388 48665 54404
rect 48599 54386 48615 54388
rect 48342 54356 48368 54386
rect 48568 54356 48615 54386
rect 48599 54354 48615 54356
rect 48649 54354 48665 54388
rect 48599 54338 48665 54354
rect 48599 54078 48665 54094
rect 48599 54076 48615 54078
rect 48342 54046 48368 54076
rect 48568 54046 48615 54076
rect 48599 54044 48615 54046
rect 48649 54044 48665 54078
rect 48599 54028 48665 54044
rect 52772 54388 52838 54404
rect 52772 54354 52788 54388
rect 52822 54386 52838 54388
rect 52822 54356 52860 54386
rect 53060 54356 53086 54386
rect 52822 54354 52838 54356
rect 52772 54338 52838 54354
rect 52772 54078 52838 54094
rect 52772 54044 52788 54078
rect 52822 54076 52838 54078
rect 52822 54046 52860 54076
rect 53060 54046 53086 54076
rect 52822 54044 52838 54046
rect 52772 54028 52838 54044
rect 53589 54388 53655 54404
rect 53589 54386 53605 54388
rect 53332 54356 53358 54386
rect 53558 54356 53605 54386
rect 53589 54354 53605 54356
rect 53639 54354 53655 54388
rect 53589 54338 53655 54354
rect 53589 54078 53655 54094
rect 53589 54076 53605 54078
rect 53332 54046 53358 54076
rect 53558 54046 53605 54076
rect 53589 54044 53605 54046
rect 53639 54044 53655 54078
rect 53589 54028 53655 54044
rect 57762 54388 57828 54404
rect 57762 54354 57778 54388
rect 57812 54386 57828 54388
rect 57812 54356 57850 54386
rect 58050 54356 58076 54386
rect 57812 54354 57828 54356
rect 57762 54338 57828 54354
rect 57762 54078 57828 54094
rect 57762 54044 57778 54078
rect 57812 54076 57828 54078
rect 57812 54046 57850 54076
rect 58050 54046 58076 54076
rect 57812 54044 57828 54046
rect 57762 54028 57828 54044
rect 58579 54388 58645 54404
rect 58579 54386 58595 54388
rect 58322 54356 58348 54386
rect 58548 54356 58595 54386
rect 58579 54354 58595 54356
rect 58629 54354 58645 54388
rect 58579 54338 58645 54354
rect 58579 54078 58645 54094
rect 58579 54076 58595 54078
rect 58322 54046 58348 54076
rect 58548 54046 58595 54076
rect 58579 54044 58595 54046
rect 58629 54044 58645 54078
rect 58579 54028 58645 54044
rect 62752 54388 62818 54404
rect 62752 54354 62768 54388
rect 62802 54386 62818 54388
rect 62802 54356 62840 54386
rect 63040 54356 63066 54386
rect 62802 54354 62818 54356
rect 62752 54338 62818 54354
rect 62752 54078 62818 54094
rect 62752 54044 62768 54078
rect 62802 54076 62818 54078
rect 62802 54046 62840 54076
rect 63040 54046 63066 54076
rect 62802 54044 62818 54046
rect 62752 54028 62818 54044
rect 63569 54388 63635 54404
rect 63569 54386 63585 54388
rect 63312 54356 63338 54386
rect 63538 54356 63585 54386
rect 63569 54354 63585 54356
rect 63619 54354 63635 54388
rect 63569 54338 63635 54354
rect 63569 54078 63635 54094
rect 63569 54076 63585 54078
rect 63312 54046 63338 54076
rect 63538 54046 63585 54076
rect 63569 54044 63585 54046
rect 63619 54044 63635 54078
rect 63569 54028 63635 54044
rect 67742 54388 67808 54404
rect 67742 54354 67758 54388
rect 67792 54386 67808 54388
rect 67792 54356 67830 54386
rect 68030 54356 68056 54386
rect 67792 54354 67808 54356
rect 67742 54338 67808 54354
rect 67742 54078 67808 54094
rect 67742 54044 67758 54078
rect 67792 54076 67808 54078
rect 67792 54046 67830 54076
rect 68030 54046 68056 54076
rect 67792 54044 67808 54046
rect 67742 54028 67808 54044
rect 68559 54388 68625 54404
rect 68559 54386 68575 54388
rect 68302 54356 68328 54386
rect 68528 54356 68575 54386
rect 68559 54354 68575 54356
rect 68609 54354 68625 54388
rect 68559 54338 68625 54354
rect 68559 54078 68625 54094
rect 68559 54076 68575 54078
rect 68302 54046 68328 54076
rect 68528 54046 68575 54076
rect 68559 54044 68575 54046
rect 68609 54044 68625 54078
rect 68559 54028 68625 54044
rect 72732 54388 72798 54404
rect 72732 54354 72748 54388
rect 72782 54386 72798 54388
rect 72782 54356 72820 54386
rect 73020 54356 73046 54386
rect 72782 54354 72798 54356
rect 72732 54338 72798 54354
rect 72732 54078 72798 54094
rect 72732 54044 72748 54078
rect 72782 54076 72798 54078
rect 72782 54046 72820 54076
rect 73020 54046 73046 54076
rect 72782 54044 72798 54046
rect 72732 54028 72798 54044
rect 73549 54388 73615 54404
rect 73549 54386 73565 54388
rect 73292 54356 73318 54386
rect 73518 54356 73565 54386
rect 73549 54354 73565 54356
rect 73599 54354 73615 54388
rect 73549 54338 73615 54354
rect 73549 54078 73615 54094
rect 73549 54076 73565 54078
rect 73292 54046 73318 54076
rect 73518 54046 73565 54076
rect 73549 54044 73565 54046
rect 73599 54044 73615 54078
rect 73549 54028 73615 54044
rect 77722 54388 77788 54404
rect 77722 54354 77738 54388
rect 77772 54386 77788 54388
rect 77772 54356 77810 54386
rect 78010 54356 78036 54386
rect 77772 54354 77788 54356
rect 77722 54338 77788 54354
rect 77722 54078 77788 54094
rect 77722 54044 77738 54078
rect 77772 54076 77788 54078
rect 77772 54046 77810 54076
rect 78010 54046 78036 54076
rect 77772 54044 77788 54046
rect 77722 54028 77788 54044
rect 78539 54388 78605 54404
rect 78539 54386 78555 54388
rect 78282 54356 78308 54386
rect 78508 54356 78555 54386
rect 78539 54354 78555 54356
rect 78589 54354 78605 54388
rect 78539 54338 78605 54354
rect 78539 54078 78605 54094
rect 78539 54076 78555 54078
rect 78282 54046 78308 54076
rect 78508 54046 78555 54076
rect 78539 54044 78555 54046
rect 78589 54044 78605 54078
rect 78539 54028 78605 54044
rect 2872 52678 2938 52694
rect 2872 52644 2888 52678
rect 2922 52676 2938 52678
rect 2922 52646 2960 52676
rect 3160 52646 3186 52676
rect 2922 52644 2938 52646
rect 2872 52628 2938 52644
rect 2872 52368 2938 52384
rect 2872 52334 2888 52368
rect 2922 52366 2938 52368
rect 2922 52336 2960 52366
rect 3160 52336 3186 52366
rect 2922 52334 2938 52336
rect 2872 52318 2938 52334
rect 3689 52678 3755 52694
rect 3689 52676 3705 52678
rect 3432 52646 3458 52676
rect 3658 52646 3705 52676
rect 3689 52644 3705 52646
rect 3739 52644 3755 52678
rect 3689 52628 3755 52644
rect 3689 52368 3755 52384
rect 3689 52366 3705 52368
rect 3432 52336 3458 52366
rect 3658 52336 3705 52366
rect 3689 52334 3705 52336
rect 3739 52334 3755 52368
rect 3689 52318 3755 52334
rect 7862 52678 7928 52694
rect 7862 52644 7878 52678
rect 7912 52676 7928 52678
rect 7912 52646 7950 52676
rect 8150 52646 8176 52676
rect 7912 52644 7928 52646
rect 7862 52628 7928 52644
rect 7862 52368 7928 52384
rect 7862 52334 7878 52368
rect 7912 52366 7928 52368
rect 7912 52336 7950 52366
rect 8150 52336 8176 52366
rect 7912 52334 7928 52336
rect 7862 52318 7928 52334
rect 8679 52678 8745 52694
rect 8679 52676 8695 52678
rect 8422 52646 8448 52676
rect 8648 52646 8695 52676
rect 8679 52644 8695 52646
rect 8729 52644 8745 52678
rect 8679 52628 8745 52644
rect 8679 52368 8745 52384
rect 8679 52366 8695 52368
rect 8422 52336 8448 52366
rect 8648 52336 8695 52366
rect 8679 52334 8695 52336
rect 8729 52334 8745 52368
rect 8679 52318 8745 52334
rect 12852 52678 12918 52694
rect 12852 52644 12868 52678
rect 12902 52676 12918 52678
rect 12902 52646 12940 52676
rect 13140 52646 13166 52676
rect 12902 52644 12918 52646
rect 12852 52628 12918 52644
rect 12852 52368 12918 52384
rect 12852 52334 12868 52368
rect 12902 52366 12918 52368
rect 12902 52336 12940 52366
rect 13140 52336 13166 52366
rect 12902 52334 12918 52336
rect 12852 52318 12918 52334
rect 13669 52678 13735 52694
rect 13669 52676 13685 52678
rect 13412 52646 13438 52676
rect 13638 52646 13685 52676
rect 13669 52644 13685 52646
rect 13719 52644 13735 52678
rect 13669 52628 13735 52644
rect 13669 52368 13735 52384
rect 13669 52366 13685 52368
rect 13412 52336 13438 52366
rect 13638 52336 13685 52366
rect 13669 52334 13685 52336
rect 13719 52334 13735 52368
rect 13669 52318 13735 52334
rect 17842 52678 17908 52694
rect 17842 52644 17858 52678
rect 17892 52676 17908 52678
rect 17892 52646 17930 52676
rect 18130 52646 18156 52676
rect 17892 52644 17908 52646
rect 17842 52628 17908 52644
rect 17842 52368 17908 52384
rect 17842 52334 17858 52368
rect 17892 52366 17908 52368
rect 17892 52336 17930 52366
rect 18130 52336 18156 52366
rect 17892 52334 17908 52336
rect 17842 52318 17908 52334
rect 18659 52678 18725 52694
rect 18659 52676 18675 52678
rect 18402 52646 18428 52676
rect 18628 52646 18675 52676
rect 18659 52644 18675 52646
rect 18709 52644 18725 52678
rect 18659 52628 18725 52644
rect 18659 52368 18725 52384
rect 18659 52366 18675 52368
rect 18402 52336 18428 52366
rect 18628 52336 18675 52366
rect 18659 52334 18675 52336
rect 18709 52334 18725 52368
rect 18659 52318 18725 52334
rect 22832 52678 22898 52694
rect 22832 52644 22848 52678
rect 22882 52676 22898 52678
rect 22882 52646 22920 52676
rect 23120 52646 23146 52676
rect 22882 52644 22898 52646
rect 22832 52628 22898 52644
rect 22832 52368 22898 52384
rect 22832 52334 22848 52368
rect 22882 52366 22898 52368
rect 22882 52336 22920 52366
rect 23120 52336 23146 52366
rect 22882 52334 22898 52336
rect 22832 52318 22898 52334
rect 23649 52678 23715 52694
rect 23649 52676 23665 52678
rect 23392 52646 23418 52676
rect 23618 52646 23665 52676
rect 23649 52644 23665 52646
rect 23699 52644 23715 52678
rect 23649 52628 23715 52644
rect 23649 52368 23715 52384
rect 23649 52366 23665 52368
rect 23392 52336 23418 52366
rect 23618 52336 23665 52366
rect 23649 52334 23665 52336
rect 23699 52334 23715 52368
rect 23649 52318 23715 52334
rect 27822 52678 27888 52694
rect 27822 52644 27838 52678
rect 27872 52676 27888 52678
rect 27872 52646 27910 52676
rect 28110 52646 28136 52676
rect 27872 52644 27888 52646
rect 27822 52628 27888 52644
rect 27822 52368 27888 52384
rect 27822 52334 27838 52368
rect 27872 52366 27888 52368
rect 27872 52336 27910 52366
rect 28110 52336 28136 52366
rect 27872 52334 27888 52336
rect 27822 52318 27888 52334
rect 28639 52678 28705 52694
rect 28639 52676 28655 52678
rect 28382 52646 28408 52676
rect 28608 52646 28655 52676
rect 28639 52644 28655 52646
rect 28689 52644 28705 52678
rect 28639 52628 28705 52644
rect 28639 52368 28705 52384
rect 28639 52366 28655 52368
rect 28382 52336 28408 52366
rect 28608 52336 28655 52366
rect 28639 52334 28655 52336
rect 28689 52334 28705 52368
rect 28639 52318 28705 52334
rect 32812 52678 32878 52694
rect 32812 52644 32828 52678
rect 32862 52676 32878 52678
rect 32862 52646 32900 52676
rect 33100 52646 33126 52676
rect 32862 52644 32878 52646
rect 32812 52628 32878 52644
rect 32812 52368 32878 52384
rect 32812 52334 32828 52368
rect 32862 52366 32878 52368
rect 32862 52336 32900 52366
rect 33100 52336 33126 52366
rect 32862 52334 32878 52336
rect 32812 52318 32878 52334
rect 33629 52678 33695 52694
rect 33629 52676 33645 52678
rect 33372 52646 33398 52676
rect 33598 52646 33645 52676
rect 33629 52644 33645 52646
rect 33679 52644 33695 52678
rect 33629 52628 33695 52644
rect 33629 52368 33695 52384
rect 33629 52366 33645 52368
rect 33372 52336 33398 52366
rect 33598 52336 33645 52366
rect 33629 52334 33645 52336
rect 33679 52334 33695 52368
rect 33629 52318 33695 52334
rect 37802 52678 37868 52694
rect 37802 52644 37818 52678
rect 37852 52676 37868 52678
rect 37852 52646 37890 52676
rect 38090 52646 38116 52676
rect 37852 52644 37868 52646
rect 37802 52628 37868 52644
rect 37802 52368 37868 52384
rect 37802 52334 37818 52368
rect 37852 52366 37868 52368
rect 37852 52336 37890 52366
rect 38090 52336 38116 52366
rect 37852 52334 37868 52336
rect 37802 52318 37868 52334
rect 38619 52678 38685 52694
rect 38619 52676 38635 52678
rect 38362 52646 38388 52676
rect 38588 52646 38635 52676
rect 38619 52644 38635 52646
rect 38669 52644 38685 52678
rect 38619 52628 38685 52644
rect 38619 52368 38685 52384
rect 38619 52366 38635 52368
rect 38362 52336 38388 52366
rect 38588 52336 38635 52366
rect 38619 52334 38635 52336
rect 38669 52334 38685 52368
rect 38619 52318 38685 52334
rect 42792 52678 42858 52694
rect 42792 52644 42808 52678
rect 42842 52676 42858 52678
rect 42842 52646 42880 52676
rect 43080 52646 43106 52676
rect 42842 52644 42858 52646
rect 42792 52628 42858 52644
rect 42792 52368 42858 52384
rect 42792 52334 42808 52368
rect 42842 52366 42858 52368
rect 42842 52336 42880 52366
rect 43080 52336 43106 52366
rect 42842 52334 42858 52336
rect 42792 52318 42858 52334
rect 43609 52678 43675 52694
rect 43609 52676 43625 52678
rect 43352 52646 43378 52676
rect 43578 52646 43625 52676
rect 43609 52644 43625 52646
rect 43659 52644 43675 52678
rect 43609 52628 43675 52644
rect 43609 52368 43675 52384
rect 43609 52366 43625 52368
rect 43352 52336 43378 52366
rect 43578 52336 43625 52366
rect 43609 52334 43625 52336
rect 43659 52334 43675 52368
rect 43609 52318 43675 52334
rect 47782 52678 47848 52694
rect 47782 52644 47798 52678
rect 47832 52676 47848 52678
rect 47832 52646 47870 52676
rect 48070 52646 48096 52676
rect 47832 52644 47848 52646
rect 47782 52628 47848 52644
rect 47782 52368 47848 52384
rect 47782 52334 47798 52368
rect 47832 52366 47848 52368
rect 47832 52336 47870 52366
rect 48070 52336 48096 52366
rect 47832 52334 47848 52336
rect 47782 52318 47848 52334
rect 48599 52678 48665 52694
rect 48599 52676 48615 52678
rect 48342 52646 48368 52676
rect 48568 52646 48615 52676
rect 48599 52644 48615 52646
rect 48649 52644 48665 52678
rect 48599 52628 48665 52644
rect 48599 52368 48665 52384
rect 48599 52366 48615 52368
rect 48342 52336 48368 52366
rect 48568 52336 48615 52366
rect 48599 52334 48615 52336
rect 48649 52334 48665 52368
rect 48599 52318 48665 52334
rect 52772 52678 52838 52694
rect 52772 52644 52788 52678
rect 52822 52676 52838 52678
rect 52822 52646 52860 52676
rect 53060 52646 53086 52676
rect 52822 52644 52838 52646
rect 52772 52628 52838 52644
rect 52772 52368 52838 52384
rect 52772 52334 52788 52368
rect 52822 52366 52838 52368
rect 52822 52336 52860 52366
rect 53060 52336 53086 52366
rect 52822 52334 52838 52336
rect 52772 52318 52838 52334
rect 53589 52678 53655 52694
rect 53589 52676 53605 52678
rect 53332 52646 53358 52676
rect 53558 52646 53605 52676
rect 53589 52644 53605 52646
rect 53639 52644 53655 52678
rect 53589 52628 53655 52644
rect 53589 52368 53655 52384
rect 53589 52366 53605 52368
rect 53332 52336 53358 52366
rect 53558 52336 53605 52366
rect 53589 52334 53605 52336
rect 53639 52334 53655 52368
rect 53589 52318 53655 52334
rect 57762 52678 57828 52694
rect 57762 52644 57778 52678
rect 57812 52676 57828 52678
rect 57812 52646 57850 52676
rect 58050 52646 58076 52676
rect 57812 52644 57828 52646
rect 57762 52628 57828 52644
rect 57762 52368 57828 52384
rect 57762 52334 57778 52368
rect 57812 52366 57828 52368
rect 57812 52336 57850 52366
rect 58050 52336 58076 52366
rect 57812 52334 57828 52336
rect 57762 52318 57828 52334
rect 58579 52678 58645 52694
rect 58579 52676 58595 52678
rect 58322 52646 58348 52676
rect 58548 52646 58595 52676
rect 58579 52644 58595 52646
rect 58629 52644 58645 52678
rect 58579 52628 58645 52644
rect 58579 52368 58645 52384
rect 58579 52366 58595 52368
rect 58322 52336 58348 52366
rect 58548 52336 58595 52366
rect 58579 52334 58595 52336
rect 58629 52334 58645 52368
rect 58579 52318 58645 52334
rect 62752 52678 62818 52694
rect 62752 52644 62768 52678
rect 62802 52676 62818 52678
rect 62802 52646 62840 52676
rect 63040 52646 63066 52676
rect 62802 52644 62818 52646
rect 62752 52628 62818 52644
rect 62752 52368 62818 52384
rect 62752 52334 62768 52368
rect 62802 52366 62818 52368
rect 62802 52336 62840 52366
rect 63040 52336 63066 52366
rect 62802 52334 62818 52336
rect 62752 52318 62818 52334
rect 63569 52678 63635 52694
rect 63569 52676 63585 52678
rect 63312 52646 63338 52676
rect 63538 52646 63585 52676
rect 63569 52644 63585 52646
rect 63619 52644 63635 52678
rect 63569 52628 63635 52644
rect 63569 52368 63635 52384
rect 63569 52366 63585 52368
rect 63312 52336 63338 52366
rect 63538 52336 63585 52366
rect 63569 52334 63585 52336
rect 63619 52334 63635 52368
rect 63569 52318 63635 52334
rect 67742 52678 67808 52694
rect 67742 52644 67758 52678
rect 67792 52676 67808 52678
rect 67792 52646 67830 52676
rect 68030 52646 68056 52676
rect 67792 52644 67808 52646
rect 67742 52628 67808 52644
rect 67742 52368 67808 52384
rect 67742 52334 67758 52368
rect 67792 52366 67808 52368
rect 67792 52336 67830 52366
rect 68030 52336 68056 52366
rect 67792 52334 67808 52336
rect 67742 52318 67808 52334
rect 68559 52678 68625 52694
rect 68559 52676 68575 52678
rect 68302 52646 68328 52676
rect 68528 52646 68575 52676
rect 68559 52644 68575 52646
rect 68609 52644 68625 52678
rect 68559 52628 68625 52644
rect 68559 52368 68625 52384
rect 68559 52366 68575 52368
rect 68302 52336 68328 52366
rect 68528 52336 68575 52366
rect 68559 52334 68575 52336
rect 68609 52334 68625 52368
rect 68559 52318 68625 52334
rect 72732 52678 72798 52694
rect 72732 52644 72748 52678
rect 72782 52676 72798 52678
rect 72782 52646 72820 52676
rect 73020 52646 73046 52676
rect 72782 52644 72798 52646
rect 72732 52628 72798 52644
rect 72732 52368 72798 52384
rect 72732 52334 72748 52368
rect 72782 52366 72798 52368
rect 72782 52336 72820 52366
rect 73020 52336 73046 52366
rect 72782 52334 72798 52336
rect 72732 52318 72798 52334
rect 73549 52678 73615 52694
rect 73549 52676 73565 52678
rect 73292 52646 73318 52676
rect 73518 52646 73565 52676
rect 73549 52644 73565 52646
rect 73599 52644 73615 52678
rect 73549 52628 73615 52644
rect 73549 52368 73615 52384
rect 73549 52366 73565 52368
rect 73292 52336 73318 52366
rect 73518 52336 73565 52366
rect 73549 52334 73565 52336
rect 73599 52334 73615 52368
rect 73549 52318 73615 52334
rect 77722 52678 77788 52694
rect 77722 52644 77738 52678
rect 77772 52676 77788 52678
rect 77772 52646 77810 52676
rect 78010 52646 78036 52676
rect 77772 52644 77788 52646
rect 77722 52628 77788 52644
rect 77722 52368 77788 52384
rect 77722 52334 77738 52368
rect 77772 52366 77788 52368
rect 77772 52336 77810 52366
rect 78010 52336 78036 52366
rect 77772 52334 77788 52336
rect 77722 52318 77788 52334
rect 78539 52678 78605 52694
rect 78539 52676 78555 52678
rect 78282 52646 78308 52676
rect 78508 52646 78555 52676
rect 78539 52644 78555 52646
rect 78589 52644 78605 52678
rect 78539 52628 78605 52644
rect 78539 52368 78605 52384
rect 78539 52366 78555 52368
rect 78282 52336 78308 52366
rect 78508 52336 78555 52366
rect 78539 52334 78555 52336
rect 78589 52334 78605 52368
rect 78539 52318 78605 52334
rect 2872 50968 2938 50984
rect 2872 50934 2888 50968
rect 2922 50966 2938 50968
rect 2922 50936 2960 50966
rect 3160 50936 3186 50966
rect 2922 50934 2938 50936
rect 2872 50918 2938 50934
rect 2872 50658 2938 50674
rect 2872 50624 2888 50658
rect 2922 50656 2938 50658
rect 2922 50626 2960 50656
rect 3160 50626 3186 50656
rect 2922 50624 2938 50626
rect 2872 50608 2938 50624
rect 3689 50968 3755 50984
rect 3689 50966 3705 50968
rect 3432 50936 3458 50966
rect 3658 50936 3705 50966
rect 3689 50934 3705 50936
rect 3739 50934 3755 50968
rect 3689 50918 3755 50934
rect 3689 50658 3755 50674
rect 3689 50656 3705 50658
rect 3432 50626 3458 50656
rect 3658 50626 3705 50656
rect 3689 50624 3705 50626
rect 3739 50624 3755 50658
rect 3689 50608 3755 50624
rect 7862 50968 7928 50984
rect 7862 50934 7878 50968
rect 7912 50966 7928 50968
rect 7912 50936 7950 50966
rect 8150 50936 8176 50966
rect 7912 50934 7928 50936
rect 7862 50918 7928 50934
rect 7862 50658 7928 50674
rect 7862 50624 7878 50658
rect 7912 50656 7928 50658
rect 7912 50626 7950 50656
rect 8150 50626 8176 50656
rect 7912 50624 7928 50626
rect 7862 50608 7928 50624
rect 8679 50968 8745 50984
rect 8679 50966 8695 50968
rect 8422 50936 8448 50966
rect 8648 50936 8695 50966
rect 8679 50934 8695 50936
rect 8729 50934 8745 50968
rect 8679 50918 8745 50934
rect 8679 50658 8745 50674
rect 8679 50656 8695 50658
rect 8422 50626 8448 50656
rect 8648 50626 8695 50656
rect 8679 50624 8695 50626
rect 8729 50624 8745 50658
rect 8679 50608 8745 50624
rect 12852 50968 12918 50984
rect 12852 50934 12868 50968
rect 12902 50966 12918 50968
rect 12902 50936 12940 50966
rect 13140 50936 13166 50966
rect 12902 50934 12918 50936
rect 12852 50918 12918 50934
rect 12852 50658 12918 50674
rect 12852 50624 12868 50658
rect 12902 50656 12918 50658
rect 12902 50626 12940 50656
rect 13140 50626 13166 50656
rect 12902 50624 12918 50626
rect 12852 50608 12918 50624
rect 13669 50968 13735 50984
rect 13669 50966 13685 50968
rect 13412 50936 13438 50966
rect 13638 50936 13685 50966
rect 13669 50934 13685 50936
rect 13719 50934 13735 50968
rect 13669 50918 13735 50934
rect 13669 50658 13735 50674
rect 13669 50656 13685 50658
rect 13412 50626 13438 50656
rect 13638 50626 13685 50656
rect 13669 50624 13685 50626
rect 13719 50624 13735 50658
rect 13669 50608 13735 50624
rect 17842 50968 17908 50984
rect 17842 50934 17858 50968
rect 17892 50966 17908 50968
rect 17892 50936 17930 50966
rect 18130 50936 18156 50966
rect 17892 50934 17908 50936
rect 17842 50918 17908 50934
rect 17842 50658 17908 50674
rect 17842 50624 17858 50658
rect 17892 50656 17908 50658
rect 17892 50626 17930 50656
rect 18130 50626 18156 50656
rect 17892 50624 17908 50626
rect 17842 50608 17908 50624
rect 18659 50968 18725 50984
rect 18659 50966 18675 50968
rect 18402 50936 18428 50966
rect 18628 50936 18675 50966
rect 18659 50934 18675 50936
rect 18709 50934 18725 50968
rect 18659 50918 18725 50934
rect 18659 50658 18725 50674
rect 18659 50656 18675 50658
rect 18402 50626 18428 50656
rect 18628 50626 18675 50656
rect 18659 50624 18675 50626
rect 18709 50624 18725 50658
rect 18659 50608 18725 50624
rect 22832 50968 22898 50984
rect 22832 50934 22848 50968
rect 22882 50966 22898 50968
rect 22882 50936 22920 50966
rect 23120 50936 23146 50966
rect 22882 50934 22898 50936
rect 22832 50918 22898 50934
rect 22832 50658 22898 50674
rect 22832 50624 22848 50658
rect 22882 50656 22898 50658
rect 22882 50626 22920 50656
rect 23120 50626 23146 50656
rect 22882 50624 22898 50626
rect 22832 50608 22898 50624
rect 23649 50968 23715 50984
rect 23649 50966 23665 50968
rect 23392 50936 23418 50966
rect 23618 50936 23665 50966
rect 23649 50934 23665 50936
rect 23699 50934 23715 50968
rect 23649 50918 23715 50934
rect 23649 50658 23715 50674
rect 23649 50656 23665 50658
rect 23392 50626 23418 50656
rect 23618 50626 23665 50656
rect 23649 50624 23665 50626
rect 23699 50624 23715 50658
rect 23649 50608 23715 50624
rect 27822 50968 27888 50984
rect 27822 50934 27838 50968
rect 27872 50966 27888 50968
rect 27872 50936 27910 50966
rect 28110 50936 28136 50966
rect 27872 50934 27888 50936
rect 27822 50918 27888 50934
rect 27822 50658 27888 50674
rect 27822 50624 27838 50658
rect 27872 50656 27888 50658
rect 27872 50626 27910 50656
rect 28110 50626 28136 50656
rect 27872 50624 27888 50626
rect 27822 50608 27888 50624
rect 28639 50968 28705 50984
rect 28639 50966 28655 50968
rect 28382 50936 28408 50966
rect 28608 50936 28655 50966
rect 28639 50934 28655 50936
rect 28689 50934 28705 50968
rect 28639 50918 28705 50934
rect 28639 50658 28705 50674
rect 28639 50656 28655 50658
rect 28382 50626 28408 50656
rect 28608 50626 28655 50656
rect 28639 50624 28655 50626
rect 28689 50624 28705 50658
rect 28639 50608 28705 50624
rect 32812 50968 32878 50984
rect 32812 50934 32828 50968
rect 32862 50966 32878 50968
rect 32862 50936 32900 50966
rect 33100 50936 33126 50966
rect 32862 50934 32878 50936
rect 32812 50918 32878 50934
rect 32812 50658 32878 50674
rect 32812 50624 32828 50658
rect 32862 50656 32878 50658
rect 32862 50626 32900 50656
rect 33100 50626 33126 50656
rect 32862 50624 32878 50626
rect 32812 50608 32878 50624
rect 33629 50968 33695 50984
rect 33629 50966 33645 50968
rect 33372 50936 33398 50966
rect 33598 50936 33645 50966
rect 33629 50934 33645 50936
rect 33679 50934 33695 50968
rect 33629 50918 33695 50934
rect 33629 50658 33695 50674
rect 33629 50656 33645 50658
rect 33372 50626 33398 50656
rect 33598 50626 33645 50656
rect 33629 50624 33645 50626
rect 33679 50624 33695 50658
rect 33629 50608 33695 50624
rect 37802 50968 37868 50984
rect 37802 50934 37818 50968
rect 37852 50966 37868 50968
rect 37852 50936 37890 50966
rect 38090 50936 38116 50966
rect 37852 50934 37868 50936
rect 37802 50918 37868 50934
rect 37802 50658 37868 50674
rect 37802 50624 37818 50658
rect 37852 50656 37868 50658
rect 37852 50626 37890 50656
rect 38090 50626 38116 50656
rect 37852 50624 37868 50626
rect 37802 50608 37868 50624
rect 38619 50968 38685 50984
rect 38619 50966 38635 50968
rect 38362 50936 38388 50966
rect 38588 50936 38635 50966
rect 38619 50934 38635 50936
rect 38669 50934 38685 50968
rect 38619 50918 38685 50934
rect 38619 50658 38685 50674
rect 38619 50656 38635 50658
rect 38362 50626 38388 50656
rect 38588 50626 38635 50656
rect 38619 50624 38635 50626
rect 38669 50624 38685 50658
rect 38619 50608 38685 50624
rect 42792 50968 42858 50984
rect 42792 50934 42808 50968
rect 42842 50966 42858 50968
rect 42842 50936 42880 50966
rect 43080 50936 43106 50966
rect 42842 50934 42858 50936
rect 42792 50918 42858 50934
rect 42792 50658 42858 50674
rect 42792 50624 42808 50658
rect 42842 50656 42858 50658
rect 42842 50626 42880 50656
rect 43080 50626 43106 50656
rect 42842 50624 42858 50626
rect 42792 50608 42858 50624
rect 43609 50968 43675 50984
rect 43609 50966 43625 50968
rect 43352 50936 43378 50966
rect 43578 50936 43625 50966
rect 43609 50934 43625 50936
rect 43659 50934 43675 50968
rect 43609 50918 43675 50934
rect 43609 50658 43675 50674
rect 43609 50656 43625 50658
rect 43352 50626 43378 50656
rect 43578 50626 43625 50656
rect 43609 50624 43625 50626
rect 43659 50624 43675 50658
rect 43609 50608 43675 50624
rect 47782 50968 47848 50984
rect 47782 50934 47798 50968
rect 47832 50966 47848 50968
rect 47832 50936 47870 50966
rect 48070 50936 48096 50966
rect 47832 50934 47848 50936
rect 47782 50918 47848 50934
rect 47782 50658 47848 50674
rect 47782 50624 47798 50658
rect 47832 50656 47848 50658
rect 47832 50626 47870 50656
rect 48070 50626 48096 50656
rect 47832 50624 47848 50626
rect 47782 50608 47848 50624
rect 48599 50968 48665 50984
rect 48599 50966 48615 50968
rect 48342 50936 48368 50966
rect 48568 50936 48615 50966
rect 48599 50934 48615 50936
rect 48649 50934 48665 50968
rect 48599 50918 48665 50934
rect 48599 50658 48665 50674
rect 48599 50656 48615 50658
rect 48342 50626 48368 50656
rect 48568 50626 48615 50656
rect 48599 50624 48615 50626
rect 48649 50624 48665 50658
rect 48599 50608 48665 50624
rect 52772 50968 52838 50984
rect 52772 50934 52788 50968
rect 52822 50966 52838 50968
rect 52822 50936 52860 50966
rect 53060 50936 53086 50966
rect 52822 50934 52838 50936
rect 52772 50918 52838 50934
rect 52772 50658 52838 50674
rect 52772 50624 52788 50658
rect 52822 50656 52838 50658
rect 52822 50626 52860 50656
rect 53060 50626 53086 50656
rect 52822 50624 52838 50626
rect 52772 50608 52838 50624
rect 53589 50968 53655 50984
rect 53589 50966 53605 50968
rect 53332 50936 53358 50966
rect 53558 50936 53605 50966
rect 53589 50934 53605 50936
rect 53639 50934 53655 50968
rect 53589 50918 53655 50934
rect 53589 50658 53655 50674
rect 53589 50656 53605 50658
rect 53332 50626 53358 50656
rect 53558 50626 53605 50656
rect 53589 50624 53605 50626
rect 53639 50624 53655 50658
rect 53589 50608 53655 50624
rect 57762 50968 57828 50984
rect 57762 50934 57778 50968
rect 57812 50966 57828 50968
rect 57812 50936 57850 50966
rect 58050 50936 58076 50966
rect 57812 50934 57828 50936
rect 57762 50918 57828 50934
rect 57762 50658 57828 50674
rect 57762 50624 57778 50658
rect 57812 50656 57828 50658
rect 57812 50626 57850 50656
rect 58050 50626 58076 50656
rect 57812 50624 57828 50626
rect 57762 50608 57828 50624
rect 58579 50968 58645 50984
rect 58579 50966 58595 50968
rect 58322 50936 58348 50966
rect 58548 50936 58595 50966
rect 58579 50934 58595 50936
rect 58629 50934 58645 50968
rect 58579 50918 58645 50934
rect 58579 50658 58645 50674
rect 58579 50656 58595 50658
rect 58322 50626 58348 50656
rect 58548 50626 58595 50656
rect 58579 50624 58595 50626
rect 58629 50624 58645 50658
rect 58579 50608 58645 50624
rect 62752 50968 62818 50984
rect 62752 50934 62768 50968
rect 62802 50966 62818 50968
rect 62802 50936 62840 50966
rect 63040 50936 63066 50966
rect 62802 50934 62818 50936
rect 62752 50918 62818 50934
rect 62752 50658 62818 50674
rect 62752 50624 62768 50658
rect 62802 50656 62818 50658
rect 62802 50626 62840 50656
rect 63040 50626 63066 50656
rect 62802 50624 62818 50626
rect 62752 50608 62818 50624
rect 63569 50968 63635 50984
rect 63569 50966 63585 50968
rect 63312 50936 63338 50966
rect 63538 50936 63585 50966
rect 63569 50934 63585 50936
rect 63619 50934 63635 50968
rect 63569 50918 63635 50934
rect 63569 50658 63635 50674
rect 63569 50656 63585 50658
rect 63312 50626 63338 50656
rect 63538 50626 63585 50656
rect 63569 50624 63585 50626
rect 63619 50624 63635 50658
rect 63569 50608 63635 50624
rect 67742 50968 67808 50984
rect 67742 50934 67758 50968
rect 67792 50966 67808 50968
rect 67792 50936 67830 50966
rect 68030 50936 68056 50966
rect 67792 50934 67808 50936
rect 67742 50918 67808 50934
rect 67742 50658 67808 50674
rect 67742 50624 67758 50658
rect 67792 50656 67808 50658
rect 67792 50626 67830 50656
rect 68030 50626 68056 50656
rect 67792 50624 67808 50626
rect 67742 50608 67808 50624
rect 68559 50968 68625 50984
rect 68559 50966 68575 50968
rect 68302 50936 68328 50966
rect 68528 50936 68575 50966
rect 68559 50934 68575 50936
rect 68609 50934 68625 50968
rect 68559 50918 68625 50934
rect 68559 50658 68625 50674
rect 68559 50656 68575 50658
rect 68302 50626 68328 50656
rect 68528 50626 68575 50656
rect 68559 50624 68575 50626
rect 68609 50624 68625 50658
rect 68559 50608 68625 50624
rect 72732 50968 72798 50984
rect 72732 50934 72748 50968
rect 72782 50966 72798 50968
rect 72782 50936 72820 50966
rect 73020 50936 73046 50966
rect 72782 50934 72798 50936
rect 72732 50918 72798 50934
rect 72732 50658 72798 50674
rect 72732 50624 72748 50658
rect 72782 50656 72798 50658
rect 72782 50626 72820 50656
rect 73020 50626 73046 50656
rect 72782 50624 72798 50626
rect 72732 50608 72798 50624
rect 73549 50968 73615 50984
rect 73549 50966 73565 50968
rect 73292 50936 73318 50966
rect 73518 50936 73565 50966
rect 73549 50934 73565 50936
rect 73599 50934 73615 50968
rect 73549 50918 73615 50934
rect 73549 50658 73615 50674
rect 73549 50656 73565 50658
rect 73292 50626 73318 50656
rect 73518 50626 73565 50656
rect 73549 50624 73565 50626
rect 73599 50624 73615 50658
rect 73549 50608 73615 50624
rect 77722 50968 77788 50984
rect 77722 50934 77738 50968
rect 77772 50966 77788 50968
rect 77772 50936 77810 50966
rect 78010 50936 78036 50966
rect 77772 50934 77788 50936
rect 77722 50918 77788 50934
rect 77722 50658 77788 50674
rect 77722 50624 77738 50658
rect 77772 50656 77788 50658
rect 77772 50626 77810 50656
rect 78010 50626 78036 50656
rect 77772 50624 77788 50626
rect 77722 50608 77788 50624
rect 78539 50968 78605 50984
rect 78539 50966 78555 50968
rect 78282 50936 78308 50966
rect 78508 50936 78555 50966
rect 78539 50934 78555 50936
rect 78589 50934 78605 50968
rect 78539 50918 78605 50934
rect 78539 50658 78605 50674
rect 78539 50656 78555 50658
rect 78282 50626 78308 50656
rect 78508 50626 78555 50656
rect 78539 50624 78555 50626
rect 78589 50624 78605 50658
rect 78539 50608 78605 50624
rect 2872 49258 2938 49274
rect 2872 49224 2888 49258
rect 2922 49256 2938 49258
rect 2922 49226 2960 49256
rect 3160 49226 3186 49256
rect 2922 49224 2938 49226
rect 2872 49208 2938 49224
rect 2872 48948 2938 48964
rect 2872 48914 2888 48948
rect 2922 48946 2938 48948
rect 2922 48916 2960 48946
rect 3160 48916 3186 48946
rect 2922 48914 2938 48916
rect 2872 48898 2938 48914
rect 3689 49258 3755 49274
rect 3689 49256 3705 49258
rect 3432 49226 3458 49256
rect 3658 49226 3705 49256
rect 3689 49224 3705 49226
rect 3739 49224 3755 49258
rect 3689 49208 3755 49224
rect 3689 48948 3755 48964
rect 3689 48946 3705 48948
rect 3432 48916 3458 48946
rect 3658 48916 3705 48946
rect 3689 48914 3705 48916
rect 3739 48914 3755 48948
rect 3689 48898 3755 48914
rect 7862 49258 7928 49274
rect 7862 49224 7878 49258
rect 7912 49256 7928 49258
rect 7912 49226 7950 49256
rect 8150 49226 8176 49256
rect 7912 49224 7928 49226
rect 7862 49208 7928 49224
rect 7862 48948 7928 48964
rect 7862 48914 7878 48948
rect 7912 48946 7928 48948
rect 7912 48916 7950 48946
rect 8150 48916 8176 48946
rect 7912 48914 7928 48916
rect 7862 48898 7928 48914
rect 8679 49258 8745 49274
rect 8679 49256 8695 49258
rect 8422 49226 8448 49256
rect 8648 49226 8695 49256
rect 8679 49224 8695 49226
rect 8729 49224 8745 49258
rect 8679 49208 8745 49224
rect 8679 48948 8745 48964
rect 8679 48946 8695 48948
rect 8422 48916 8448 48946
rect 8648 48916 8695 48946
rect 8679 48914 8695 48916
rect 8729 48914 8745 48948
rect 8679 48898 8745 48914
rect 12852 49258 12918 49274
rect 12852 49224 12868 49258
rect 12902 49256 12918 49258
rect 12902 49226 12940 49256
rect 13140 49226 13166 49256
rect 12902 49224 12918 49226
rect 12852 49208 12918 49224
rect 12852 48948 12918 48964
rect 12852 48914 12868 48948
rect 12902 48946 12918 48948
rect 12902 48916 12940 48946
rect 13140 48916 13166 48946
rect 12902 48914 12918 48916
rect 12852 48898 12918 48914
rect 13669 49258 13735 49274
rect 13669 49256 13685 49258
rect 13412 49226 13438 49256
rect 13638 49226 13685 49256
rect 13669 49224 13685 49226
rect 13719 49224 13735 49258
rect 13669 49208 13735 49224
rect 13669 48948 13735 48964
rect 13669 48946 13685 48948
rect 13412 48916 13438 48946
rect 13638 48916 13685 48946
rect 13669 48914 13685 48916
rect 13719 48914 13735 48948
rect 13669 48898 13735 48914
rect 17842 49258 17908 49274
rect 17842 49224 17858 49258
rect 17892 49256 17908 49258
rect 17892 49226 17930 49256
rect 18130 49226 18156 49256
rect 17892 49224 17908 49226
rect 17842 49208 17908 49224
rect 17842 48948 17908 48964
rect 17842 48914 17858 48948
rect 17892 48946 17908 48948
rect 17892 48916 17930 48946
rect 18130 48916 18156 48946
rect 17892 48914 17908 48916
rect 17842 48898 17908 48914
rect 18659 49258 18725 49274
rect 18659 49256 18675 49258
rect 18402 49226 18428 49256
rect 18628 49226 18675 49256
rect 18659 49224 18675 49226
rect 18709 49224 18725 49258
rect 18659 49208 18725 49224
rect 18659 48948 18725 48964
rect 18659 48946 18675 48948
rect 18402 48916 18428 48946
rect 18628 48916 18675 48946
rect 18659 48914 18675 48916
rect 18709 48914 18725 48948
rect 18659 48898 18725 48914
rect 22832 49258 22898 49274
rect 22832 49224 22848 49258
rect 22882 49256 22898 49258
rect 22882 49226 22920 49256
rect 23120 49226 23146 49256
rect 22882 49224 22898 49226
rect 22832 49208 22898 49224
rect 22832 48948 22898 48964
rect 22832 48914 22848 48948
rect 22882 48946 22898 48948
rect 22882 48916 22920 48946
rect 23120 48916 23146 48946
rect 22882 48914 22898 48916
rect 22832 48898 22898 48914
rect 23649 49258 23715 49274
rect 23649 49256 23665 49258
rect 23392 49226 23418 49256
rect 23618 49226 23665 49256
rect 23649 49224 23665 49226
rect 23699 49224 23715 49258
rect 23649 49208 23715 49224
rect 23649 48948 23715 48964
rect 23649 48946 23665 48948
rect 23392 48916 23418 48946
rect 23618 48916 23665 48946
rect 23649 48914 23665 48916
rect 23699 48914 23715 48948
rect 23649 48898 23715 48914
rect 27822 49258 27888 49274
rect 27822 49224 27838 49258
rect 27872 49256 27888 49258
rect 27872 49226 27910 49256
rect 28110 49226 28136 49256
rect 27872 49224 27888 49226
rect 27822 49208 27888 49224
rect 27822 48948 27888 48964
rect 27822 48914 27838 48948
rect 27872 48946 27888 48948
rect 27872 48916 27910 48946
rect 28110 48916 28136 48946
rect 27872 48914 27888 48916
rect 27822 48898 27888 48914
rect 28639 49258 28705 49274
rect 28639 49256 28655 49258
rect 28382 49226 28408 49256
rect 28608 49226 28655 49256
rect 28639 49224 28655 49226
rect 28689 49224 28705 49258
rect 28639 49208 28705 49224
rect 28639 48948 28705 48964
rect 28639 48946 28655 48948
rect 28382 48916 28408 48946
rect 28608 48916 28655 48946
rect 28639 48914 28655 48916
rect 28689 48914 28705 48948
rect 28639 48898 28705 48914
rect 32812 49258 32878 49274
rect 32812 49224 32828 49258
rect 32862 49256 32878 49258
rect 32862 49226 32900 49256
rect 33100 49226 33126 49256
rect 32862 49224 32878 49226
rect 32812 49208 32878 49224
rect 32812 48948 32878 48964
rect 32812 48914 32828 48948
rect 32862 48946 32878 48948
rect 32862 48916 32900 48946
rect 33100 48916 33126 48946
rect 32862 48914 32878 48916
rect 32812 48898 32878 48914
rect 33629 49258 33695 49274
rect 33629 49256 33645 49258
rect 33372 49226 33398 49256
rect 33598 49226 33645 49256
rect 33629 49224 33645 49226
rect 33679 49224 33695 49258
rect 33629 49208 33695 49224
rect 33629 48948 33695 48964
rect 33629 48946 33645 48948
rect 33372 48916 33398 48946
rect 33598 48916 33645 48946
rect 33629 48914 33645 48916
rect 33679 48914 33695 48948
rect 33629 48898 33695 48914
rect 37802 49258 37868 49274
rect 37802 49224 37818 49258
rect 37852 49256 37868 49258
rect 37852 49226 37890 49256
rect 38090 49226 38116 49256
rect 37852 49224 37868 49226
rect 37802 49208 37868 49224
rect 37802 48948 37868 48964
rect 37802 48914 37818 48948
rect 37852 48946 37868 48948
rect 37852 48916 37890 48946
rect 38090 48916 38116 48946
rect 37852 48914 37868 48916
rect 37802 48898 37868 48914
rect 38619 49258 38685 49274
rect 38619 49256 38635 49258
rect 38362 49226 38388 49256
rect 38588 49226 38635 49256
rect 38619 49224 38635 49226
rect 38669 49224 38685 49258
rect 38619 49208 38685 49224
rect 38619 48948 38685 48964
rect 38619 48946 38635 48948
rect 38362 48916 38388 48946
rect 38588 48916 38635 48946
rect 38619 48914 38635 48916
rect 38669 48914 38685 48948
rect 38619 48898 38685 48914
rect 42792 49258 42858 49274
rect 42792 49224 42808 49258
rect 42842 49256 42858 49258
rect 42842 49226 42880 49256
rect 43080 49226 43106 49256
rect 42842 49224 42858 49226
rect 42792 49208 42858 49224
rect 42792 48948 42858 48964
rect 42792 48914 42808 48948
rect 42842 48946 42858 48948
rect 42842 48916 42880 48946
rect 43080 48916 43106 48946
rect 42842 48914 42858 48916
rect 42792 48898 42858 48914
rect 43609 49258 43675 49274
rect 43609 49256 43625 49258
rect 43352 49226 43378 49256
rect 43578 49226 43625 49256
rect 43609 49224 43625 49226
rect 43659 49224 43675 49258
rect 43609 49208 43675 49224
rect 43609 48948 43675 48964
rect 43609 48946 43625 48948
rect 43352 48916 43378 48946
rect 43578 48916 43625 48946
rect 43609 48914 43625 48916
rect 43659 48914 43675 48948
rect 43609 48898 43675 48914
rect 47782 49258 47848 49274
rect 47782 49224 47798 49258
rect 47832 49256 47848 49258
rect 47832 49226 47870 49256
rect 48070 49226 48096 49256
rect 47832 49224 47848 49226
rect 47782 49208 47848 49224
rect 47782 48948 47848 48964
rect 47782 48914 47798 48948
rect 47832 48946 47848 48948
rect 47832 48916 47870 48946
rect 48070 48916 48096 48946
rect 47832 48914 47848 48916
rect 47782 48898 47848 48914
rect 48599 49258 48665 49274
rect 48599 49256 48615 49258
rect 48342 49226 48368 49256
rect 48568 49226 48615 49256
rect 48599 49224 48615 49226
rect 48649 49224 48665 49258
rect 48599 49208 48665 49224
rect 48599 48948 48665 48964
rect 48599 48946 48615 48948
rect 48342 48916 48368 48946
rect 48568 48916 48615 48946
rect 48599 48914 48615 48916
rect 48649 48914 48665 48948
rect 48599 48898 48665 48914
rect 52772 49258 52838 49274
rect 52772 49224 52788 49258
rect 52822 49256 52838 49258
rect 52822 49226 52860 49256
rect 53060 49226 53086 49256
rect 52822 49224 52838 49226
rect 52772 49208 52838 49224
rect 52772 48948 52838 48964
rect 52772 48914 52788 48948
rect 52822 48946 52838 48948
rect 52822 48916 52860 48946
rect 53060 48916 53086 48946
rect 52822 48914 52838 48916
rect 52772 48898 52838 48914
rect 53589 49258 53655 49274
rect 53589 49256 53605 49258
rect 53332 49226 53358 49256
rect 53558 49226 53605 49256
rect 53589 49224 53605 49226
rect 53639 49224 53655 49258
rect 53589 49208 53655 49224
rect 53589 48948 53655 48964
rect 53589 48946 53605 48948
rect 53332 48916 53358 48946
rect 53558 48916 53605 48946
rect 53589 48914 53605 48916
rect 53639 48914 53655 48948
rect 53589 48898 53655 48914
rect 57762 49258 57828 49274
rect 57762 49224 57778 49258
rect 57812 49256 57828 49258
rect 57812 49226 57850 49256
rect 58050 49226 58076 49256
rect 57812 49224 57828 49226
rect 57762 49208 57828 49224
rect 57762 48948 57828 48964
rect 57762 48914 57778 48948
rect 57812 48946 57828 48948
rect 57812 48916 57850 48946
rect 58050 48916 58076 48946
rect 57812 48914 57828 48916
rect 57762 48898 57828 48914
rect 58579 49258 58645 49274
rect 58579 49256 58595 49258
rect 58322 49226 58348 49256
rect 58548 49226 58595 49256
rect 58579 49224 58595 49226
rect 58629 49224 58645 49258
rect 58579 49208 58645 49224
rect 58579 48948 58645 48964
rect 58579 48946 58595 48948
rect 58322 48916 58348 48946
rect 58548 48916 58595 48946
rect 58579 48914 58595 48916
rect 58629 48914 58645 48948
rect 58579 48898 58645 48914
rect 62752 49258 62818 49274
rect 62752 49224 62768 49258
rect 62802 49256 62818 49258
rect 62802 49226 62840 49256
rect 63040 49226 63066 49256
rect 62802 49224 62818 49226
rect 62752 49208 62818 49224
rect 62752 48948 62818 48964
rect 62752 48914 62768 48948
rect 62802 48946 62818 48948
rect 62802 48916 62840 48946
rect 63040 48916 63066 48946
rect 62802 48914 62818 48916
rect 62752 48898 62818 48914
rect 63569 49258 63635 49274
rect 63569 49256 63585 49258
rect 63312 49226 63338 49256
rect 63538 49226 63585 49256
rect 63569 49224 63585 49226
rect 63619 49224 63635 49258
rect 63569 49208 63635 49224
rect 63569 48948 63635 48964
rect 63569 48946 63585 48948
rect 63312 48916 63338 48946
rect 63538 48916 63585 48946
rect 63569 48914 63585 48916
rect 63619 48914 63635 48948
rect 63569 48898 63635 48914
rect 67742 49258 67808 49274
rect 67742 49224 67758 49258
rect 67792 49256 67808 49258
rect 67792 49226 67830 49256
rect 68030 49226 68056 49256
rect 67792 49224 67808 49226
rect 67742 49208 67808 49224
rect 67742 48948 67808 48964
rect 67742 48914 67758 48948
rect 67792 48946 67808 48948
rect 67792 48916 67830 48946
rect 68030 48916 68056 48946
rect 67792 48914 67808 48916
rect 67742 48898 67808 48914
rect 68559 49258 68625 49274
rect 68559 49256 68575 49258
rect 68302 49226 68328 49256
rect 68528 49226 68575 49256
rect 68559 49224 68575 49226
rect 68609 49224 68625 49258
rect 68559 49208 68625 49224
rect 68559 48948 68625 48964
rect 68559 48946 68575 48948
rect 68302 48916 68328 48946
rect 68528 48916 68575 48946
rect 68559 48914 68575 48916
rect 68609 48914 68625 48948
rect 68559 48898 68625 48914
rect 72732 49258 72798 49274
rect 72732 49224 72748 49258
rect 72782 49256 72798 49258
rect 72782 49226 72820 49256
rect 73020 49226 73046 49256
rect 72782 49224 72798 49226
rect 72732 49208 72798 49224
rect 72732 48948 72798 48964
rect 72732 48914 72748 48948
rect 72782 48946 72798 48948
rect 72782 48916 72820 48946
rect 73020 48916 73046 48946
rect 72782 48914 72798 48916
rect 72732 48898 72798 48914
rect 73549 49258 73615 49274
rect 73549 49256 73565 49258
rect 73292 49226 73318 49256
rect 73518 49226 73565 49256
rect 73549 49224 73565 49226
rect 73599 49224 73615 49258
rect 73549 49208 73615 49224
rect 73549 48948 73615 48964
rect 73549 48946 73565 48948
rect 73292 48916 73318 48946
rect 73518 48916 73565 48946
rect 73549 48914 73565 48916
rect 73599 48914 73615 48948
rect 73549 48898 73615 48914
rect 77722 49258 77788 49274
rect 77722 49224 77738 49258
rect 77772 49256 77788 49258
rect 77772 49226 77810 49256
rect 78010 49226 78036 49256
rect 77772 49224 77788 49226
rect 77722 49208 77788 49224
rect 77722 48948 77788 48964
rect 77722 48914 77738 48948
rect 77772 48946 77788 48948
rect 77772 48916 77810 48946
rect 78010 48916 78036 48946
rect 77772 48914 77788 48916
rect 77722 48898 77788 48914
rect 78539 49258 78605 49274
rect 78539 49256 78555 49258
rect 78282 49226 78308 49256
rect 78508 49226 78555 49256
rect 78539 49224 78555 49226
rect 78589 49224 78605 49258
rect 78539 49208 78605 49224
rect 78539 48948 78605 48964
rect 78539 48946 78555 48948
rect 78282 48916 78308 48946
rect 78508 48916 78555 48946
rect 78539 48914 78555 48916
rect 78589 48914 78605 48948
rect 78539 48898 78605 48914
rect 2872 47548 2938 47564
rect 2872 47514 2888 47548
rect 2922 47546 2938 47548
rect 2922 47516 2960 47546
rect 3160 47516 3186 47546
rect 2922 47514 2938 47516
rect 2872 47498 2938 47514
rect 2872 47238 2938 47254
rect 2872 47204 2888 47238
rect 2922 47236 2938 47238
rect 2922 47206 2960 47236
rect 3160 47206 3186 47236
rect 2922 47204 2938 47206
rect 2872 47188 2938 47204
rect 3689 47548 3755 47564
rect 3689 47546 3705 47548
rect 3432 47516 3458 47546
rect 3658 47516 3705 47546
rect 3689 47514 3705 47516
rect 3739 47514 3755 47548
rect 3689 47498 3755 47514
rect 3689 47238 3755 47254
rect 3689 47236 3705 47238
rect 3432 47206 3458 47236
rect 3658 47206 3705 47236
rect 3689 47204 3705 47206
rect 3739 47204 3755 47238
rect 3689 47188 3755 47204
rect 7862 47548 7928 47564
rect 7862 47514 7878 47548
rect 7912 47546 7928 47548
rect 7912 47516 7950 47546
rect 8150 47516 8176 47546
rect 7912 47514 7928 47516
rect 7862 47498 7928 47514
rect 7862 47238 7928 47254
rect 7862 47204 7878 47238
rect 7912 47236 7928 47238
rect 7912 47206 7950 47236
rect 8150 47206 8176 47236
rect 7912 47204 7928 47206
rect 7862 47188 7928 47204
rect 8679 47548 8745 47564
rect 8679 47546 8695 47548
rect 8422 47516 8448 47546
rect 8648 47516 8695 47546
rect 8679 47514 8695 47516
rect 8729 47514 8745 47548
rect 8679 47498 8745 47514
rect 8679 47238 8745 47254
rect 8679 47236 8695 47238
rect 8422 47206 8448 47236
rect 8648 47206 8695 47236
rect 8679 47204 8695 47206
rect 8729 47204 8745 47238
rect 8679 47188 8745 47204
rect 12852 47548 12918 47564
rect 12852 47514 12868 47548
rect 12902 47546 12918 47548
rect 12902 47516 12940 47546
rect 13140 47516 13166 47546
rect 12902 47514 12918 47516
rect 12852 47498 12918 47514
rect 12852 47238 12918 47254
rect 12852 47204 12868 47238
rect 12902 47236 12918 47238
rect 12902 47206 12940 47236
rect 13140 47206 13166 47236
rect 12902 47204 12918 47206
rect 12852 47188 12918 47204
rect 13669 47548 13735 47564
rect 13669 47546 13685 47548
rect 13412 47516 13438 47546
rect 13638 47516 13685 47546
rect 13669 47514 13685 47516
rect 13719 47514 13735 47548
rect 13669 47498 13735 47514
rect 13669 47238 13735 47254
rect 13669 47236 13685 47238
rect 13412 47206 13438 47236
rect 13638 47206 13685 47236
rect 13669 47204 13685 47206
rect 13719 47204 13735 47238
rect 13669 47188 13735 47204
rect 17842 47548 17908 47564
rect 17842 47514 17858 47548
rect 17892 47546 17908 47548
rect 17892 47516 17930 47546
rect 18130 47516 18156 47546
rect 17892 47514 17908 47516
rect 17842 47498 17908 47514
rect 17842 47238 17908 47254
rect 17842 47204 17858 47238
rect 17892 47236 17908 47238
rect 17892 47206 17930 47236
rect 18130 47206 18156 47236
rect 17892 47204 17908 47206
rect 17842 47188 17908 47204
rect 18659 47548 18725 47564
rect 18659 47546 18675 47548
rect 18402 47516 18428 47546
rect 18628 47516 18675 47546
rect 18659 47514 18675 47516
rect 18709 47514 18725 47548
rect 18659 47498 18725 47514
rect 18659 47238 18725 47254
rect 18659 47236 18675 47238
rect 18402 47206 18428 47236
rect 18628 47206 18675 47236
rect 18659 47204 18675 47206
rect 18709 47204 18725 47238
rect 18659 47188 18725 47204
rect 22832 47548 22898 47564
rect 22832 47514 22848 47548
rect 22882 47546 22898 47548
rect 22882 47516 22920 47546
rect 23120 47516 23146 47546
rect 22882 47514 22898 47516
rect 22832 47498 22898 47514
rect 22832 47238 22898 47254
rect 22832 47204 22848 47238
rect 22882 47236 22898 47238
rect 22882 47206 22920 47236
rect 23120 47206 23146 47236
rect 22882 47204 22898 47206
rect 22832 47188 22898 47204
rect 23649 47548 23715 47564
rect 23649 47546 23665 47548
rect 23392 47516 23418 47546
rect 23618 47516 23665 47546
rect 23649 47514 23665 47516
rect 23699 47514 23715 47548
rect 23649 47498 23715 47514
rect 23649 47238 23715 47254
rect 23649 47236 23665 47238
rect 23392 47206 23418 47236
rect 23618 47206 23665 47236
rect 23649 47204 23665 47206
rect 23699 47204 23715 47238
rect 23649 47188 23715 47204
rect 27822 47548 27888 47564
rect 27822 47514 27838 47548
rect 27872 47546 27888 47548
rect 27872 47516 27910 47546
rect 28110 47516 28136 47546
rect 27872 47514 27888 47516
rect 27822 47498 27888 47514
rect 27822 47238 27888 47254
rect 27822 47204 27838 47238
rect 27872 47236 27888 47238
rect 27872 47206 27910 47236
rect 28110 47206 28136 47236
rect 27872 47204 27888 47206
rect 27822 47188 27888 47204
rect 28639 47548 28705 47564
rect 28639 47546 28655 47548
rect 28382 47516 28408 47546
rect 28608 47516 28655 47546
rect 28639 47514 28655 47516
rect 28689 47514 28705 47548
rect 28639 47498 28705 47514
rect 28639 47238 28705 47254
rect 28639 47236 28655 47238
rect 28382 47206 28408 47236
rect 28608 47206 28655 47236
rect 28639 47204 28655 47206
rect 28689 47204 28705 47238
rect 28639 47188 28705 47204
rect 32812 47548 32878 47564
rect 32812 47514 32828 47548
rect 32862 47546 32878 47548
rect 32862 47516 32900 47546
rect 33100 47516 33126 47546
rect 32862 47514 32878 47516
rect 32812 47498 32878 47514
rect 32812 47238 32878 47254
rect 32812 47204 32828 47238
rect 32862 47236 32878 47238
rect 32862 47206 32900 47236
rect 33100 47206 33126 47236
rect 32862 47204 32878 47206
rect 32812 47188 32878 47204
rect 33629 47548 33695 47564
rect 33629 47546 33645 47548
rect 33372 47516 33398 47546
rect 33598 47516 33645 47546
rect 33629 47514 33645 47516
rect 33679 47514 33695 47548
rect 33629 47498 33695 47514
rect 33629 47238 33695 47254
rect 33629 47236 33645 47238
rect 33372 47206 33398 47236
rect 33598 47206 33645 47236
rect 33629 47204 33645 47206
rect 33679 47204 33695 47238
rect 33629 47188 33695 47204
rect 37802 47548 37868 47564
rect 37802 47514 37818 47548
rect 37852 47546 37868 47548
rect 37852 47516 37890 47546
rect 38090 47516 38116 47546
rect 37852 47514 37868 47516
rect 37802 47498 37868 47514
rect 37802 47238 37868 47254
rect 37802 47204 37818 47238
rect 37852 47236 37868 47238
rect 37852 47206 37890 47236
rect 38090 47206 38116 47236
rect 37852 47204 37868 47206
rect 37802 47188 37868 47204
rect 38619 47548 38685 47564
rect 38619 47546 38635 47548
rect 38362 47516 38388 47546
rect 38588 47516 38635 47546
rect 38619 47514 38635 47516
rect 38669 47514 38685 47548
rect 38619 47498 38685 47514
rect 38619 47238 38685 47254
rect 38619 47236 38635 47238
rect 38362 47206 38388 47236
rect 38588 47206 38635 47236
rect 38619 47204 38635 47206
rect 38669 47204 38685 47238
rect 38619 47188 38685 47204
rect 42792 47548 42858 47564
rect 42792 47514 42808 47548
rect 42842 47546 42858 47548
rect 42842 47516 42880 47546
rect 43080 47516 43106 47546
rect 42842 47514 42858 47516
rect 42792 47498 42858 47514
rect 42792 47238 42858 47254
rect 42792 47204 42808 47238
rect 42842 47236 42858 47238
rect 42842 47206 42880 47236
rect 43080 47206 43106 47236
rect 42842 47204 42858 47206
rect 42792 47188 42858 47204
rect 43609 47548 43675 47564
rect 43609 47546 43625 47548
rect 43352 47516 43378 47546
rect 43578 47516 43625 47546
rect 43609 47514 43625 47516
rect 43659 47514 43675 47548
rect 43609 47498 43675 47514
rect 43609 47238 43675 47254
rect 43609 47236 43625 47238
rect 43352 47206 43378 47236
rect 43578 47206 43625 47236
rect 43609 47204 43625 47206
rect 43659 47204 43675 47238
rect 43609 47188 43675 47204
rect 47782 47548 47848 47564
rect 47782 47514 47798 47548
rect 47832 47546 47848 47548
rect 47832 47516 47870 47546
rect 48070 47516 48096 47546
rect 47832 47514 47848 47516
rect 47782 47498 47848 47514
rect 47782 47238 47848 47254
rect 47782 47204 47798 47238
rect 47832 47236 47848 47238
rect 47832 47206 47870 47236
rect 48070 47206 48096 47236
rect 47832 47204 47848 47206
rect 47782 47188 47848 47204
rect 48599 47548 48665 47564
rect 48599 47546 48615 47548
rect 48342 47516 48368 47546
rect 48568 47516 48615 47546
rect 48599 47514 48615 47516
rect 48649 47514 48665 47548
rect 48599 47498 48665 47514
rect 48599 47238 48665 47254
rect 48599 47236 48615 47238
rect 48342 47206 48368 47236
rect 48568 47206 48615 47236
rect 48599 47204 48615 47206
rect 48649 47204 48665 47238
rect 48599 47188 48665 47204
rect 52772 47548 52838 47564
rect 52772 47514 52788 47548
rect 52822 47546 52838 47548
rect 52822 47516 52860 47546
rect 53060 47516 53086 47546
rect 52822 47514 52838 47516
rect 52772 47498 52838 47514
rect 52772 47238 52838 47254
rect 52772 47204 52788 47238
rect 52822 47236 52838 47238
rect 52822 47206 52860 47236
rect 53060 47206 53086 47236
rect 52822 47204 52838 47206
rect 52772 47188 52838 47204
rect 53589 47548 53655 47564
rect 53589 47546 53605 47548
rect 53332 47516 53358 47546
rect 53558 47516 53605 47546
rect 53589 47514 53605 47516
rect 53639 47514 53655 47548
rect 53589 47498 53655 47514
rect 53589 47238 53655 47254
rect 53589 47236 53605 47238
rect 53332 47206 53358 47236
rect 53558 47206 53605 47236
rect 53589 47204 53605 47206
rect 53639 47204 53655 47238
rect 53589 47188 53655 47204
rect 57762 47548 57828 47564
rect 57762 47514 57778 47548
rect 57812 47546 57828 47548
rect 57812 47516 57850 47546
rect 58050 47516 58076 47546
rect 57812 47514 57828 47516
rect 57762 47498 57828 47514
rect 57762 47238 57828 47254
rect 57762 47204 57778 47238
rect 57812 47236 57828 47238
rect 57812 47206 57850 47236
rect 58050 47206 58076 47236
rect 57812 47204 57828 47206
rect 57762 47188 57828 47204
rect 58579 47548 58645 47564
rect 58579 47546 58595 47548
rect 58322 47516 58348 47546
rect 58548 47516 58595 47546
rect 58579 47514 58595 47516
rect 58629 47514 58645 47548
rect 58579 47498 58645 47514
rect 58579 47238 58645 47254
rect 58579 47236 58595 47238
rect 58322 47206 58348 47236
rect 58548 47206 58595 47236
rect 58579 47204 58595 47206
rect 58629 47204 58645 47238
rect 58579 47188 58645 47204
rect 62752 47548 62818 47564
rect 62752 47514 62768 47548
rect 62802 47546 62818 47548
rect 62802 47516 62840 47546
rect 63040 47516 63066 47546
rect 62802 47514 62818 47516
rect 62752 47498 62818 47514
rect 62752 47238 62818 47254
rect 62752 47204 62768 47238
rect 62802 47236 62818 47238
rect 62802 47206 62840 47236
rect 63040 47206 63066 47236
rect 62802 47204 62818 47206
rect 62752 47188 62818 47204
rect 63569 47548 63635 47564
rect 63569 47546 63585 47548
rect 63312 47516 63338 47546
rect 63538 47516 63585 47546
rect 63569 47514 63585 47516
rect 63619 47514 63635 47548
rect 63569 47498 63635 47514
rect 63569 47238 63635 47254
rect 63569 47236 63585 47238
rect 63312 47206 63338 47236
rect 63538 47206 63585 47236
rect 63569 47204 63585 47206
rect 63619 47204 63635 47238
rect 63569 47188 63635 47204
rect 67742 47548 67808 47564
rect 67742 47514 67758 47548
rect 67792 47546 67808 47548
rect 67792 47516 67830 47546
rect 68030 47516 68056 47546
rect 67792 47514 67808 47516
rect 67742 47498 67808 47514
rect 67742 47238 67808 47254
rect 67742 47204 67758 47238
rect 67792 47236 67808 47238
rect 67792 47206 67830 47236
rect 68030 47206 68056 47236
rect 67792 47204 67808 47206
rect 67742 47188 67808 47204
rect 68559 47548 68625 47564
rect 68559 47546 68575 47548
rect 68302 47516 68328 47546
rect 68528 47516 68575 47546
rect 68559 47514 68575 47516
rect 68609 47514 68625 47548
rect 68559 47498 68625 47514
rect 68559 47238 68625 47254
rect 68559 47236 68575 47238
rect 68302 47206 68328 47236
rect 68528 47206 68575 47236
rect 68559 47204 68575 47206
rect 68609 47204 68625 47238
rect 68559 47188 68625 47204
rect 72732 47548 72798 47564
rect 72732 47514 72748 47548
rect 72782 47546 72798 47548
rect 72782 47516 72820 47546
rect 73020 47516 73046 47546
rect 72782 47514 72798 47516
rect 72732 47498 72798 47514
rect 72732 47238 72798 47254
rect 72732 47204 72748 47238
rect 72782 47236 72798 47238
rect 72782 47206 72820 47236
rect 73020 47206 73046 47236
rect 72782 47204 72798 47206
rect 72732 47188 72798 47204
rect 73549 47548 73615 47564
rect 73549 47546 73565 47548
rect 73292 47516 73318 47546
rect 73518 47516 73565 47546
rect 73549 47514 73565 47516
rect 73599 47514 73615 47548
rect 73549 47498 73615 47514
rect 73549 47238 73615 47254
rect 73549 47236 73565 47238
rect 73292 47206 73318 47236
rect 73518 47206 73565 47236
rect 73549 47204 73565 47206
rect 73599 47204 73615 47238
rect 73549 47188 73615 47204
rect 77722 47548 77788 47564
rect 77722 47514 77738 47548
rect 77772 47546 77788 47548
rect 77772 47516 77810 47546
rect 78010 47516 78036 47546
rect 77772 47514 77788 47516
rect 77722 47498 77788 47514
rect 77722 47238 77788 47254
rect 77722 47204 77738 47238
rect 77772 47236 77788 47238
rect 77772 47206 77810 47236
rect 78010 47206 78036 47236
rect 77772 47204 77788 47206
rect 77722 47188 77788 47204
rect 78539 47548 78605 47564
rect 78539 47546 78555 47548
rect 78282 47516 78308 47546
rect 78508 47516 78555 47546
rect 78539 47514 78555 47516
rect 78589 47514 78605 47548
rect 78539 47498 78605 47514
rect 78539 47238 78605 47254
rect 78539 47236 78555 47238
rect 78282 47206 78308 47236
rect 78508 47206 78555 47236
rect 78539 47204 78555 47206
rect 78589 47204 78605 47238
rect 78539 47188 78605 47204
rect 2872 45838 2938 45854
rect 2872 45804 2888 45838
rect 2922 45836 2938 45838
rect 2922 45806 2960 45836
rect 3160 45806 3186 45836
rect 2922 45804 2938 45806
rect 2872 45788 2938 45804
rect 2872 45528 2938 45544
rect 2872 45494 2888 45528
rect 2922 45526 2938 45528
rect 2922 45496 2960 45526
rect 3160 45496 3186 45526
rect 2922 45494 2938 45496
rect 2872 45478 2938 45494
rect 3689 45838 3755 45854
rect 3689 45836 3705 45838
rect 3432 45806 3458 45836
rect 3658 45806 3705 45836
rect 3689 45804 3705 45806
rect 3739 45804 3755 45838
rect 3689 45788 3755 45804
rect 3689 45528 3755 45544
rect 3689 45526 3705 45528
rect 3432 45496 3458 45526
rect 3658 45496 3705 45526
rect 3689 45494 3705 45496
rect 3739 45494 3755 45528
rect 3689 45478 3755 45494
rect 7862 45838 7928 45854
rect 7862 45804 7878 45838
rect 7912 45836 7928 45838
rect 7912 45806 7950 45836
rect 8150 45806 8176 45836
rect 7912 45804 7928 45806
rect 7862 45788 7928 45804
rect 7862 45528 7928 45544
rect 7862 45494 7878 45528
rect 7912 45526 7928 45528
rect 7912 45496 7950 45526
rect 8150 45496 8176 45526
rect 7912 45494 7928 45496
rect 7862 45478 7928 45494
rect 8679 45838 8745 45854
rect 8679 45836 8695 45838
rect 8422 45806 8448 45836
rect 8648 45806 8695 45836
rect 8679 45804 8695 45806
rect 8729 45804 8745 45838
rect 8679 45788 8745 45804
rect 8679 45528 8745 45544
rect 8679 45526 8695 45528
rect 8422 45496 8448 45526
rect 8648 45496 8695 45526
rect 8679 45494 8695 45496
rect 8729 45494 8745 45528
rect 8679 45478 8745 45494
rect 12852 45838 12918 45854
rect 12852 45804 12868 45838
rect 12902 45836 12918 45838
rect 12902 45806 12940 45836
rect 13140 45806 13166 45836
rect 12902 45804 12918 45806
rect 12852 45788 12918 45804
rect 12852 45528 12918 45544
rect 12852 45494 12868 45528
rect 12902 45526 12918 45528
rect 12902 45496 12940 45526
rect 13140 45496 13166 45526
rect 12902 45494 12918 45496
rect 12852 45478 12918 45494
rect 13669 45838 13735 45854
rect 13669 45836 13685 45838
rect 13412 45806 13438 45836
rect 13638 45806 13685 45836
rect 13669 45804 13685 45806
rect 13719 45804 13735 45838
rect 13669 45788 13735 45804
rect 13669 45528 13735 45544
rect 13669 45526 13685 45528
rect 13412 45496 13438 45526
rect 13638 45496 13685 45526
rect 13669 45494 13685 45496
rect 13719 45494 13735 45528
rect 13669 45478 13735 45494
rect 17842 45838 17908 45854
rect 17842 45804 17858 45838
rect 17892 45836 17908 45838
rect 17892 45806 17930 45836
rect 18130 45806 18156 45836
rect 17892 45804 17908 45806
rect 17842 45788 17908 45804
rect 17842 45528 17908 45544
rect 17842 45494 17858 45528
rect 17892 45526 17908 45528
rect 17892 45496 17930 45526
rect 18130 45496 18156 45526
rect 17892 45494 17908 45496
rect 17842 45478 17908 45494
rect 18659 45838 18725 45854
rect 18659 45836 18675 45838
rect 18402 45806 18428 45836
rect 18628 45806 18675 45836
rect 18659 45804 18675 45806
rect 18709 45804 18725 45838
rect 18659 45788 18725 45804
rect 18659 45528 18725 45544
rect 18659 45526 18675 45528
rect 18402 45496 18428 45526
rect 18628 45496 18675 45526
rect 18659 45494 18675 45496
rect 18709 45494 18725 45528
rect 18659 45478 18725 45494
rect 22832 45838 22898 45854
rect 22832 45804 22848 45838
rect 22882 45836 22898 45838
rect 22882 45806 22920 45836
rect 23120 45806 23146 45836
rect 22882 45804 22898 45806
rect 22832 45788 22898 45804
rect 22832 45528 22898 45544
rect 22832 45494 22848 45528
rect 22882 45526 22898 45528
rect 22882 45496 22920 45526
rect 23120 45496 23146 45526
rect 22882 45494 22898 45496
rect 22832 45478 22898 45494
rect 23649 45838 23715 45854
rect 23649 45836 23665 45838
rect 23392 45806 23418 45836
rect 23618 45806 23665 45836
rect 23649 45804 23665 45806
rect 23699 45804 23715 45838
rect 23649 45788 23715 45804
rect 23649 45528 23715 45544
rect 23649 45526 23665 45528
rect 23392 45496 23418 45526
rect 23618 45496 23665 45526
rect 23649 45494 23665 45496
rect 23699 45494 23715 45528
rect 23649 45478 23715 45494
rect 27822 45838 27888 45854
rect 27822 45804 27838 45838
rect 27872 45836 27888 45838
rect 27872 45806 27910 45836
rect 28110 45806 28136 45836
rect 27872 45804 27888 45806
rect 27822 45788 27888 45804
rect 27822 45528 27888 45544
rect 27822 45494 27838 45528
rect 27872 45526 27888 45528
rect 27872 45496 27910 45526
rect 28110 45496 28136 45526
rect 27872 45494 27888 45496
rect 27822 45478 27888 45494
rect 28639 45838 28705 45854
rect 28639 45836 28655 45838
rect 28382 45806 28408 45836
rect 28608 45806 28655 45836
rect 28639 45804 28655 45806
rect 28689 45804 28705 45838
rect 28639 45788 28705 45804
rect 28639 45528 28705 45544
rect 28639 45526 28655 45528
rect 28382 45496 28408 45526
rect 28608 45496 28655 45526
rect 28639 45494 28655 45496
rect 28689 45494 28705 45528
rect 28639 45478 28705 45494
rect 32812 45838 32878 45854
rect 32812 45804 32828 45838
rect 32862 45836 32878 45838
rect 32862 45806 32900 45836
rect 33100 45806 33126 45836
rect 32862 45804 32878 45806
rect 32812 45788 32878 45804
rect 32812 45528 32878 45544
rect 32812 45494 32828 45528
rect 32862 45526 32878 45528
rect 32862 45496 32900 45526
rect 33100 45496 33126 45526
rect 32862 45494 32878 45496
rect 32812 45478 32878 45494
rect 33629 45838 33695 45854
rect 33629 45836 33645 45838
rect 33372 45806 33398 45836
rect 33598 45806 33645 45836
rect 33629 45804 33645 45806
rect 33679 45804 33695 45838
rect 33629 45788 33695 45804
rect 33629 45528 33695 45544
rect 33629 45526 33645 45528
rect 33372 45496 33398 45526
rect 33598 45496 33645 45526
rect 33629 45494 33645 45496
rect 33679 45494 33695 45528
rect 33629 45478 33695 45494
rect 37802 45838 37868 45854
rect 37802 45804 37818 45838
rect 37852 45836 37868 45838
rect 37852 45806 37890 45836
rect 38090 45806 38116 45836
rect 37852 45804 37868 45806
rect 37802 45788 37868 45804
rect 37802 45528 37868 45544
rect 37802 45494 37818 45528
rect 37852 45526 37868 45528
rect 37852 45496 37890 45526
rect 38090 45496 38116 45526
rect 37852 45494 37868 45496
rect 37802 45478 37868 45494
rect 38619 45838 38685 45854
rect 38619 45836 38635 45838
rect 38362 45806 38388 45836
rect 38588 45806 38635 45836
rect 38619 45804 38635 45806
rect 38669 45804 38685 45838
rect 38619 45788 38685 45804
rect 38619 45528 38685 45544
rect 38619 45526 38635 45528
rect 38362 45496 38388 45526
rect 38588 45496 38635 45526
rect 38619 45494 38635 45496
rect 38669 45494 38685 45528
rect 38619 45478 38685 45494
rect 42792 45838 42858 45854
rect 42792 45804 42808 45838
rect 42842 45836 42858 45838
rect 42842 45806 42880 45836
rect 43080 45806 43106 45836
rect 42842 45804 42858 45806
rect 42792 45788 42858 45804
rect 42792 45528 42858 45544
rect 42792 45494 42808 45528
rect 42842 45526 42858 45528
rect 42842 45496 42880 45526
rect 43080 45496 43106 45526
rect 42842 45494 42858 45496
rect 42792 45478 42858 45494
rect 43609 45838 43675 45854
rect 43609 45836 43625 45838
rect 43352 45806 43378 45836
rect 43578 45806 43625 45836
rect 43609 45804 43625 45806
rect 43659 45804 43675 45838
rect 43609 45788 43675 45804
rect 43609 45528 43675 45544
rect 43609 45526 43625 45528
rect 43352 45496 43378 45526
rect 43578 45496 43625 45526
rect 43609 45494 43625 45496
rect 43659 45494 43675 45528
rect 43609 45478 43675 45494
rect 47782 45838 47848 45854
rect 47782 45804 47798 45838
rect 47832 45836 47848 45838
rect 47832 45806 47870 45836
rect 48070 45806 48096 45836
rect 47832 45804 47848 45806
rect 47782 45788 47848 45804
rect 47782 45528 47848 45544
rect 47782 45494 47798 45528
rect 47832 45526 47848 45528
rect 47832 45496 47870 45526
rect 48070 45496 48096 45526
rect 47832 45494 47848 45496
rect 47782 45478 47848 45494
rect 48599 45838 48665 45854
rect 48599 45836 48615 45838
rect 48342 45806 48368 45836
rect 48568 45806 48615 45836
rect 48599 45804 48615 45806
rect 48649 45804 48665 45838
rect 48599 45788 48665 45804
rect 48599 45528 48665 45544
rect 48599 45526 48615 45528
rect 48342 45496 48368 45526
rect 48568 45496 48615 45526
rect 48599 45494 48615 45496
rect 48649 45494 48665 45528
rect 48599 45478 48665 45494
rect 52772 45838 52838 45854
rect 52772 45804 52788 45838
rect 52822 45836 52838 45838
rect 52822 45806 52860 45836
rect 53060 45806 53086 45836
rect 52822 45804 52838 45806
rect 52772 45788 52838 45804
rect 52772 45528 52838 45544
rect 52772 45494 52788 45528
rect 52822 45526 52838 45528
rect 52822 45496 52860 45526
rect 53060 45496 53086 45526
rect 52822 45494 52838 45496
rect 52772 45478 52838 45494
rect 53589 45838 53655 45854
rect 53589 45836 53605 45838
rect 53332 45806 53358 45836
rect 53558 45806 53605 45836
rect 53589 45804 53605 45806
rect 53639 45804 53655 45838
rect 53589 45788 53655 45804
rect 53589 45528 53655 45544
rect 53589 45526 53605 45528
rect 53332 45496 53358 45526
rect 53558 45496 53605 45526
rect 53589 45494 53605 45496
rect 53639 45494 53655 45528
rect 53589 45478 53655 45494
rect 57762 45838 57828 45854
rect 57762 45804 57778 45838
rect 57812 45836 57828 45838
rect 57812 45806 57850 45836
rect 58050 45806 58076 45836
rect 57812 45804 57828 45806
rect 57762 45788 57828 45804
rect 57762 45528 57828 45544
rect 57762 45494 57778 45528
rect 57812 45526 57828 45528
rect 57812 45496 57850 45526
rect 58050 45496 58076 45526
rect 57812 45494 57828 45496
rect 57762 45478 57828 45494
rect 58579 45838 58645 45854
rect 58579 45836 58595 45838
rect 58322 45806 58348 45836
rect 58548 45806 58595 45836
rect 58579 45804 58595 45806
rect 58629 45804 58645 45838
rect 58579 45788 58645 45804
rect 58579 45528 58645 45544
rect 58579 45526 58595 45528
rect 58322 45496 58348 45526
rect 58548 45496 58595 45526
rect 58579 45494 58595 45496
rect 58629 45494 58645 45528
rect 58579 45478 58645 45494
rect 62752 45838 62818 45854
rect 62752 45804 62768 45838
rect 62802 45836 62818 45838
rect 62802 45806 62840 45836
rect 63040 45806 63066 45836
rect 62802 45804 62818 45806
rect 62752 45788 62818 45804
rect 62752 45528 62818 45544
rect 62752 45494 62768 45528
rect 62802 45526 62818 45528
rect 62802 45496 62840 45526
rect 63040 45496 63066 45526
rect 62802 45494 62818 45496
rect 62752 45478 62818 45494
rect 63569 45838 63635 45854
rect 63569 45836 63585 45838
rect 63312 45806 63338 45836
rect 63538 45806 63585 45836
rect 63569 45804 63585 45806
rect 63619 45804 63635 45838
rect 63569 45788 63635 45804
rect 63569 45528 63635 45544
rect 63569 45526 63585 45528
rect 63312 45496 63338 45526
rect 63538 45496 63585 45526
rect 63569 45494 63585 45496
rect 63619 45494 63635 45528
rect 63569 45478 63635 45494
rect 67742 45838 67808 45854
rect 67742 45804 67758 45838
rect 67792 45836 67808 45838
rect 67792 45806 67830 45836
rect 68030 45806 68056 45836
rect 67792 45804 67808 45806
rect 67742 45788 67808 45804
rect 67742 45528 67808 45544
rect 67742 45494 67758 45528
rect 67792 45526 67808 45528
rect 67792 45496 67830 45526
rect 68030 45496 68056 45526
rect 67792 45494 67808 45496
rect 67742 45478 67808 45494
rect 68559 45838 68625 45854
rect 68559 45836 68575 45838
rect 68302 45806 68328 45836
rect 68528 45806 68575 45836
rect 68559 45804 68575 45806
rect 68609 45804 68625 45838
rect 68559 45788 68625 45804
rect 68559 45528 68625 45544
rect 68559 45526 68575 45528
rect 68302 45496 68328 45526
rect 68528 45496 68575 45526
rect 68559 45494 68575 45496
rect 68609 45494 68625 45528
rect 68559 45478 68625 45494
rect 72732 45838 72798 45854
rect 72732 45804 72748 45838
rect 72782 45836 72798 45838
rect 72782 45806 72820 45836
rect 73020 45806 73046 45836
rect 72782 45804 72798 45806
rect 72732 45788 72798 45804
rect 72732 45528 72798 45544
rect 72732 45494 72748 45528
rect 72782 45526 72798 45528
rect 72782 45496 72820 45526
rect 73020 45496 73046 45526
rect 72782 45494 72798 45496
rect 72732 45478 72798 45494
rect 73549 45838 73615 45854
rect 73549 45836 73565 45838
rect 73292 45806 73318 45836
rect 73518 45806 73565 45836
rect 73549 45804 73565 45806
rect 73599 45804 73615 45838
rect 73549 45788 73615 45804
rect 73549 45528 73615 45544
rect 73549 45526 73565 45528
rect 73292 45496 73318 45526
rect 73518 45496 73565 45526
rect 73549 45494 73565 45496
rect 73599 45494 73615 45528
rect 73549 45478 73615 45494
rect 77722 45838 77788 45854
rect 77722 45804 77738 45838
rect 77772 45836 77788 45838
rect 77772 45806 77810 45836
rect 78010 45806 78036 45836
rect 77772 45804 77788 45806
rect 77722 45788 77788 45804
rect 77722 45528 77788 45544
rect 77722 45494 77738 45528
rect 77772 45526 77788 45528
rect 77772 45496 77810 45526
rect 78010 45496 78036 45526
rect 77772 45494 77788 45496
rect 77722 45478 77788 45494
rect 78539 45838 78605 45854
rect 78539 45836 78555 45838
rect 78282 45806 78308 45836
rect 78508 45806 78555 45836
rect 78539 45804 78555 45806
rect 78589 45804 78605 45838
rect 78539 45788 78605 45804
rect 78539 45528 78605 45544
rect 78539 45526 78555 45528
rect 78282 45496 78308 45526
rect 78508 45496 78555 45526
rect 78539 45494 78555 45496
rect 78589 45494 78605 45528
rect 78539 45478 78605 45494
rect 2872 44128 2938 44144
rect 2872 44094 2888 44128
rect 2922 44126 2938 44128
rect 2922 44096 2960 44126
rect 3160 44096 3186 44126
rect 2922 44094 2938 44096
rect 2872 44078 2938 44094
rect 2872 43818 2938 43834
rect 2872 43784 2888 43818
rect 2922 43816 2938 43818
rect 2922 43786 2960 43816
rect 3160 43786 3186 43816
rect 2922 43784 2938 43786
rect 2872 43768 2938 43784
rect 3689 44128 3755 44144
rect 3689 44126 3705 44128
rect 3432 44096 3458 44126
rect 3658 44096 3705 44126
rect 3689 44094 3705 44096
rect 3739 44094 3755 44128
rect 3689 44078 3755 44094
rect 3689 43818 3755 43834
rect 3689 43816 3705 43818
rect 3432 43786 3458 43816
rect 3658 43786 3705 43816
rect 3689 43784 3705 43786
rect 3739 43784 3755 43818
rect 3689 43768 3755 43784
rect 7862 44128 7928 44144
rect 7862 44094 7878 44128
rect 7912 44126 7928 44128
rect 7912 44096 7950 44126
rect 8150 44096 8176 44126
rect 7912 44094 7928 44096
rect 7862 44078 7928 44094
rect 7862 43818 7928 43834
rect 7862 43784 7878 43818
rect 7912 43816 7928 43818
rect 7912 43786 7950 43816
rect 8150 43786 8176 43816
rect 7912 43784 7928 43786
rect 7862 43768 7928 43784
rect 8679 44128 8745 44144
rect 8679 44126 8695 44128
rect 8422 44096 8448 44126
rect 8648 44096 8695 44126
rect 8679 44094 8695 44096
rect 8729 44094 8745 44128
rect 8679 44078 8745 44094
rect 8679 43818 8745 43834
rect 8679 43816 8695 43818
rect 8422 43786 8448 43816
rect 8648 43786 8695 43816
rect 8679 43784 8695 43786
rect 8729 43784 8745 43818
rect 8679 43768 8745 43784
rect 12852 44128 12918 44144
rect 12852 44094 12868 44128
rect 12902 44126 12918 44128
rect 12902 44096 12940 44126
rect 13140 44096 13166 44126
rect 12902 44094 12918 44096
rect 12852 44078 12918 44094
rect 12852 43818 12918 43834
rect 12852 43784 12868 43818
rect 12902 43816 12918 43818
rect 12902 43786 12940 43816
rect 13140 43786 13166 43816
rect 12902 43784 12918 43786
rect 12852 43768 12918 43784
rect 13669 44128 13735 44144
rect 13669 44126 13685 44128
rect 13412 44096 13438 44126
rect 13638 44096 13685 44126
rect 13669 44094 13685 44096
rect 13719 44094 13735 44128
rect 13669 44078 13735 44094
rect 13669 43818 13735 43834
rect 13669 43816 13685 43818
rect 13412 43786 13438 43816
rect 13638 43786 13685 43816
rect 13669 43784 13685 43786
rect 13719 43784 13735 43818
rect 13669 43768 13735 43784
rect 17842 44128 17908 44144
rect 17842 44094 17858 44128
rect 17892 44126 17908 44128
rect 17892 44096 17930 44126
rect 18130 44096 18156 44126
rect 17892 44094 17908 44096
rect 17842 44078 17908 44094
rect 17842 43818 17908 43834
rect 17842 43784 17858 43818
rect 17892 43816 17908 43818
rect 17892 43786 17930 43816
rect 18130 43786 18156 43816
rect 17892 43784 17908 43786
rect 17842 43768 17908 43784
rect 18659 44128 18725 44144
rect 18659 44126 18675 44128
rect 18402 44096 18428 44126
rect 18628 44096 18675 44126
rect 18659 44094 18675 44096
rect 18709 44094 18725 44128
rect 18659 44078 18725 44094
rect 18659 43818 18725 43834
rect 18659 43816 18675 43818
rect 18402 43786 18428 43816
rect 18628 43786 18675 43816
rect 18659 43784 18675 43786
rect 18709 43784 18725 43818
rect 18659 43768 18725 43784
rect 22832 44128 22898 44144
rect 22832 44094 22848 44128
rect 22882 44126 22898 44128
rect 22882 44096 22920 44126
rect 23120 44096 23146 44126
rect 22882 44094 22898 44096
rect 22832 44078 22898 44094
rect 22832 43818 22898 43834
rect 22832 43784 22848 43818
rect 22882 43816 22898 43818
rect 22882 43786 22920 43816
rect 23120 43786 23146 43816
rect 22882 43784 22898 43786
rect 22832 43768 22898 43784
rect 23649 44128 23715 44144
rect 23649 44126 23665 44128
rect 23392 44096 23418 44126
rect 23618 44096 23665 44126
rect 23649 44094 23665 44096
rect 23699 44094 23715 44128
rect 23649 44078 23715 44094
rect 23649 43818 23715 43834
rect 23649 43816 23665 43818
rect 23392 43786 23418 43816
rect 23618 43786 23665 43816
rect 23649 43784 23665 43786
rect 23699 43784 23715 43818
rect 23649 43768 23715 43784
rect 27822 44128 27888 44144
rect 27822 44094 27838 44128
rect 27872 44126 27888 44128
rect 27872 44096 27910 44126
rect 28110 44096 28136 44126
rect 27872 44094 27888 44096
rect 27822 44078 27888 44094
rect 27822 43818 27888 43834
rect 27822 43784 27838 43818
rect 27872 43816 27888 43818
rect 27872 43786 27910 43816
rect 28110 43786 28136 43816
rect 27872 43784 27888 43786
rect 27822 43768 27888 43784
rect 28639 44128 28705 44144
rect 28639 44126 28655 44128
rect 28382 44096 28408 44126
rect 28608 44096 28655 44126
rect 28639 44094 28655 44096
rect 28689 44094 28705 44128
rect 28639 44078 28705 44094
rect 28639 43818 28705 43834
rect 28639 43816 28655 43818
rect 28382 43786 28408 43816
rect 28608 43786 28655 43816
rect 28639 43784 28655 43786
rect 28689 43784 28705 43818
rect 28639 43768 28705 43784
rect 32812 44128 32878 44144
rect 32812 44094 32828 44128
rect 32862 44126 32878 44128
rect 32862 44096 32900 44126
rect 33100 44096 33126 44126
rect 32862 44094 32878 44096
rect 32812 44078 32878 44094
rect 32812 43818 32878 43834
rect 32812 43784 32828 43818
rect 32862 43816 32878 43818
rect 32862 43786 32900 43816
rect 33100 43786 33126 43816
rect 32862 43784 32878 43786
rect 32812 43768 32878 43784
rect 33629 44128 33695 44144
rect 33629 44126 33645 44128
rect 33372 44096 33398 44126
rect 33598 44096 33645 44126
rect 33629 44094 33645 44096
rect 33679 44094 33695 44128
rect 33629 44078 33695 44094
rect 33629 43818 33695 43834
rect 33629 43816 33645 43818
rect 33372 43786 33398 43816
rect 33598 43786 33645 43816
rect 33629 43784 33645 43786
rect 33679 43784 33695 43818
rect 33629 43768 33695 43784
rect 37802 44128 37868 44144
rect 37802 44094 37818 44128
rect 37852 44126 37868 44128
rect 37852 44096 37890 44126
rect 38090 44096 38116 44126
rect 37852 44094 37868 44096
rect 37802 44078 37868 44094
rect 37802 43818 37868 43834
rect 37802 43784 37818 43818
rect 37852 43816 37868 43818
rect 37852 43786 37890 43816
rect 38090 43786 38116 43816
rect 37852 43784 37868 43786
rect 37802 43768 37868 43784
rect 38619 44128 38685 44144
rect 38619 44126 38635 44128
rect 38362 44096 38388 44126
rect 38588 44096 38635 44126
rect 38619 44094 38635 44096
rect 38669 44094 38685 44128
rect 38619 44078 38685 44094
rect 38619 43818 38685 43834
rect 38619 43816 38635 43818
rect 38362 43786 38388 43816
rect 38588 43786 38635 43816
rect 38619 43784 38635 43786
rect 38669 43784 38685 43818
rect 38619 43768 38685 43784
rect 42792 44128 42858 44144
rect 42792 44094 42808 44128
rect 42842 44126 42858 44128
rect 42842 44096 42880 44126
rect 43080 44096 43106 44126
rect 42842 44094 42858 44096
rect 42792 44078 42858 44094
rect 42792 43818 42858 43834
rect 42792 43784 42808 43818
rect 42842 43816 42858 43818
rect 42842 43786 42880 43816
rect 43080 43786 43106 43816
rect 42842 43784 42858 43786
rect 42792 43768 42858 43784
rect 43609 44128 43675 44144
rect 43609 44126 43625 44128
rect 43352 44096 43378 44126
rect 43578 44096 43625 44126
rect 43609 44094 43625 44096
rect 43659 44094 43675 44128
rect 43609 44078 43675 44094
rect 43609 43818 43675 43834
rect 43609 43816 43625 43818
rect 43352 43786 43378 43816
rect 43578 43786 43625 43816
rect 43609 43784 43625 43786
rect 43659 43784 43675 43818
rect 43609 43768 43675 43784
rect 47782 44128 47848 44144
rect 47782 44094 47798 44128
rect 47832 44126 47848 44128
rect 47832 44096 47870 44126
rect 48070 44096 48096 44126
rect 47832 44094 47848 44096
rect 47782 44078 47848 44094
rect 47782 43818 47848 43834
rect 47782 43784 47798 43818
rect 47832 43816 47848 43818
rect 47832 43786 47870 43816
rect 48070 43786 48096 43816
rect 47832 43784 47848 43786
rect 47782 43768 47848 43784
rect 48599 44128 48665 44144
rect 48599 44126 48615 44128
rect 48342 44096 48368 44126
rect 48568 44096 48615 44126
rect 48599 44094 48615 44096
rect 48649 44094 48665 44128
rect 48599 44078 48665 44094
rect 48599 43818 48665 43834
rect 48599 43816 48615 43818
rect 48342 43786 48368 43816
rect 48568 43786 48615 43816
rect 48599 43784 48615 43786
rect 48649 43784 48665 43818
rect 48599 43768 48665 43784
rect 52772 44128 52838 44144
rect 52772 44094 52788 44128
rect 52822 44126 52838 44128
rect 52822 44096 52860 44126
rect 53060 44096 53086 44126
rect 52822 44094 52838 44096
rect 52772 44078 52838 44094
rect 52772 43818 52838 43834
rect 52772 43784 52788 43818
rect 52822 43816 52838 43818
rect 52822 43786 52860 43816
rect 53060 43786 53086 43816
rect 52822 43784 52838 43786
rect 52772 43768 52838 43784
rect 53589 44128 53655 44144
rect 53589 44126 53605 44128
rect 53332 44096 53358 44126
rect 53558 44096 53605 44126
rect 53589 44094 53605 44096
rect 53639 44094 53655 44128
rect 53589 44078 53655 44094
rect 53589 43818 53655 43834
rect 53589 43816 53605 43818
rect 53332 43786 53358 43816
rect 53558 43786 53605 43816
rect 53589 43784 53605 43786
rect 53639 43784 53655 43818
rect 53589 43768 53655 43784
rect 57762 44128 57828 44144
rect 57762 44094 57778 44128
rect 57812 44126 57828 44128
rect 57812 44096 57850 44126
rect 58050 44096 58076 44126
rect 57812 44094 57828 44096
rect 57762 44078 57828 44094
rect 57762 43818 57828 43834
rect 57762 43784 57778 43818
rect 57812 43816 57828 43818
rect 57812 43786 57850 43816
rect 58050 43786 58076 43816
rect 57812 43784 57828 43786
rect 57762 43768 57828 43784
rect 58579 44128 58645 44144
rect 58579 44126 58595 44128
rect 58322 44096 58348 44126
rect 58548 44096 58595 44126
rect 58579 44094 58595 44096
rect 58629 44094 58645 44128
rect 58579 44078 58645 44094
rect 58579 43818 58645 43834
rect 58579 43816 58595 43818
rect 58322 43786 58348 43816
rect 58548 43786 58595 43816
rect 58579 43784 58595 43786
rect 58629 43784 58645 43818
rect 58579 43768 58645 43784
rect 62752 44128 62818 44144
rect 62752 44094 62768 44128
rect 62802 44126 62818 44128
rect 62802 44096 62840 44126
rect 63040 44096 63066 44126
rect 62802 44094 62818 44096
rect 62752 44078 62818 44094
rect 62752 43818 62818 43834
rect 62752 43784 62768 43818
rect 62802 43816 62818 43818
rect 62802 43786 62840 43816
rect 63040 43786 63066 43816
rect 62802 43784 62818 43786
rect 62752 43768 62818 43784
rect 63569 44128 63635 44144
rect 63569 44126 63585 44128
rect 63312 44096 63338 44126
rect 63538 44096 63585 44126
rect 63569 44094 63585 44096
rect 63619 44094 63635 44128
rect 63569 44078 63635 44094
rect 63569 43818 63635 43834
rect 63569 43816 63585 43818
rect 63312 43786 63338 43816
rect 63538 43786 63585 43816
rect 63569 43784 63585 43786
rect 63619 43784 63635 43818
rect 63569 43768 63635 43784
rect 67742 44128 67808 44144
rect 67742 44094 67758 44128
rect 67792 44126 67808 44128
rect 67792 44096 67830 44126
rect 68030 44096 68056 44126
rect 67792 44094 67808 44096
rect 67742 44078 67808 44094
rect 67742 43818 67808 43834
rect 67742 43784 67758 43818
rect 67792 43816 67808 43818
rect 67792 43786 67830 43816
rect 68030 43786 68056 43816
rect 67792 43784 67808 43786
rect 67742 43768 67808 43784
rect 68559 44128 68625 44144
rect 68559 44126 68575 44128
rect 68302 44096 68328 44126
rect 68528 44096 68575 44126
rect 68559 44094 68575 44096
rect 68609 44094 68625 44128
rect 68559 44078 68625 44094
rect 68559 43818 68625 43834
rect 68559 43816 68575 43818
rect 68302 43786 68328 43816
rect 68528 43786 68575 43816
rect 68559 43784 68575 43786
rect 68609 43784 68625 43818
rect 68559 43768 68625 43784
rect 72732 44128 72798 44144
rect 72732 44094 72748 44128
rect 72782 44126 72798 44128
rect 72782 44096 72820 44126
rect 73020 44096 73046 44126
rect 72782 44094 72798 44096
rect 72732 44078 72798 44094
rect 72732 43818 72798 43834
rect 72732 43784 72748 43818
rect 72782 43816 72798 43818
rect 72782 43786 72820 43816
rect 73020 43786 73046 43816
rect 72782 43784 72798 43786
rect 72732 43768 72798 43784
rect 73549 44128 73615 44144
rect 73549 44126 73565 44128
rect 73292 44096 73318 44126
rect 73518 44096 73565 44126
rect 73549 44094 73565 44096
rect 73599 44094 73615 44128
rect 73549 44078 73615 44094
rect 73549 43818 73615 43834
rect 73549 43816 73565 43818
rect 73292 43786 73318 43816
rect 73518 43786 73565 43816
rect 73549 43784 73565 43786
rect 73599 43784 73615 43818
rect 73549 43768 73615 43784
rect 77722 44128 77788 44144
rect 77722 44094 77738 44128
rect 77772 44126 77788 44128
rect 77772 44096 77810 44126
rect 78010 44096 78036 44126
rect 77772 44094 77788 44096
rect 77722 44078 77788 44094
rect 77722 43818 77788 43834
rect 77722 43784 77738 43818
rect 77772 43816 77788 43818
rect 77772 43786 77810 43816
rect 78010 43786 78036 43816
rect 77772 43784 77788 43786
rect 77722 43768 77788 43784
rect 78539 44128 78605 44144
rect 78539 44126 78555 44128
rect 78282 44096 78308 44126
rect 78508 44096 78555 44126
rect 78539 44094 78555 44096
rect 78589 44094 78605 44128
rect 78539 44078 78605 44094
rect 78539 43818 78605 43834
rect 78539 43816 78555 43818
rect 78282 43786 78308 43816
rect 78508 43786 78555 43816
rect 78539 43784 78555 43786
rect 78589 43784 78605 43818
rect 78539 43768 78605 43784
rect 2872 42418 2938 42434
rect 2872 42384 2888 42418
rect 2922 42416 2938 42418
rect 2922 42386 2960 42416
rect 3160 42386 3186 42416
rect 2922 42384 2938 42386
rect 2872 42368 2938 42384
rect 2872 42108 2938 42124
rect 2872 42074 2888 42108
rect 2922 42106 2938 42108
rect 2922 42076 2960 42106
rect 3160 42076 3186 42106
rect 2922 42074 2938 42076
rect 2872 42058 2938 42074
rect 3689 42418 3755 42434
rect 3689 42416 3705 42418
rect 3432 42386 3458 42416
rect 3658 42386 3705 42416
rect 3689 42384 3705 42386
rect 3739 42384 3755 42418
rect 3689 42368 3755 42384
rect 3689 42108 3755 42124
rect 3689 42106 3705 42108
rect 3432 42076 3458 42106
rect 3658 42076 3705 42106
rect 3689 42074 3705 42076
rect 3739 42074 3755 42108
rect 3689 42058 3755 42074
rect 7862 42418 7928 42434
rect 7862 42384 7878 42418
rect 7912 42416 7928 42418
rect 7912 42386 7950 42416
rect 8150 42386 8176 42416
rect 7912 42384 7928 42386
rect 7862 42368 7928 42384
rect 7862 42108 7928 42124
rect 7862 42074 7878 42108
rect 7912 42106 7928 42108
rect 7912 42076 7950 42106
rect 8150 42076 8176 42106
rect 7912 42074 7928 42076
rect 7862 42058 7928 42074
rect 8679 42418 8745 42434
rect 8679 42416 8695 42418
rect 8422 42386 8448 42416
rect 8648 42386 8695 42416
rect 8679 42384 8695 42386
rect 8729 42384 8745 42418
rect 8679 42368 8745 42384
rect 8679 42108 8745 42124
rect 8679 42106 8695 42108
rect 8422 42076 8448 42106
rect 8648 42076 8695 42106
rect 8679 42074 8695 42076
rect 8729 42074 8745 42108
rect 8679 42058 8745 42074
rect 12852 42418 12918 42434
rect 12852 42384 12868 42418
rect 12902 42416 12918 42418
rect 12902 42386 12940 42416
rect 13140 42386 13166 42416
rect 12902 42384 12918 42386
rect 12852 42368 12918 42384
rect 12852 42108 12918 42124
rect 12852 42074 12868 42108
rect 12902 42106 12918 42108
rect 12902 42076 12940 42106
rect 13140 42076 13166 42106
rect 12902 42074 12918 42076
rect 12852 42058 12918 42074
rect 13669 42418 13735 42434
rect 13669 42416 13685 42418
rect 13412 42386 13438 42416
rect 13638 42386 13685 42416
rect 13669 42384 13685 42386
rect 13719 42384 13735 42418
rect 13669 42368 13735 42384
rect 13669 42108 13735 42124
rect 13669 42106 13685 42108
rect 13412 42076 13438 42106
rect 13638 42076 13685 42106
rect 13669 42074 13685 42076
rect 13719 42074 13735 42108
rect 13669 42058 13735 42074
rect 17842 42418 17908 42434
rect 17842 42384 17858 42418
rect 17892 42416 17908 42418
rect 17892 42386 17930 42416
rect 18130 42386 18156 42416
rect 17892 42384 17908 42386
rect 17842 42368 17908 42384
rect 17842 42108 17908 42124
rect 17842 42074 17858 42108
rect 17892 42106 17908 42108
rect 17892 42076 17930 42106
rect 18130 42076 18156 42106
rect 17892 42074 17908 42076
rect 17842 42058 17908 42074
rect 18659 42418 18725 42434
rect 18659 42416 18675 42418
rect 18402 42386 18428 42416
rect 18628 42386 18675 42416
rect 18659 42384 18675 42386
rect 18709 42384 18725 42418
rect 18659 42368 18725 42384
rect 18659 42108 18725 42124
rect 18659 42106 18675 42108
rect 18402 42076 18428 42106
rect 18628 42076 18675 42106
rect 18659 42074 18675 42076
rect 18709 42074 18725 42108
rect 18659 42058 18725 42074
rect 22832 42418 22898 42434
rect 22832 42384 22848 42418
rect 22882 42416 22898 42418
rect 22882 42386 22920 42416
rect 23120 42386 23146 42416
rect 22882 42384 22898 42386
rect 22832 42368 22898 42384
rect 22832 42108 22898 42124
rect 22832 42074 22848 42108
rect 22882 42106 22898 42108
rect 22882 42076 22920 42106
rect 23120 42076 23146 42106
rect 22882 42074 22898 42076
rect 22832 42058 22898 42074
rect 23649 42418 23715 42434
rect 23649 42416 23665 42418
rect 23392 42386 23418 42416
rect 23618 42386 23665 42416
rect 23649 42384 23665 42386
rect 23699 42384 23715 42418
rect 23649 42368 23715 42384
rect 23649 42108 23715 42124
rect 23649 42106 23665 42108
rect 23392 42076 23418 42106
rect 23618 42076 23665 42106
rect 23649 42074 23665 42076
rect 23699 42074 23715 42108
rect 23649 42058 23715 42074
rect 27822 42418 27888 42434
rect 27822 42384 27838 42418
rect 27872 42416 27888 42418
rect 27872 42386 27910 42416
rect 28110 42386 28136 42416
rect 27872 42384 27888 42386
rect 27822 42368 27888 42384
rect 27822 42108 27888 42124
rect 27822 42074 27838 42108
rect 27872 42106 27888 42108
rect 27872 42076 27910 42106
rect 28110 42076 28136 42106
rect 27872 42074 27888 42076
rect 27822 42058 27888 42074
rect 28639 42418 28705 42434
rect 28639 42416 28655 42418
rect 28382 42386 28408 42416
rect 28608 42386 28655 42416
rect 28639 42384 28655 42386
rect 28689 42384 28705 42418
rect 28639 42368 28705 42384
rect 28639 42108 28705 42124
rect 28639 42106 28655 42108
rect 28382 42076 28408 42106
rect 28608 42076 28655 42106
rect 28639 42074 28655 42076
rect 28689 42074 28705 42108
rect 28639 42058 28705 42074
rect 32812 42418 32878 42434
rect 32812 42384 32828 42418
rect 32862 42416 32878 42418
rect 32862 42386 32900 42416
rect 33100 42386 33126 42416
rect 32862 42384 32878 42386
rect 32812 42368 32878 42384
rect 32812 42108 32878 42124
rect 32812 42074 32828 42108
rect 32862 42106 32878 42108
rect 32862 42076 32900 42106
rect 33100 42076 33126 42106
rect 32862 42074 32878 42076
rect 32812 42058 32878 42074
rect 33629 42418 33695 42434
rect 33629 42416 33645 42418
rect 33372 42386 33398 42416
rect 33598 42386 33645 42416
rect 33629 42384 33645 42386
rect 33679 42384 33695 42418
rect 33629 42368 33695 42384
rect 33629 42108 33695 42124
rect 33629 42106 33645 42108
rect 33372 42076 33398 42106
rect 33598 42076 33645 42106
rect 33629 42074 33645 42076
rect 33679 42074 33695 42108
rect 33629 42058 33695 42074
rect 37802 42418 37868 42434
rect 37802 42384 37818 42418
rect 37852 42416 37868 42418
rect 37852 42386 37890 42416
rect 38090 42386 38116 42416
rect 37852 42384 37868 42386
rect 37802 42368 37868 42384
rect 37802 42108 37868 42124
rect 37802 42074 37818 42108
rect 37852 42106 37868 42108
rect 37852 42076 37890 42106
rect 38090 42076 38116 42106
rect 37852 42074 37868 42076
rect 37802 42058 37868 42074
rect 38619 42418 38685 42434
rect 38619 42416 38635 42418
rect 38362 42386 38388 42416
rect 38588 42386 38635 42416
rect 38619 42384 38635 42386
rect 38669 42384 38685 42418
rect 38619 42368 38685 42384
rect 38619 42108 38685 42124
rect 38619 42106 38635 42108
rect 38362 42076 38388 42106
rect 38588 42076 38635 42106
rect 38619 42074 38635 42076
rect 38669 42074 38685 42108
rect 38619 42058 38685 42074
rect 42792 42418 42858 42434
rect 42792 42384 42808 42418
rect 42842 42416 42858 42418
rect 42842 42386 42880 42416
rect 43080 42386 43106 42416
rect 42842 42384 42858 42386
rect 42792 42368 42858 42384
rect 42792 42108 42858 42124
rect 42792 42074 42808 42108
rect 42842 42106 42858 42108
rect 42842 42076 42880 42106
rect 43080 42076 43106 42106
rect 42842 42074 42858 42076
rect 42792 42058 42858 42074
rect 43609 42418 43675 42434
rect 43609 42416 43625 42418
rect 43352 42386 43378 42416
rect 43578 42386 43625 42416
rect 43609 42384 43625 42386
rect 43659 42384 43675 42418
rect 43609 42368 43675 42384
rect 43609 42108 43675 42124
rect 43609 42106 43625 42108
rect 43352 42076 43378 42106
rect 43578 42076 43625 42106
rect 43609 42074 43625 42076
rect 43659 42074 43675 42108
rect 43609 42058 43675 42074
rect 47782 42418 47848 42434
rect 47782 42384 47798 42418
rect 47832 42416 47848 42418
rect 47832 42386 47870 42416
rect 48070 42386 48096 42416
rect 47832 42384 47848 42386
rect 47782 42368 47848 42384
rect 47782 42108 47848 42124
rect 47782 42074 47798 42108
rect 47832 42106 47848 42108
rect 47832 42076 47870 42106
rect 48070 42076 48096 42106
rect 47832 42074 47848 42076
rect 47782 42058 47848 42074
rect 48599 42418 48665 42434
rect 48599 42416 48615 42418
rect 48342 42386 48368 42416
rect 48568 42386 48615 42416
rect 48599 42384 48615 42386
rect 48649 42384 48665 42418
rect 48599 42368 48665 42384
rect 48599 42108 48665 42124
rect 48599 42106 48615 42108
rect 48342 42076 48368 42106
rect 48568 42076 48615 42106
rect 48599 42074 48615 42076
rect 48649 42074 48665 42108
rect 48599 42058 48665 42074
rect 52772 42418 52838 42434
rect 52772 42384 52788 42418
rect 52822 42416 52838 42418
rect 52822 42386 52860 42416
rect 53060 42386 53086 42416
rect 52822 42384 52838 42386
rect 52772 42368 52838 42384
rect 52772 42108 52838 42124
rect 52772 42074 52788 42108
rect 52822 42106 52838 42108
rect 52822 42076 52860 42106
rect 53060 42076 53086 42106
rect 52822 42074 52838 42076
rect 52772 42058 52838 42074
rect 53589 42418 53655 42434
rect 53589 42416 53605 42418
rect 53332 42386 53358 42416
rect 53558 42386 53605 42416
rect 53589 42384 53605 42386
rect 53639 42384 53655 42418
rect 53589 42368 53655 42384
rect 53589 42108 53655 42124
rect 53589 42106 53605 42108
rect 53332 42076 53358 42106
rect 53558 42076 53605 42106
rect 53589 42074 53605 42076
rect 53639 42074 53655 42108
rect 53589 42058 53655 42074
rect 57762 42418 57828 42434
rect 57762 42384 57778 42418
rect 57812 42416 57828 42418
rect 57812 42386 57850 42416
rect 58050 42386 58076 42416
rect 57812 42384 57828 42386
rect 57762 42368 57828 42384
rect 57762 42108 57828 42124
rect 57762 42074 57778 42108
rect 57812 42106 57828 42108
rect 57812 42076 57850 42106
rect 58050 42076 58076 42106
rect 57812 42074 57828 42076
rect 57762 42058 57828 42074
rect 58579 42418 58645 42434
rect 58579 42416 58595 42418
rect 58322 42386 58348 42416
rect 58548 42386 58595 42416
rect 58579 42384 58595 42386
rect 58629 42384 58645 42418
rect 58579 42368 58645 42384
rect 58579 42108 58645 42124
rect 58579 42106 58595 42108
rect 58322 42076 58348 42106
rect 58548 42076 58595 42106
rect 58579 42074 58595 42076
rect 58629 42074 58645 42108
rect 58579 42058 58645 42074
rect 62752 42418 62818 42434
rect 62752 42384 62768 42418
rect 62802 42416 62818 42418
rect 62802 42386 62840 42416
rect 63040 42386 63066 42416
rect 62802 42384 62818 42386
rect 62752 42368 62818 42384
rect 62752 42108 62818 42124
rect 62752 42074 62768 42108
rect 62802 42106 62818 42108
rect 62802 42076 62840 42106
rect 63040 42076 63066 42106
rect 62802 42074 62818 42076
rect 62752 42058 62818 42074
rect 63569 42418 63635 42434
rect 63569 42416 63585 42418
rect 63312 42386 63338 42416
rect 63538 42386 63585 42416
rect 63569 42384 63585 42386
rect 63619 42384 63635 42418
rect 63569 42368 63635 42384
rect 63569 42108 63635 42124
rect 63569 42106 63585 42108
rect 63312 42076 63338 42106
rect 63538 42076 63585 42106
rect 63569 42074 63585 42076
rect 63619 42074 63635 42108
rect 63569 42058 63635 42074
rect 67742 42418 67808 42434
rect 67742 42384 67758 42418
rect 67792 42416 67808 42418
rect 67792 42386 67830 42416
rect 68030 42386 68056 42416
rect 67792 42384 67808 42386
rect 67742 42368 67808 42384
rect 67742 42108 67808 42124
rect 67742 42074 67758 42108
rect 67792 42106 67808 42108
rect 67792 42076 67830 42106
rect 68030 42076 68056 42106
rect 67792 42074 67808 42076
rect 67742 42058 67808 42074
rect 68559 42418 68625 42434
rect 68559 42416 68575 42418
rect 68302 42386 68328 42416
rect 68528 42386 68575 42416
rect 68559 42384 68575 42386
rect 68609 42384 68625 42418
rect 68559 42368 68625 42384
rect 68559 42108 68625 42124
rect 68559 42106 68575 42108
rect 68302 42076 68328 42106
rect 68528 42076 68575 42106
rect 68559 42074 68575 42076
rect 68609 42074 68625 42108
rect 68559 42058 68625 42074
rect 72732 42418 72798 42434
rect 72732 42384 72748 42418
rect 72782 42416 72798 42418
rect 72782 42386 72820 42416
rect 73020 42386 73046 42416
rect 72782 42384 72798 42386
rect 72732 42368 72798 42384
rect 72732 42108 72798 42124
rect 72732 42074 72748 42108
rect 72782 42106 72798 42108
rect 72782 42076 72820 42106
rect 73020 42076 73046 42106
rect 72782 42074 72798 42076
rect 72732 42058 72798 42074
rect 73549 42418 73615 42434
rect 73549 42416 73565 42418
rect 73292 42386 73318 42416
rect 73518 42386 73565 42416
rect 73549 42384 73565 42386
rect 73599 42384 73615 42418
rect 73549 42368 73615 42384
rect 73549 42108 73615 42124
rect 73549 42106 73565 42108
rect 73292 42076 73318 42106
rect 73518 42076 73565 42106
rect 73549 42074 73565 42076
rect 73599 42074 73615 42108
rect 73549 42058 73615 42074
rect 77722 42418 77788 42434
rect 77722 42384 77738 42418
rect 77772 42416 77788 42418
rect 77772 42386 77810 42416
rect 78010 42386 78036 42416
rect 77772 42384 77788 42386
rect 77722 42368 77788 42384
rect 77722 42108 77788 42124
rect 77722 42074 77738 42108
rect 77772 42106 77788 42108
rect 77772 42076 77810 42106
rect 78010 42076 78036 42106
rect 77772 42074 77788 42076
rect 77722 42058 77788 42074
rect 78539 42418 78605 42434
rect 78539 42416 78555 42418
rect 78282 42386 78308 42416
rect 78508 42386 78555 42416
rect 78539 42384 78555 42386
rect 78589 42384 78605 42418
rect 78539 42368 78605 42384
rect 78539 42108 78605 42124
rect 78539 42106 78555 42108
rect 78282 42076 78308 42106
rect 78508 42076 78555 42106
rect 78539 42074 78555 42076
rect 78589 42074 78605 42108
rect 78539 42058 78605 42074
rect 2872 40708 2938 40724
rect 2872 40674 2888 40708
rect 2922 40706 2938 40708
rect 2922 40676 2960 40706
rect 3160 40676 3186 40706
rect 2922 40674 2938 40676
rect 2872 40658 2938 40674
rect 2872 40398 2938 40414
rect 2872 40364 2888 40398
rect 2922 40396 2938 40398
rect 2922 40366 2960 40396
rect 3160 40366 3186 40396
rect 2922 40364 2938 40366
rect 2872 40348 2938 40364
rect 3689 40708 3755 40724
rect 3689 40706 3705 40708
rect 3432 40676 3458 40706
rect 3658 40676 3705 40706
rect 3689 40674 3705 40676
rect 3739 40674 3755 40708
rect 3689 40658 3755 40674
rect 3689 40398 3755 40414
rect 3689 40396 3705 40398
rect 3432 40366 3458 40396
rect 3658 40366 3705 40396
rect 3689 40364 3705 40366
rect 3739 40364 3755 40398
rect 3689 40348 3755 40364
rect 7862 40708 7928 40724
rect 7862 40674 7878 40708
rect 7912 40706 7928 40708
rect 7912 40676 7950 40706
rect 8150 40676 8176 40706
rect 7912 40674 7928 40676
rect 7862 40658 7928 40674
rect 7862 40398 7928 40414
rect 7862 40364 7878 40398
rect 7912 40396 7928 40398
rect 7912 40366 7950 40396
rect 8150 40366 8176 40396
rect 7912 40364 7928 40366
rect 7862 40348 7928 40364
rect 8679 40708 8745 40724
rect 8679 40706 8695 40708
rect 8422 40676 8448 40706
rect 8648 40676 8695 40706
rect 8679 40674 8695 40676
rect 8729 40674 8745 40708
rect 8679 40658 8745 40674
rect 8679 40398 8745 40414
rect 8679 40396 8695 40398
rect 8422 40366 8448 40396
rect 8648 40366 8695 40396
rect 8679 40364 8695 40366
rect 8729 40364 8745 40398
rect 8679 40348 8745 40364
rect 12852 40708 12918 40724
rect 12852 40674 12868 40708
rect 12902 40706 12918 40708
rect 12902 40676 12940 40706
rect 13140 40676 13166 40706
rect 12902 40674 12918 40676
rect 12852 40658 12918 40674
rect 12852 40398 12918 40414
rect 12852 40364 12868 40398
rect 12902 40396 12918 40398
rect 12902 40366 12940 40396
rect 13140 40366 13166 40396
rect 12902 40364 12918 40366
rect 12852 40348 12918 40364
rect 13669 40708 13735 40724
rect 13669 40706 13685 40708
rect 13412 40676 13438 40706
rect 13638 40676 13685 40706
rect 13669 40674 13685 40676
rect 13719 40674 13735 40708
rect 13669 40658 13735 40674
rect 13669 40398 13735 40414
rect 13669 40396 13685 40398
rect 13412 40366 13438 40396
rect 13638 40366 13685 40396
rect 13669 40364 13685 40366
rect 13719 40364 13735 40398
rect 13669 40348 13735 40364
rect 17842 40708 17908 40724
rect 17842 40674 17858 40708
rect 17892 40706 17908 40708
rect 17892 40676 17930 40706
rect 18130 40676 18156 40706
rect 17892 40674 17908 40676
rect 17842 40658 17908 40674
rect 17842 40398 17908 40414
rect 17842 40364 17858 40398
rect 17892 40396 17908 40398
rect 17892 40366 17930 40396
rect 18130 40366 18156 40396
rect 17892 40364 17908 40366
rect 17842 40348 17908 40364
rect 18659 40708 18725 40724
rect 18659 40706 18675 40708
rect 18402 40676 18428 40706
rect 18628 40676 18675 40706
rect 18659 40674 18675 40676
rect 18709 40674 18725 40708
rect 18659 40658 18725 40674
rect 18659 40398 18725 40414
rect 18659 40396 18675 40398
rect 18402 40366 18428 40396
rect 18628 40366 18675 40396
rect 18659 40364 18675 40366
rect 18709 40364 18725 40398
rect 18659 40348 18725 40364
rect 22832 40708 22898 40724
rect 22832 40674 22848 40708
rect 22882 40706 22898 40708
rect 22882 40676 22920 40706
rect 23120 40676 23146 40706
rect 22882 40674 22898 40676
rect 22832 40658 22898 40674
rect 22832 40398 22898 40414
rect 22832 40364 22848 40398
rect 22882 40396 22898 40398
rect 22882 40366 22920 40396
rect 23120 40366 23146 40396
rect 22882 40364 22898 40366
rect 22832 40348 22898 40364
rect 23649 40708 23715 40724
rect 23649 40706 23665 40708
rect 23392 40676 23418 40706
rect 23618 40676 23665 40706
rect 23649 40674 23665 40676
rect 23699 40674 23715 40708
rect 23649 40658 23715 40674
rect 23649 40398 23715 40414
rect 23649 40396 23665 40398
rect 23392 40366 23418 40396
rect 23618 40366 23665 40396
rect 23649 40364 23665 40366
rect 23699 40364 23715 40398
rect 23649 40348 23715 40364
rect 27822 40708 27888 40724
rect 27822 40674 27838 40708
rect 27872 40706 27888 40708
rect 27872 40676 27910 40706
rect 28110 40676 28136 40706
rect 27872 40674 27888 40676
rect 27822 40658 27888 40674
rect 27822 40398 27888 40414
rect 27822 40364 27838 40398
rect 27872 40396 27888 40398
rect 27872 40366 27910 40396
rect 28110 40366 28136 40396
rect 27872 40364 27888 40366
rect 27822 40348 27888 40364
rect 28639 40708 28705 40724
rect 28639 40706 28655 40708
rect 28382 40676 28408 40706
rect 28608 40676 28655 40706
rect 28639 40674 28655 40676
rect 28689 40674 28705 40708
rect 28639 40658 28705 40674
rect 28639 40398 28705 40414
rect 28639 40396 28655 40398
rect 28382 40366 28408 40396
rect 28608 40366 28655 40396
rect 28639 40364 28655 40366
rect 28689 40364 28705 40398
rect 28639 40348 28705 40364
rect 32812 40708 32878 40724
rect 32812 40674 32828 40708
rect 32862 40706 32878 40708
rect 32862 40676 32900 40706
rect 33100 40676 33126 40706
rect 32862 40674 32878 40676
rect 32812 40658 32878 40674
rect 32812 40398 32878 40414
rect 32812 40364 32828 40398
rect 32862 40396 32878 40398
rect 32862 40366 32900 40396
rect 33100 40366 33126 40396
rect 32862 40364 32878 40366
rect 32812 40348 32878 40364
rect 33629 40708 33695 40724
rect 33629 40706 33645 40708
rect 33372 40676 33398 40706
rect 33598 40676 33645 40706
rect 33629 40674 33645 40676
rect 33679 40674 33695 40708
rect 33629 40658 33695 40674
rect 33629 40398 33695 40414
rect 33629 40396 33645 40398
rect 33372 40366 33398 40396
rect 33598 40366 33645 40396
rect 33629 40364 33645 40366
rect 33679 40364 33695 40398
rect 33629 40348 33695 40364
rect 37802 40708 37868 40724
rect 37802 40674 37818 40708
rect 37852 40706 37868 40708
rect 37852 40676 37890 40706
rect 38090 40676 38116 40706
rect 37852 40674 37868 40676
rect 37802 40658 37868 40674
rect 37802 40398 37868 40414
rect 37802 40364 37818 40398
rect 37852 40396 37868 40398
rect 37852 40366 37890 40396
rect 38090 40366 38116 40396
rect 37852 40364 37868 40366
rect 37802 40348 37868 40364
rect 38619 40708 38685 40724
rect 38619 40706 38635 40708
rect 38362 40676 38388 40706
rect 38588 40676 38635 40706
rect 38619 40674 38635 40676
rect 38669 40674 38685 40708
rect 38619 40658 38685 40674
rect 38619 40398 38685 40414
rect 38619 40396 38635 40398
rect 38362 40366 38388 40396
rect 38588 40366 38635 40396
rect 38619 40364 38635 40366
rect 38669 40364 38685 40398
rect 38619 40348 38685 40364
rect 42792 40708 42858 40724
rect 42792 40674 42808 40708
rect 42842 40706 42858 40708
rect 42842 40676 42880 40706
rect 43080 40676 43106 40706
rect 42842 40674 42858 40676
rect 42792 40658 42858 40674
rect 42792 40398 42858 40414
rect 42792 40364 42808 40398
rect 42842 40396 42858 40398
rect 42842 40366 42880 40396
rect 43080 40366 43106 40396
rect 42842 40364 42858 40366
rect 42792 40348 42858 40364
rect 43609 40708 43675 40724
rect 43609 40706 43625 40708
rect 43352 40676 43378 40706
rect 43578 40676 43625 40706
rect 43609 40674 43625 40676
rect 43659 40674 43675 40708
rect 43609 40658 43675 40674
rect 43609 40398 43675 40414
rect 43609 40396 43625 40398
rect 43352 40366 43378 40396
rect 43578 40366 43625 40396
rect 43609 40364 43625 40366
rect 43659 40364 43675 40398
rect 43609 40348 43675 40364
rect 47782 40708 47848 40724
rect 47782 40674 47798 40708
rect 47832 40706 47848 40708
rect 47832 40676 47870 40706
rect 48070 40676 48096 40706
rect 47832 40674 47848 40676
rect 47782 40658 47848 40674
rect 47782 40398 47848 40414
rect 47782 40364 47798 40398
rect 47832 40396 47848 40398
rect 47832 40366 47870 40396
rect 48070 40366 48096 40396
rect 47832 40364 47848 40366
rect 47782 40348 47848 40364
rect 48599 40708 48665 40724
rect 48599 40706 48615 40708
rect 48342 40676 48368 40706
rect 48568 40676 48615 40706
rect 48599 40674 48615 40676
rect 48649 40674 48665 40708
rect 48599 40658 48665 40674
rect 48599 40398 48665 40414
rect 48599 40396 48615 40398
rect 48342 40366 48368 40396
rect 48568 40366 48615 40396
rect 48599 40364 48615 40366
rect 48649 40364 48665 40398
rect 48599 40348 48665 40364
rect 52772 40708 52838 40724
rect 52772 40674 52788 40708
rect 52822 40706 52838 40708
rect 52822 40676 52860 40706
rect 53060 40676 53086 40706
rect 52822 40674 52838 40676
rect 52772 40658 52838 40674
rect 52772 40398 52838 40414
rect 52772 40364 52788 40398
rect 52822 40396 52838 40398
rect 52822 40366 52860 40396
rect 53060 40366 53086 40396
rect 52822 40364 52838 40366
rect 52772 40348 52838 40364
rect 53589 40708 53655 40724
rect 53589 40706 53605 40708
rect 53332 40676 53358 40706
rect 53558 40676 53605 40706
rect 53589 40674 53605 40676
rect 53639 40674 53655 40708
rect 53589 40658 53655 40674
rect 53589 40398 53655 40414
rect 53589 40396 53605 40398
rect 53332 40366 53358 40396
rect 53558 40366 53605 40396
rect 53589 40364 53605 40366
rect 53639 40364 53655 40398
rect 53589 40348 53655 40364
rect 57762 40708 57828 40724
rect 57762 40674 57778 40708
rect 57812 40706 57828 40708
rect 57812 40676 57850 40706
rect 58050 40676 58076 40706
rect 57812 40674 57828 40676
rect 57762 40658 57828 40674
rect 57762 40398 57828 40414
rect 57762 40364 57778 40398
rect 57812 40396 57828 40398
rect 57812 40366 57850 40396
rect 58050 40366 58076 40396
rect 57812 40364 57828 40366
rect 57762 40348 57828 40364
rect 58579 40708 58645 40724
rect 58579 40706 58595 40708
rect 58322 40676 58348 40706
rect 58548 40676 58595 40706
rect 58579 40674 58595 40676
rect 58629 40674 58645 40708
rect 58579 40658 58645 40674
rect 58579 40398 58645 40414
rect 58579 40396 58595 40398
rect 58322 40366 58348 40396
rect 58548 40366 58595 40396
rect 58579 40364 58595 40366
rect 58629 40364 58645 40398
rect 58579 40348 58645 40364
rect 62752 40708 62818 40724
rect 62752 40674 62768 40708
rect 62802 40706 62818 40708
rect 62802 40676 62840 40706
rect 63040 40676 63066 40706
rect 62802 40674 62818 40676
rect 62752 40658 62818 40674
rect 62752 40398 62818 40414
rect 62752 40364 62768 40398
rect 62802 40396 62818 40398
rect 62802 40366 62840 40396
rect 63040 40366 63066 40396
rect 62802 40364 62818 40366
rect 62752 40348 62818 40364
rect 63569 40708 63635 40724
rect 63569 40706 63585 40708
rect 63312 40676 63338 40706
rect 63538 40676 63585 40706
rect 63569 40674 63585 40676
rect 63619 40674 63635 40708
rect 63569 40658 63635 40674
rect 63569 40398 63635 40414
rect 63569 40396 63585 40398
rect 63312 40366 63338 40396
rect 63538 40366 63585 40396
rect 63569 40364 63585 40366
rect 63619 40364 63635 40398
rect 63569 40348 63635 40364
rect 67742 40708 67808 40724
rect 67742 40674 67758 40708
rect 67792 40706 67808 40708
rect 67792 40676 67830 40706
rect 68030 40676 68056 40706
rect 67792 40674 67808 40676
rect 67742 40658 67808 40674
rect 67742 40398 67808 40414
rect 67742 40364 67758 40398
rect 67792 40396 67808 40398
rect 67792 40366 67830 40396
rect 68030 40366 68056 40396
rect 67792 40364 67808 40366
rect 67742 40348 67808 40364
rect 68559 40708 68625 40724
rect 68559 40706 68575 40708
rect 68302 40676 68328 40706
rect 68528 40676 68575 40706
rect 68559 40674 68575 40676
rect 68609 40674 68625 40708
rect 68559 40658 68625 40674
rect 68559 40398 68625 40414
rect 68559 40396 68575 40398
rect 68302 40366 68328 40396
rect 68528 40366 68575 40396
rect 68559 40364 68575 40366
rect 68609 40364 68625 40398
rect 68559 40348 68625 40364
rect 72732 40708 72798 40724
rect 72732 40674 72748 40708
rect 72782 40706 72798 40708
rect 72782 40676 72820 40706
rect 73020 40676 73046 40706
rect 72782 40674 72798 40676
rect 72732 40658 72798 40674
rect 72732 40398 72798 40414
rect 72732 40364 72748 40398
rect 72782 40396 72798 40398
rect 72782 40366 72820 40396
rect 73020 40366 73046 40396
rect 72782 40364 72798 40366
rect 72732 40348 72798 40364
rect 73549 40708 73615 40724
rect 73549 40706 73565 40708
rect 73292 40676 73318 40706
rect 73518 40676 73565 40706
rect 73549 40674 73565 40676
rect 73599 40674 73615 40708
rect 73549 40658 73615 40674
rect 73549 40398 73615 40414
rect 73549 40396 73565 40398
rect 73292 40366 73318 40396
rect 73518 40366 73565 40396
rect 73549 40364 73565 40366
rect 73599 40364 73615 40398
rect 73549 40348 73615 40364
rect 77722 40708 77788 40724
rect 77722 40674 77738 40708
rect 77772 40706 77788 40708
rect 77772 40676 77810 40706
rect 78010 40676 78036 40706
rect 77772 40674 77788 40676
rect 77722 40658 77788 40674
rect 77722 40398 77788 40414
rect 77722 40364 77738 40398
rect 77772 40396 77788 40398
rect 77772 40366 77810 40396
rect 78010 40366 78036 40396
rect 77772 40364 77788 40366
rect 77722 40348 77788 40364
rect 78539 40708 78605 40724
rect 78539 40706 78555 40708
rect 78282 40676 78308 40706
rect 78508 40676 78555 40706
rect 78539 40674 78555 40676
rect 78589 40674 78605 40708
rect 78539 40658 78605 40674
rect 78539 40398 78605 40414
rect 78539 40396 78555 40398
rect 78282 40366 78308 40396
rect 78508 40366 78555 40396
rect 78539 40364 78555 40366
rect 78589 40364 78605 40398
rect 78539 40348 78605 40364
<< polycont >>
rect 2888 66324 2922 66358
rect 2888 66014 2922 66048
rect 3705 66324 3739 66358
rect 3705 66014 3739 66048
rect 7878 66324 7912 66358
rect 7878 66014 7912 66048
rect 8695 66324 8729 66358
rect 8695 66014 8729 66048
rect 12868 66324 12902 66358
rect 12868 66014 12902 66048
rect 13685 66324 13719 66358
rect 13685 66014 13719 66048
rect 17858 66324 17892 66358
rect 17858 66014 17892 66048
rect 18675 66324 18709 66358
rect 18675 66014 18709 66048
rect 22848 66324 22882 66358
rect 22848 66014 22882 66048
rect 23665 66324 23699 66358
rect 23665 66014 23699 66048
rect 27838 66324 27872 66358
rect 27838 66014 27872 66048
rect 28655 66324 28689 66358
rect 28655 66014 28689 66048
rect 32828 66324 32862 66358
rect 32828 66014 32862 66048
rect 33645 66324 33679 66358
rect 33645 66014 33679 66048
rect 37818 66324 37852 66358
rect 37818 66014 37852 66048
rect 38635 66324 38669 66358
rect 38635 66014 38669 66048
rect 42808 66324 42842 66358
rect 42808 66014 42842 66048
rect 43625 66324 43659 66358
rect 43625 66014 43659 66048
rect 47798 66324 47832 66358
rect 47798 66014 47832 66048
rect 48615 66324 48649 66358
rect 48615 66014 48649 66048
rect 52788 66324 52822 66358
rect 52788 66014 52822 66048
rect 53605 66324 53639 66358
rect 53605 66014 53639 66048
rect 57778 66324 57812 66358
rect 57778 66014 57812 66048
rect 58595 66324 58629 66358
rect 58595 66014 58629 66048
rect 62768 66324 62802 66358
rect 62768 66014 62802 66048
rect 63585 66324 63619 66358
rect 63585 66014 63619 66048
rect 67758 66324 67792 66358
rect 67758 66014 67792 66048
rect 68575 66324 68609 66358
rect 68575 66014 68609 66048
rect 72748 66324 72782 66358
rect 72748 66014 72782 66048
rect 73565 66324 73599 66358
rect 73565 66014 73599 66048
rect 77738 66324 77772 66358
rect 77738 66014 77772 66048
rect 78555 66324 78589 66358
rect 78555 66014 78589 66048
rect 2888 64614 2922 64648
rect 2888 64304 2922 64338
rect 3705 64614 3739 64648
rect 3705 64304 3739 64338
rect 7878 64614 7912 64648
rect 7878 64304 7912 64338
rect 8695 64614 8729 64648
rect 8695 64304 8729 64338
rect 12868 64614 12902 64648
rect 12868 64304 12902 64338
rect 13685 64614 13719 64648
rect 13685 64304 13719 64338
rect 17858 64614 17892 64648
rect 17858 64304 17892 64338
rect 18675 64614 18709 64648
rect 18675 64304 18709 64338
rect 22848 64614 22882 64648
rect 22848 64304 22882 64338
rect 23665 64614 23699 64648
rect 23665 64304 23699 64338
rect 27838 64614 27872 64648
rect 27838 64304 27872 64338
rect 28655 64614 28689 64648
rect 28655 64304 28689 64338
rect 32828 64614 32862 64648
rect 32828 64304 32862 64338
rect 33645 64614 33679 64648
rect 33645 64304 33679 64338
rect 37818 64614 37852 64648
rect 37818 64304 37852 64338
rect 38635 64614 38669 64648
rect 38635 64304 38669 64338
rect 42808 64614 42842 64648
rect 42808 64304 42842 64338
rect 43625 64614 43659 64648
rect 43625 64304 43659 64338
rect 47798 64614 47832 64648
rect 47798 64304 47832 64338
rect 48615 64614 48649 64648
rect 48615 64304 48649 64338
rect 52788 64614 52822 64648
rect 52788 64304 52822 64338
rect 53605 64614 53639 64648
rect 53605 64304 53639 64338
rect 57778 64614 57812 64648
rect 57778 64304 57812 64338
rect 58595 64614 58629 64648
rect 58595 64304 58629 64338
rect 62768 64614 62802 64648
rect 62768 64304 62802 64338
rect 63585 64614 63619 64648
rect 63585 64304 63619 64338
rect 67758 64614 67792 64648
rect 67758 64304 67792 64338
rect 68575 64614 68609 64648
rect 68575 64304 68609 64338
rect 72748 64614 72782 64648
rect 72748 64304 72782 64338
rect 73565 64614 73599 64648
rect 73565 64304 73599 64338
rect 77738 64614 77772 64648
rect 77738 64304 77772 64338
rect 78555 64614 78589 64648
rect 78555 64304 78589 64338
rect 2888 62904 2922 62938
rect 2888 62594 2922 62628
rect 3705 62904 3739 62938
rect 3705 62594 3739 62628
rect 7878 62904 7912 62938
rect 7878 62594 7912 62628
rect 8695 62904 8729 62938
rect 8695 62594 8729 62628
rect 12868 62904 12902 62938
rect 12868 62594 12902 62628
rect 13685 62904 13719 62938
rect 13685 62594 13719 62628
rect 17858 62904 17892 62938
rect 17858 62594 17892 62628
rect 18675 62904 18709 62938
rect 18675 62594 18709 62628
rect 22848 62904 22882 62938
rect 22848 62594 22882 62628
rect 23665 62904 23699 62938
rect 23665 62594 23699 62628
rect 27838 62904 27872 62938
rect 27838 62594 27872 62628
rect 28655 62904 28689 62938
rect 28655 62594 28689 62628
rect 32828 62904 32862 62938
rect 32828 62594 32862 62628
rect 33645 62904 33679 62938
rect 33645 62594 33679 62628
rect 37818 62904 37852 62938
rect 37818 62594 37852 62628
rect 38635 62904 38669 62938
rect 38635 62594 38669 62628
rect 42808 62904 42842 62938
rect 42808 62594 42842 62628
rect 43625 62904 43659 62938
rect 43625 62594 43659 62628
rect 47798 62904 47832 62938
rect 47798 62594 47832 62628
rect 48615 62904 48649 62938
rect 48615 62594 48649 62628
rect 52788 62904 52822 62938
rect 52788 62594 52822 62628
rect 53605 62904 53639 62938
rect 53605 62594 53639 62628
rect 57778 62904 57812 62938
rect 57778 62594 57812 62628
rect 58595 62904 58629 62938
rect 58595 62594 58629 62628
rect 62768 62904 62802 62938
rect 62768 62594 62802 62628
rect 63585 62904 63619 62938
rect 63585 62594 63619 62628
rect 67758 62904 67792 62938
rect 67758 62594 67792 62628
rect 68575 62904 68609 62938
rect 68575 62594 68609 62628
rect 72748 62904 72782 62938
rect 72748 62594 72782 62628
rect 73565 62904 73599 62938
rect 73565 62594 73599 62628
rect 77738 62904 77772 62938
rect 77738 62594 77772 62628
rect 78555 62904 78589 62938
rect 78555 62594 78589 62628
rect 2888 61194 2922 61228
rect 2888 60884 2922 60918
rect 3705 61194 3739 61228
rect 3705 60884 3739 60918
rect 7878 61194 7912 61228
rect 7878 60884 7912 60918
rect 8695 61194 8729 61228
rect 8695 60884 8729 60918
rect 12868 61194 12902 61228
rect 12868 60884 12902 60918
rect 13685 61194 13719 61228
rect 13685 60884 13719 60918
rect 17858 61194 17892 61228
rect 17858 60884 17892 60918
rect 18675 61194 18709 61228
rect 18675 60884 18709 60918
rect 22848 61194 22882 61228
rect 22848 60884 22882 60918
rect 23665 61194 23699 61228
rect 23665 60884 23699 60918
rect 27838 61194 27872 61228
rect 27838 60884 27872 60918
rect 28655 61194 28689 61228
rect 28655 60884 28689 60918
rect 32828 61194 32862 61228
rect 32828 60884 32862 60918
rect 33645 61194 33679 61228
rect 33645 60884 33679 60918
rect 37818 61194 37852 61228
rect 37818 60884 37852 60918
rect 38635 61194 38669 61228
rect 38635 60884 38669 60918
rect 42808 61194 42842 61228
rect 42808 60884 42842 60918
rect 43625 61194 43659 61228
rect 43625 60884 43659 60918
rect 47798 61194 47832 61228
rect 47798 60884 47832 60918
rect 48615 61194 48649 61228
rect 48615 60884 48649 60918
rect 52788 61194 52822 61228
rect 52788 60884 52822 60918
rect 53605 61194 53639 61228
rect 53605 60884 53639 60918
rect 57778 61194 57812 61228
rect 57778 60884 57812 60918
rect 58595 61194 58629 61228
rect 58595 60884 58629 60918
rect 62768 61194 62802 61228
rect 62768 60884 62802 60918
rect 63585 61194 63619 61228
rect 63585 60884 63619 60918
rect 67758 61194 67792 61228
rect 67758 60884 67792 60918
rect 68575 61194 68609 61228
rect 68575 60884 68609 60918
rect 72748 61194 72782 61228
rect 72748 60884 72782 60918
rect 73565 61194 73599 61228
rect 73565 60884 73599 60918
rect 77738 61194 77772 61228
rect 77738 60884 77772 60918
rect 78555 61194 78589 61228
rect 78555 60884 78589 60918
rect 2888 59484 2922 59518
rect 2888 59174 2922 59208
rect 3705 59484 3739 59518
rect 3705 59174 3739 59208
rect 7878 59484 7912 59518
rect 7878 59174 7912 59208
rect 8695 59484 8729 59518
rect 8695 59174 8729 59208
rect 12868 59484 12902 59518
rect 12868 59174 12902 59208
rect 13685 59484 13719 59518
rect 13685 59174 13719 59208
rect 17858 59484 17892 59518
rect 17858 59174 17892 59208
rect 18675 59484 18709 59518
rect 18675 59174 18709 59208
rect 22848 59484 22882 59518
rect 22848 59174 22882 59208
rect 23665 59484 23699 59518
rect 23665 59174 23699 59208
rect 27838 59484 27872 59518
rect 27838 59174 27872 59208
rect 28655 59484 28689 59518
rect 28655 59174 28689 59208
rect 32828 59484 32862 59518
rect 32828 59174 32862 59208
rect 33645 59484 33679 59518
rect 33645 59174 33679 59208
rect 37818 59484 37852 59518
rect 37818 59174 37852 59208
rect 38635 59484 38669 59518
rect 38635 59174 38669 59208
rect 42808 59484 42842 59518
rect 42808 59174 42842 59208
rect 43625 59484 43659 59518
rect 43625 59174 43659 59208
rect 47798 59484 47832 59518
rect 47798 59174 47832 59208
rect 48615 59484 48649 59518
rect 48615 59174 48649 59208
rect 52788 59484 52822 59518
rect 52788 59174 52822 59208
rect 53605 59484 53639 59518
rect 53605 59174 53639 59208
rect 57778 59484 57812 59518
rect 57778 59174 57812 59208
rect 58595 59484 58629 59518
rect 58595 59174 58629 59208
rect 62768 59484 62802 59518
rect 62768 59174 62802 59208
rect 63585 59484 63619 59518
rect 63585 59174 63619 59208
rect 67758 59484 67792 59518
rect 67758 59174 67792 59208
rect 68575 59484 68609 59518
rect 68575 59174 68609 59208
rect 72748 59484 72782 59518
rect 72748 59174 72782 59208
rect 73565 59484 73599 59518
rect 73565 59174 73599 59208
rect 77738 59484 77772 59518
rect 77738 59174 77772 59208
rect 78555 59484 78589 59518
rect 78555 59174 78589 59208
rect 2888 57774 2922 57808
rect 2888 57464 2922 57498
rect 3705 57774 3739 57808
rect 3705 57464 3739 57498
rect 7878 57774 7912 57808
rect 7878 57464 7912 57498
rect 8695 57774 8729 57808
rect 8695 57464 8729 57498
rect 12868 57774 12902 57808
rect 12868 57464 12902 57498
rect 13685 57774 13719 57808
rect 13685 57464 13719 57498
rect 17858 57774 17892 57808
rect 17858 57464 17892 57498
rect 18675 57774 18709 57808
rect 18675 57464 18709 57498
rect 22848 57774 22882 57808
rect 22848 57464 22882 57498
rect 23665 57774 23699 57808
rect 23665 57464 23699 57498
rect 27838 57774 27872 57808
rect 27838 57464 27872 57498
rect 28655 57774 28689 57808
rect 28655 57464 28689 57498
rect 32828 57774 32862 57808
rect 32828 57464 32862 57498
rect 33645 57774 33679 57808
rect 33645 57464 33679 57498
rect 37818 57774 37852 57808
rect 37818 57464 37852 57498
rect 38635 57774 38669 57808
rect 38635 57464 38669 57498
rect 42808 57774 42842 57808
rect 42808 57464 42842 57498
rect 43625 57774 43659 57808
rect 43625 57464 43659 57498
rect 47798 57774 47832 57808
rect 47798 57464 47832 57498
rect 48615 57774 48649 57808
rect 48615 57464 48649 57498
rect 52788 57774 52822 57808
rect 52788 57464 52822 57498
rect 53605 57774 53639 57808
rect 53605 57464 53639 57498
rect 57778 57774 57812 57808
rect 57778 57464 57812 57498
rect 58595 57774 58629 57808
rect 58595 57464 58629 57498
rect 62768 57774 62802 57808
rect 62768 57464 62802 57498
rect 63585 57774 63619 57808
rect 63585 57464 63619 57498
rect 67758 57774 67792 57808
rect 67758 57464 67792 57498
rect 68575 57774 68609 57808
rect 68575 57464 68609 57498
rect 72748 57774 72782 57808
rect 72748 57464 72782 57498
rect 73565 57774 73599 57808
rect 73565 57464 73599 57498
rect 77738 57774 77772 57808
rect 77738 57464 77772 57498
rect 78555 57774 78589 57808
rect 78555 57464 78589 57498
rect 2888 56064 2922 56098
rect 2888 55754 2922 55788
rect 3705 56064 3739 56098
rect 3705 55754 3739 55788
rect 7878 56064 7912 56098
rect 7878 55754 7912 55788
rect 8695 56064 8729 56098
rect 8695 55754 8729 55788
rect 12868 56064 12902 56098
rect 12868 55754 12902 55788
rect 13685 56064 13719 56098
rect 13685 55754 13719 55788
rect 17858 56064 17892 56098
rect 17858 55754 17892 55788
rect 18675 56064 18709 56098
rect 18675 55754 18709 55788
rect 22848 56064 22882 56098
rect 22848 55754 22882 55788
rect 23665 56064 23699 56098
rect 23665 55754 23699 55788
rect 27838 56064 27872 56098
rect 27838 55754 27872 55788
rect 28655 56064 28689 56098
rect 28655 55754 28689 55788
rect 32828 56064 32862 56098
rect 32828 55754 32862 55788
rect 33645 56064 33679 56098
rect 33645 55754 33679 55788
rect 37818 56064 37852 56098
rect 37818 55754 37852 55788
rect 38635 56064 38669 56098
rect 38635 55754 38669 55788
rect 42808 56064 42842 56098
rect 42808 55754 42842 55788
rect 43625 56064 43659 56098
rect 43625 55754 43659 55788
rect 47798 56064 47832 56098
rect 47798 55754 47832 55788
rect 48615 56064 48649 56098
rect 48615 55754 48649 55788
rect 52788 56064 52822 56098
rect 52788 55754 52822 55788
rect 53605 56064 53639 56098
rect 53605 55754 53639 55788
rect 57778 56064 57812 56098
rect 57778 55754 57812 55788
rect 58595 56064 58629 56098
rect 58595 55754 58629 55788
rect 62768 56064 62802 56098
rect 62768 55754 62802 55788
rect 63585 56064 63619 56098
rect 63585 55754 63619 55788
rect 67758 56064 67792 56098
rect 67758 55754 67792 55788
rect 68575 56064 68609 56098
rect 68575 55754 68609 55788
rect 72748 56064 72782 56098
rect 72748 55754 72782 55788
rect 73565 56064 73599 56098
rect 73565 55754 73599 55788
rect 77738 56064 77772 56098
rect 77738 55754 77772 55788
rect 78555 56064 78589 56098
rect 78555 55754 78589 55788
rect 2888 54354 2922 54388
rect 2888 54044 2922 54078
rect 3705 54354 3739 54388
rect 3705 54044 3739 54078
rect 7878 54354 7912 54388
rect 7878 54044 7912 54078
rect 8695 54354 8729 54388
rect 8695 54044 8729 54078
rect 12868 54354 12902 54388
rect 12868 54044 12902 54078
rect 13685 54354 13719 54388
rect 13685 54044 13719 54078
rect 17858 54354 17892 54388
rect 17858 54044 17892 54078
rect 18675 54354 18709 54388
rect 18675 54044 18709 54078
rect 22848 54354 22882 54388
rect 22848 54044 22882 54078
rect 23665 54354 23699 54388
rect 23665 54044 23699 54078
rect 27838 54354 27872 54388
rect 27838 54044 27872 54078
rect 28655 54354 28689 54388
rect 28655 54044 28689 54078
rect 32828 54354 32862 54388
rect 32828 54044 32862 54078
rect 33645 54354 33679 54388
rect 33645 54044 33679 54078
rect 37818 54354 37852 54388
rect 37818 54044 37852 54078
rect 38635 54354 38669 54388
rect 38635 54044 38669 54078
rect 42808 54354 42842 54388
rect 42808 54044 42842 54078
rect 43625 54354 43659 54388
rect 43625 54044 43659 54078
rect 47798 54354 47832 54388
rect 47798 54044 47832 54078
rect 48615 54354 48649 54388
rect 48615 54044 48649 54078
rect 52788 54354 52822 54388
rect 52788 54044 52822 54078
rect 53605 54354 53639 54388
rect 53605 54044 53639 54078
rect 57778 54354 57812 54388
rect 57778 54044 57812 54078
rect 58595 54354 58629 54388
rect 58595 54044 58629 54078
rect 62768 54354 62802 54388
rect 62768 54044 62802 54078
rect 63585 54354 63619 54388
rect 63585 54044 63619 54078
rect 67758 54354 67792 54388
rect 67758 54044 67792 54078
rect 68575 54354 68609 54388
rect 68575 54044 68609 54078
rect 72748 54354 72782 54388
rect 72748 54044 72782 54078
rect 73565 54354 73599 54388
rect 73565 54044 73599 54078
rect 77738 54354 77772 54388
rect 77738 54044 77772 54078
rect 78555 54354 78589 54388
rect 78555 54044 78589 54078
rect 2888 52644 2922 52678
rect 2888 52334 2922 52368
rect 3705 52644 3739 52678
rect 3705 52334 3739 52368
rect 7878 52644 7912 52678
rect 7878 52334 7912 52368
rect 8695 52644 8729 52678
rect 8695 52334 8729 52368
rect 12868 52644 12902 52678
rect 12868 52334 12902 52368
rect 13685 52644 13719 52678
rect 13685 52334 13719 52368
rect 17858 52644 17892 52678
rect 17858 52334 17892 52368
rect 18675 52644 18709 52678
rect 18675 52334 18709 52368
rect 22848 52644 22882 52678
rect 22848 52334 22882 52368
rect 23665 52644 23699 52678
rect 23665 52334 23699 52368
rect 27838 52644 27872 52678
rect 27838 52334 27872 52368
rect 28655 52644 28689 52678
rect 28655 52334 28689 52368
rect 32828 52644 32862 52678
rect 32828 52334 32862 52368
rect 33645 52644 33679 52678
rect 33645 52334 33679 52368
rect 37818 52644 37852 52678
rect 37818 52334 37852 52368
rect 38635 52644 38669 52678
rect 38635 52334 38669 52368
rect 42808 52644 42842 52678
rect 42808 52334 42842 52368
rect 43625 52644 43659 52678
rect 43625 52334 43659 52368
rect 47798 52644 47832 52678
rect 47798 52334 47832 52368
rect 48615 52644 48649 52678
rect 48615 52334 48649 52368
rect 52788 52644 52822 52678
rect 52788 52334 52822 52368
rect 53605 52644 53639 52678
rect 53605 52334 53639 52368
rect 57778 52644 57812 52678
rect 57778 52334 57812 52368
rect 58595 52644 58629 52678
rect 58595 52334 58629 52368
rect 62768 52644 62802 52678
rect 62768 52334 62802 52368
rect 63585 52644 63619 52678
rect 63585 52334 63619 52368
rect 67758 52644 67792 52678
rect 67758 52334 67792 52368
rect 68575 52644 68609 52678
rect 68575 52334 68609 52368
rect 72748 52644 72782 52678
rect 72748 52334 72782 52368
rect 73565 52644 73599 52678
rect 73565 52334 73599 52368
rect 77738 52644 77772 52678
rect 77738 52334 77772 52368
rect 78555 52644 78589 52678
rect 78555 52334 78589 52368
rect 2888 50934 2922 50968
rect 2888 50624 2922 50658
rect 3705 50934 3739 50968
rect 3705 50624 3739 50658
rect 7878 50934 7912 50968
rect 7878 50624 7912 50658
rect 8695 50934 8729 50968
rect 8695 50624 8729 50658
rect 12868 50934 12902 50968
rect 12868 50624 12902 50658
rect 13685 50934 13719 50968
rect 13685 50624 13719 50658
rect 17858 50934 17892 50968
rect 17858 50624 17892 50658
rect 18675 50934 18709 50968
rect 18675 50624 18709 50658
rect 22848 50934 22882 50968
rect 22848 50624 22882 50658
rect 23665 50934 23699 50968
rect 23665 50624 23699 50658
rect 27838 50934 27872 50968
rect 27838 50624 27872 50658
rect 28655 50934 28689 50968
rect 28655 50624 28689 50658
rect 32828 50934 32862 50968
rect 32828 50624 32862 50658
rect 33645 50934 33679 50968
rect 33645 50624 33679 50658
rect 37818 50934 37852 50968
rect 37818 50624 37852 50658
rect 38635 50934 38669 50968
rect 38635 50624 38669 50658
rect 42808 50934 42842 50968
rect 42808 50624 42842 50658
rect 43625 50934 43659 50968
rect 43625 50624 43659 50658
rect 47798 50934 47832 50968
rect 47798 50624 47832 50658
rect 48615 50934 48649 50968
rect 48615 50624 48649 50658
rect 52788 50934 52822 50968
rect 52788 50624 52822 50658
rect 53605 50934 53639 50968
rect 53605 50624 53639 50658
rect 57778 50934 57812 50968
rect 57778 50624 57812 50658
rect 58595 50934 58629 50968
rect 58595 50624 58629 50658
rect 62768 50934 62802 50968
rect 62768 50624 62802 50658
rect 63585 50934 63619 50968
rect 63585 50624 63619 50658
rect 67758 50934 67792 50968
rect 67758 50624 67792 50658
rect 68575 50934 68609 50968
rect 68575 50624 68609 50658
rect 72748 50934 72782 50968
rect 72748 50624 72782 50658
rect 73565 50934 73599 50968
rect 73565 50624 73599 50658
rect 77738 50934 77772 50968
rect 77738 50624 77772 50658
rect 78555 50934 78589 50968
rect 78555 50624 78589 50658
rect 2888 49224 2922 49258
rect 2888 48914 2922 48948
rect 3705 49224 3739 49258
rect 3705 48914 3739 48948
rect 7878 49224 7912 49258
rect 7878 48914 7912 48948
rect 8695 49224 8729 49258
rect 8695 48914 8729 48948
rect 12868 49224 12902 49258
rect 12868 48914 12902 48948
rect 13685 49224 13719 49258
rect 13685 48914 13719 48948
rect 17858 49224 17892 49258
rect 17858 48914 17892 48948
rect 18675 49224 18709 49258
rect 18675 48914 18709 48948
rect 22848 49224 22882 49258
rect 22848 48914 22882 48948
rect 23665 49224 23699 49258
rect 23665 48914 23699 48948
rect 27838 49224 27872 49258
rect 27838 48914 27872 48948
rect 28655 49224 28689 49258
rect 28655 48914 28689 48948
rect 32828 49224 32862 49258
rect 32828 48914 32862 48948
rect 33645 49224 33679 49258
rect 33645 48914 33679 48948
rect 37818 49224 37852 49258
rect 37818 48914 37852 48948
rect 38635 49224 38669 49258
rect 38635 48914 38669 48948
rect 42808 49224 42842 49258
rect 42808 48914 42842 48948
rect 43625 49224 43659 49258
rect 43625 48914 43659 48948
rect 47798 49224 47832 49258
rect 47798 48914 47832 48948
rect 48615 49224 48649 49258
rect 48615 48914 48649 48948
rect 52788 49224 52822 49258
rect 52788 48914 52822 48948
rect 53605 49224 53639 49258
rect 53605 48914 53639 48948
rect 57778 49224 57812 49258
rect 57778 48914 57812 48948
rect 58595 49224 58629 49258
rect 58595 48914 58629 48948
rect 62768 49224 62802 49258
rect 62768 48914 62802 48948
rect 63585 49224 63619 49258
rect 63585 48914 63619 48948
rect 67758 49224 67792 49258
rect 67758 48914 67792 48948
rect 68575 49224 68609 49258
rect 68575 48914 68609 48948
rect 72748 49224 72782 49258
rect 72748 48914 72782 48948
rect 73565 49224 73599 49258
rect 73565 48914 73599 48948
rect 77738 49224 77772 49258
rect 77738 48914 77772 48948
rect 78555 49224 78589 49258
rect 78555 48914 78589 48948
rect 2888 47514 2922 47548
rect 2888 47204 2922 47238
rect 3705 47514 3739 47548
rect 3705 47204 3739 47238
rect 7878 47514 7912 47548
rect 7878 47204 7912 47238
rect 8695 47514 8729 47548
rect 8695 47204 8729 47238
rect 12868 47514 12902 47548
rect 12868 47204 12902 47238
rect 13685 47514 13719 47548
rect 13685 47204 13719 47238
rect 17858 47514 17892 47548
rect 17858 47204 17892 47238
rect 18675 47514 18709 47548
rect 18675 47204 18709 47238
rect 22848 47514 22882 47548
rect 22848 47204 22882 47238
rect 23665 47514 23699 47548
rect 23665 47204 23699 47238
rect 27838 47514 27872 47548
rect 27838 47204 27872 47238
rect 28655 47514 28689 47548
rect 28655 47204 28689 47238
rect 32828 47514 32862 47548
rect 32828 47204 32862 47238
rect 33645 47514 33679 47548
rect 33645 47204 33679 47238
rect 37818 47514 37852 47548
rect 37818 47204 37852 47238
rect 38635 47514 38669 47548
rect 38635 47204 38669 47238
rect 42808 47514 42842 47548
rect 42808 47204 42842 47238
rect 43625 47514 43659 47548
rect 43625 47204 43659 47238
rect 47798 47514 47832 47548
rect 47798 47204 47832 47238
rect 48615 47514 48649 47548
rect 48615 47204 48649 47238
rect 52788 47514 52822 47548
rect 52788 47204 52822 47238
rect 53605 47514 53639 47548
rect 53605 47204 53639 47238
rect 57778 47514 57812 47548
rect 57778 47204 57812 47238
rect 58595 47514 58629 47548
rect 58595 47204 58629 47238
rect 62768 47514 62802 47548
rect 62768 47204 62802 47238
rect 63585 47514 63619 47548
rect 63585 47204 63619 47238
rect 67758 47514 67792 47548
rect 67758 47204 67792 47238
rect 68575 47514 68609 47548
rect 68575 47204 68609 47238
rect 72748 47514 72782 47548
rect 72748 47204 72782 47238
rect 73565 47514 73599 47548
rect 73565 47204 73599 47238
rect 77738 47514 77772 47548
rect 77738 47204 77772 47238
rect 78555 47514 78589 47548
rect 78555 47204 78589 47238
rect 2888 45804 2922 45838
rect 2888 45494 2922 45528
rect 3705 45804 3739 45838
rect 3705 45494 3739 45528
rect 7878 45804 7912 45838
rect 7878 45494 7912 45528
rect 8695 45804 8729 45838
rect 8695 45494 8729 45528
rect 12868 45804 12902 45838
rect 12868 45494 12902 45528
rect 13685 45804 13719 45838
rect 13685 45494 13719 45528
rect 17858 45804 17892 45838
rect 17858 45494 17892 45528
rect 18675 45804 18709 45838
rect 18675 45494 18709 45528
rect 22848 45804 22882 45838
rect 22848 45494 22882 45528
rect 23665 45804 23699 45838
rect 23665 45494 23699 45528
rect 27838 45804 27872 45838
rect 27838 45494 27872 45528
rect 28655 45804 28689 45838
rect 28655 45494 28689 45528
rect 32828 45804 32862 45838
rect 32828 45494 32862 45528
rect 33645 45804 33679 45838
rect 33645 45494 33679 45528
rect 37818 45804 37852 45838
rect 37818 45494 37852 45528
rect 38635 45804 38669 45838
rect 38635 45494 38669 45528
rect 42808 45804 42842 45838
rect 42808 45494 42842 45528
rect 43625 45804 43659 45838
rect 43625 45494 43659 45528
rect 47798 45804 47832 45838
rect 47798 45494 47832 45528
rect 48615 45804 48649 45838
rect 48615 45494 48649 45528
rect 52788 45804 52822 45838
rect 52788 45494 52822 45528
rect 53605 45804 53639 45838
rect 53605 45494 53639 45528
rect 57778 45804 57812 45838
rect 57778 45494 57812 45528
rect 58595 45804 58629 45838
rect 58595 45494 58629 45528
rect 62768 45804 62802 45838
rect 62768 45494 62802 45528
rect 63585 45804 63619 45838
rect 63585 45494 63619 45528
rect 67758 45804 67792 45838
rect 67758 45494 67792 45528
rect 68575 45804 68609 45838
rect 68575 45494 68609 45528
rect 72748 45804 72782 45838
rect 72748 45494 72782 45528
rect 73565 45804 73599 45838
rect 73565 45494 73599 45528
rect 77738 45804 77772 45838
rect 77738 45494 77772 45528
rect 78555 45804 78589 45838
rect 78555 45494 78589 45528
rect 2888 44094 2922 44128
rect 2888 43784 2922 43818
rect 3705 44094 3739 44128
rect 3705 43784 3739 43818
rect 7878 44094 7912 44128
rect 7878 43784 7912 43818
rect 8695 44094 8729 44128
rect 8695 43784 8729 43818
rect 12868 44094 12902 44128
rect 12868 43784 12902 43818
rect 13685 44094 13719 44128
rect 13685 43784 13719 43818
rect 17858 44094 17892 44128
rect 17858 43784 17892 43818
rect 18675 44094 18709 44128
rect 18675 43784 18709 43818
rect 22848 44094 22882 44128
rect 22848 43784 22882 43818
rect 23665 44094 23699 44128
rect 23665 43784 23699 43818
rect 27838 44094 27872 44128
rect 27838 43784 27872 43818
rect 28655 44094 28689 44128
rect 28655 43784 28689 43818
rect 32828 44094 32862 44128
rect 32828 43784 32862 43818
rect 33645 44094 33679 44128
rect 33645 43784 33679 43818
rect 37818 44094 37852 44128
rect 37818 43784 37852 43818
rect 38635 44094 38669 44128
rect 38635 43784 38669 43818
rect 42808 44094 42842 44128
rect 42808 43784 42842 43818
rect 43625 44094 43659 44128
rect 43625 43784 43659 43818
rect 47798 44094 47832 44128
rect 47798 43784 47832 43818
rect 48615 44094 48649 44128
rect 48615 43784 48649 43818
rect 52788 44094 52822 44128
rect 52788 43784 52822 43818
rect 53605 44094 53639 44128
rect 53605 43784 53639 43818
rect 57778 44094 57812 44128
rect 57778 43784 57812 43818
rect 58595 44094 58629 44128
rect 58595 43784 58629 43818
rect 62768 44094 62802 44128
rect 62768 43784 62802 43818
rect 63585 44094 63619 44128
rect 63585 43784 63619 43818
rect 67758 44094 67792 44128
rect 67758 43784 67792 43818
rect 68575 44094 68609 44128
rect 68575 43784 68609 43818
rect 72748 44094 72782 44128
rect 72748 43784 72782 43818
rect 73565 44094 73599 44128
rect 73565 43784 73599 43818
rect 77738 44094 77772 44128
rect 77738 43784 77772 43818
rect 78555 44094 78589 44128
rect 78555 43784 78589 43818
rect 2888 42384 2922 42418
rect 2888 42074 2922 42108
rect 3705 42384 3739 42418
rect 3705 42074 3739 42108
rect 7878 42384 7912 42418
rect 7878 42074 7912 42108
rect 8695 42384 8729 42418
rect 8695 42074 8729 42108
rect 12868 42384 12902 42418
rect 12868 42074 12902 42108
rect 13685 42384 13719 42418
rect 13685 42074 13719 42108
rect 17858 42384 17892 42418
rect 17858 42074 17892 42108
rect 18675 42384 18709 42418
rect 18675 42074 18709 42108
rect 22848 42384 22882 42418
rect 22848 42074 22882 42108
rect 23665 42384 23699 42418
rect 23665 42074 23699 42108
rect 27838 42384 27872 42418
rect 27838 42074 27872 42108
rect 28655 42384 28689 42418
rect 28655 42074 28689 42108
rect 32828 42384 32862 42418
rect 32828 42074 32862 42108
rect 33645 42384 33679 42418
rect 33645 42074 33679 42108
rect 37818 42384 37852 42418
rect 37818 42074 37852 42108
rect 38635 42384 38669 42418
rect 38635 42074 38669 42108
rect 42808 42384 42842 42418
rect 42808 42074 42842 42108
rect 43625 42384 43659 42418
rect 43625 42074 43659 42108
rect 47798 42384 47832 42418
rect 47798 42074 47832 42108
rect 48615 42384 48649 42418
rect 48615 42074 48649 42108
rect 52788 42384 52822 42418
rect 52788 42074 52822 42108
rect 53605 42384 53639 42418
rect 53605 42074 53639 42108
rect 57778 42384 57812 42418
rect 57778 42074 57812 42108
rect 58595 42384 58629 42418
rect 58595 42074 58629 42108
rect 62768 42384 62802 42418
rect 62768 42074 62802 42108
rect 63585 42384 63619 42418
rect 63585 42074 63619 42108
rect 67758 42384 67792 42418
rect 67758 42074 67792 42108
rect 68575 42384 68609 42418
rect 68575 42074 68609 42108
rect 72748 42384 72782 42418
rect 72748 42074 72782 42108
rect 73565 42384 73599 42418
rect 73565 42074 73599 42108
rect 77738 42384 77772 42418
rect 77738 42074 77772 42108
rect 78555 42384 78589 42418
rect 78555 42074 78589 42108
rect 2888 40674 2922 40708
rect 2888 40364 2922 40398
rect 3705 40674 3739 40708
rect 3705 40364 3739 40398
rect 7878 40674 7912 40708
rect 7878 40364 7912 40398
rect 8695 40674 8729 40708
rect 8695 40364 8729 40398
rect 12868 40674 12902 40708
rect 12868 40364 12902 40398
rect 13685 40674 13719 40708
rect 13685 40364 13719 40398
rect 17858 40674 17892 40708
rect 17858 40364 17892 40398
rect 18675 40674 18709 40708
rect 18675 40364 18709 40398
rect 22848 40674 22882 40708
rect 22848 40364 22882 40398
rect 23665 40674 23699 40708
rect 23665 40364 23699 40398
rect 27838 40674 27872 40708
rect 27838 40364 27872 40398
rect 28655 40674 28689 40708
rect 28655 40364 28689 40398
rect 32828 40674 32862 40708
rect 32828 40364 32862 40398
rect 33645 40674 33679 40708
rect 33645 40364 33679 40398
rect 37818 40674 37852 40708
rect 37818 40364 37852 40398
rect 38635 40674 38669 40708
rect 38635 40364 38669 40398
rect 42808 40674 42842 40708
rect 42808 40364 42842 40398
rect 43625 40674 43659 40708
rect 43625 40364 43659 40398
rect 47798 40674 47832 40708
rect 47798 40364 47832 40398
rect 48615 40674 48649 40708
rect 48615 40364 48649 40398
rect 52788 40674 52822 40708
rect 52788 40364 52822 40398
rect 53605 40674 53639 40708
rect 53605 40364 53639 40398
rect 57778 40674 57812 40708
rect 57778 40364 57812 40398
rect 58595 40674 58629 40708
rect 58595 40364 58629 40398
rect 62768 40674 62802 40708
rect 62768 40364 62802 40398
rect 63585 40674 63619 40708
rect 63585 40364 63619 40398
rect 67758 40674 67792 40708
rect 67758 40364 67792 40398
rect 68575 40674 68609 40708
rect 68575 40364 68609 40398
rect 72748 40674 72782 40708
rect 72748 40364 72782 40398
rect 73565 40674 73599 40708
rect 73565 40364 73599 40398
rect 77738 40674 77772 40708
rect 77738 40364 77772 40398
rect 78555 40674 78589 40708
rect 78555 40364 78589 40398
<< locali >>
rect 2740 66470 2830 66590
rect 2740 66210 2760 66470
rect 2800 66420 2830 66470
rect 2820 66262 2830 66420
rect 3800 66470 3890 66590
rect 3800 66420 3830 66470
rect 2888 66358 2922 66374
rect 2956 66368 2972 66402
rect 3148 66368 3164 66402
rect 3454 66368 3470 66402
rect 3646 66368 3662 66402
rect 2888 66308 2922 66324
rect 3705 66358 3739 66374
rect 2956 66280 2972 66314
rect 3148 66280 3164 66314
rect 3454 66280 3470 66314
rect 3646 66280 3662 66314
rect 3705 66308 3739 66324
rect 2800 66210 2830 66262
rect 2740 66150 2830 66210
rect 2740 65910 2760 66150
rect 2800 66110 2830 66150
rect 2820 65952 2830 66110
rect 3800 66262 3808 66420
rect 3800 66230 3830 66262
rect 3870 66230 3890 66470
rect 3800 66150 3890 66230
rect 3800 66110 3830 66150
rect 2888 66048 2922 66064
rect 2956 66058 2972 66092
rect 3148 66058 3164 66092
rect 3454 66058 3470 66092
rect 3646 66058 3662 66092
rect 2888 65998 2922 66014
rect 3705 66048 3739 66064
rect 2956 65970 2972 66004
rect 3148 65970 3164 66004
rect 3454 65970 3470 66004
rect 3646 65970 3662 66004
rect 3705 65998 3739 66014
rect 2800 65910 2830 65952
rect 2740 65780 2830 65910
rect 3800 65952 3808 66110
rect 3800 65910 3830 65952
rect 3870 65910 3890 66150
rect 3800 65780 3890 65910
rect 7730 66470 7820 66590
rect 7730 66210 7750 66470
rect 7790 66420 7820 66470
rect 7810 66262 7820 66420
rect 8790 66470 8880 66590
rect 8790 66420 8820 66470
rect 7878 66358 7912 66374
rect 7946 66368 7962 66402
rect 8138 66368 8154 66402
rect 8444 66368 8460 66402
rect 8636 66368 8652 66402
rect 7878 66308 7912 66324
rect 8695 66358 8729 66374
rect 7946 66280 7962 66314
rect 8138 66280 8154 66314
rect 8444 66280 8460 66314
rect 8636 66280 8652 66314
rect 8695 66308 8729 66324
rect 7790 66210 7820 66262
rect 7730 66150 7820 66210
rect 7730 65910 7750 66150
rect 7790 66110 7820 66150
rect 7810 65952 7820 66110
rect 8790 66262 8798 66420
rect 8790 66230 8820 66262
rect 8860 66230 8880 66470
rect 8790 66150 8880 66230
rect 8790 66110 8820 66150
rect 7878 66048 7912 66064
rect 7946 66058 7962 66092
rect 8138 66058 8154 66092
rect 8444 66058 8460 66092
rect 8636 66058 8652 66092
rect 7878 65998 7912 66014
rect 8695 66048 8729 66064
rect 7946 65970 7962 66004
rect 8138 65970 8154 66004
rect 8444 65970 8460 66004
rect 8636 65970 8652 66004
rect 8695 65998 8729 66014
rect 7790 65910 7820 65952
rect 7730 65780 7820 65910
rect 8790 65952 8798 66110
rect 8790 65910 8820 65952
rect 8860 65910 8880 66150
rect 8790 65780 8880 65910
rect 12720 66470 12810 66590
rect 12720 66210 12740 66470
rect 12780 66420 12810 66470
rect 12800 66262 12810 66420
rect 13780 66470 13870 66590
rect 13780 66420 13810 66470
rect 12868 66358 12902 66374
rect 12936 66368 12952 66402
rect 13128 66368 13144 66402
rect 13434 66368 13450 66402
rect 13626 66368 13642 66402
rect 12868 66308 12902 66324
rect 13685 66358 13719 66374
rect 12936 66280 12952 66314
rect 13128 66280 13144 66314
rect 13434 66280 13450 66314
rect 13626 66280 13642 66314
rect 13685 66308 13719 66324
rect 12780 66210 12810 66262
rect 12720 66150 12810 66210
rect 12720 65910 12740 66150
rect 12780 66110 12810 66150
rect 12800 65952 12810 66110
rect 13780 66262 13788 66420
rect 13780 66230 13810 66262
rect 13850 66230 13870 66470
rect 13780 66150 13870 66230
rect 13780 66110 13810 66150
rect 12868 66048 12902 66064
rect 12936 66058 12952 66092
rect 13128 66058 13144 66092
rect 13434 66058 13450 66092
rect 13626 66058 13642 66092
rect 12868 65998 12902 66014
rect 13685 66048 13719 66064
rect 12936 65970 12952 66004
rect 13128 65970 13144 66004
rect 13434 65970 13450 66004
rect 13626 65970 13642 66004
rect 13685 65998 13719 66014
rect 12780 65910 12810 65952
rect 12720 65780 12810 65910
rect 13780 65952 13788 66110
rect 13780 65910 13810 65952
rect 13850 65910 13870 66150
rect 13780 65780 13870 65910
rect 17710 66470 17800 66590
rect 17710 66210 17730 66470
rect 17770 66420 17800 66470
rect 17790 66262 17800 66420
rect 18770 66470 18860 66590
rect 18770 66420 18800 66470
rect 17858 66358 17892 66374
rect 17926 66368 17942 66402
rect 18118 66368 18134 66402
rect 18424 66368 18440 66402
rect 18616 66368 18632 66402
rect 17858 66308 17892 66324
rect 18675 66358 18709 66374
rect 17926 66280 17942 66314
rect 18118 66280 18134 66314
rect 18424 66280 18440 66314
rect 18616 66280 18632 66314
rect 18675 66308 18709 66324
rect 17770 66210 17800 66262
rect 17710 66150 17800 66210
rect 17710 65910 17730 66150
rect 17770 66110 17800 66150
rect 17790 65952 17800 66110
rect 18770 66262 18778 66420
rect 18770 66230 18800 66262
rect 18840 66230 18860 66470
rect 18770 66150 18860 66230
rect 18770 66110 18800 66150
rect 17858 66048 17892 66064
rect 17926 66058 17942 66092
rect 18118 66058 18134 66092
rect 18424 66058 18440 66092
rect 18616 66058 18632 66092
rect 17858 65998 17892 66014
rect 18675 66048 18709 66064
rect 17926 65970 17942 66004
rect 18118 65970 18134 66004
rect 18424 65970 18440 66004
rect 18616 65970 18632 66004
rect 18675 65998 18709 66014
rect 17770 65910 17800 65952
rect 17710 65780 17800 65910
rect 18770 65952 18778 66110
rect 18770 65910 18800 65952
rect 18840 65910 18860 66150
rect 18770 65780 18860 65910
rect 22700 66470 22790 66590
rect 22700 66210 22720 66470
rect 22760 66420 22790 66470
rect 22780 66262 22790 66420
rect 23760 66470 23850 66590
rect 23760 66420 23790 66470
rect 22848 66358 22882 66374
rect 22916 66368 22932 66402
rect 23108 66368 23124 66402
rect 23414 66368 23430 66402
rect 23606 66368 23622 66402
rect 22848 66308 22882 66324
rect 23665 66358 23699 66374
rect 22916 66280 22932 66314
rect 23108 66280 23124 66314
rect 23414 66280 23430 66314
rect 23606 66280 23622 66314
rect 23665 66308 23699 66324
rect 22760 66210 22790 66262
rect 22700 66150 22790 66210
rect 22700 65910 22720 66150
rect 22760 66110 22790 66150
rect 22780 65952 22790 66110
rect 23760 66262 23768 66420
rect 23760 66230 23790 66262
rect 23830 66230 23850 66470
rect 23760 66150 23850 66230
rect 23760 66110 23790 66150
rect 22848 66048 22882 66064
rect 22916 66058 22932 66092
rect 23108 66058 23124 66092
rect 23414 66058 23430 66092
rect 23606 66058 23622 66092
rect 22848 65998 22882 66014
rect 23665 66048 23699 66064
rect 22916 65970 22932 66004
rect 23108 65970 23124 66004
rect 23414 65970 23430 66004
rect 23606 65970 23622 66004
rect 23665 65998 23699 66014
rect 22760 65910 22790 65952
rect 22700 65780 22790 65910
rect 23760 65952 23768 66110
rect 23760 65910 23790 65952
rect 23830 65910 23850 66150
rect 23760 65780 23850 65910
rect 27690 66470 27780 66590
rect 27690 66210 27710 66470
rect 27750 66420 27780 66470
rect 27770 66262 27780 66420
rect 28750 66470 28840 66590
rect 28750 66420 28780 66470
rect 27838 66358 27872 66374
rect 27906 66368 27922 66402
rect 28098 66368 28114 66402
rect 28404 66368 28420 66402
rect 28596 66368 28612 66402
rect 27838 66308 27872 66324
rect 28655 66358 28689 66374
rect 27906 66280 27922 66314
rect 28098 66280 28114 66314
rect 28404 66280 28420 66314
rect 28596 66280 28612 66314
rect 28655 66308 28689 66324
rect 27750 66210 27780 66262
rect 27690 66150 27780 66210
rect 27690 65910 27710 66150
rect 27750 66110 27780 66150
rect 27770 65952 27780 66110
rect 28750 66262 28758 66420
rect 28750 66230 28780 66262
rect 28820 66230 28840 66470
rect 28750 66150 28840 66230
rect 28750 66110 28780 66150
rect 27838 66048 27872 66064
rect 27906 66058 27922 66092
rect 28098 66058 28114 66092
rect 28404 66058 28420 66092
rect 28596 66058 28612 66092
rect 27838 65998 27872 66014
rect 28655 66048 28689 66064
rect 27906 65970 27922 66004
rect 28098 65970 28114 66004
rect 28404 65970 28420 66004
rect 28596 65970 28612 66004
rect 28655 65998 28689 66014
rect 27750 65910 27780 65952
rect 27690 65780 27780 65910
rect 28750 65952 28758 66110
rect 28750 65910 28780 65952
rect 28820 65910 28840 66150
rect 28750 65780 28840 65910
rect 32680 66470 32770 66590
rect 32680 66210 32700 66470
rect 32740 66420 32770 66470
rect 32760 66262 32770 66420
rect 33740 66470 33830 66590
rect 33740 66420 33770 66470
rect 32828 66358 32862 66374
rect 32896 66368 32912 66402
rect 33088 66368 33104 66402
rect 33394 66368 33410 66402
rect 33586 66368 33602 66402
rect 32828 66308 32862 66324
rect 33645 66358 33679 66374
rect 32896 66280 32912 66314
rect 33088 66280 33104 66314
rect 33394 66280 33410 66314
rect 33586 66280 33602 66314
rect 33645 66308 33679 66324
rect 32740 66210 32770 66262
rect 32680 66150 32770 66210
rect 32680 65910 32700 66150
rect 32740 66110 32770 66150
rect 32760 65952 32770 66110
rect 33740 66262 33748 66420
rect 33740 66230 33770 66262
rect 33810 66230 33830 66470
rect 33740 66150 33830 66230
rect 33740 66110 33770 66150
rect 32828 66048 32862 66064
rect 32896 66058 32912 66092
rect 33088 66058 33104 66092
rect 33394 66058 33410 66092
rect 33586 66058 33602 66092
rect 32828 65998 32862 66014
rect 33645 66048 33679 66064
rect 32896 65970 32912 66004
rect 33088 65970 33104 66004
rect 33394 65970 33410 66004
rect 33586 65970 33602 66004
rect 33645 65998 33679 66014
rect 32740 65910 32770 65952
rect 32680 65780 32770 65910
rect 33740 65952 33748 66110
rect 33740 65910 33770 65952
rect 33810 65910 33830 66150
rect 33740 65780 33830 65910
rect 37670 66470 37760 66590
rect 37670 66210 37690 66470
rect 37730 66420 37760 66470
rect 37750 66262 37760 66420
rect 38730 66470 38820 66590
rect 38730 66420 38760 66470
rect 37818 66358 37852 66374
rect 37886 66368 37902 66402
rect 38078 66368 38094 66402
rect 38384 66368 38400 66402
rect 38576 66368 38592 66402
rect 37818 66308 37852 66324
rect 38635 66358 38669 66374
rect 37886 66280 37902 66314
rect 38078 66280 38094 66314
rect 38384 66280 38400 66314
rect 38576 66280 38592 66314
rect 38635 66308 38669 66324
rect 37730 66210 37760 66262
rect 37670 66150 37760 66210
rect 37670 65910 37690 66150
rect 37730 66110 37760 66150
rect 37750 65952 37760 66110
rect 38730 66262 38738 66420
rect 38730 66230 38760 66262
rect 38800 66230 38820 66470
rect 38730 66150 38820 66230
rect 38730 66110 38760 66150
rect 37818 66048 37852 66064
rect 37886 66058 37902 66092
rect 38078 66058 38094 66092
rect 38384 66058 38400 66092
rect 38576 66058 38592 66092
rect 37818 65998 37852 66014
rect 38635 66048 38669 66064
rect 37886 65970 37902 66004
rect 38078 65970 38094 66004
rect 38384 65970 38400 66004
rect 38576 65970 38592 66004
rect 38635 65998 38669 66014
rect 37730 65910 37760 65952
rect 37670 65780 37760 65910
rect 38730 65952 38738 66110
rect 38730 65910 38760 65952
rect 38800 65910 38820 66150
rect 38730 65780 38820 65910
rect 42660 66470 42750 66590
rect 42660 66210 42680 66470
rect 42720 66420 42750 66470
rect 42740 66262 42750 66420
rect 43720 66470 43810 66590
rect 43720 66420 43750 66470
rect 42808 66358 42842 66374
rect 42876 66368 42892 66402
rect 43068 66368 43084 66402
rect 43374 66368 43390 66402
rect 43566 66368 43582 66402
rect 42808 66308 42842 66324
rect 43625 66358 43659 66374
rect 42876 66280 42892 66314
rect 43068 66280 43084 66314
rect 43374 66280 43390 66314
rect 43566 66280 43582 66314
rect 43625 66308 43659 66324
rect 42720 66210 42750 66262
rect 42660 66150 42750 66210
rect 42660 65910 42680 66150
rect 42720 66110 42750 66150
rect 42740 65952 42750 66110
rect 43720 66262 43728 66420
rect 43720 66230 43750 66262
rect 43790 66230 43810 66470
rect 43720 66150 43810 66230
rect 43720 66110 43750 66150
rect 42808 66048 42842 66064
rect 42876 66058 42892 66092
rect 43068 66058 43084 66092
rect 43374 66058 43390 66092
rect 43566 66058 43582 66092
rect 42808 65998 42842 66014
rect 43625 66048 43659 66064
rect 42876 65970 42892 66004
rect 43068 65970 43084 66004
rect 43374 65970 43390 66004
rect 43566 65970 43582 66004
rect 43625 65998 43659 66014
rect 42720 65910 42750 65952
rect 42660 65780 42750 65910
rect 43720 65952 43728 66110
rect 43720 65910 43750 65952
rect 43790 65910 43810 66150
rect 43720 65780 43810 65910
rect 47650 66470 47740 66590
rect 47650 66210 47670 66470
rect 47710 66420 47740 66470
rect 47730 66262 47740 66420
rect 48710 66470 48800 66590
rect 48710 66420 48740 66470
rect 47798 66358 47832 66374
rect 47866 66368 47882 66402
rect 48058 66368 48074 66402
rect 48364 66368 48380 66402
rect 48556 66368 48572 66402
rect 47798 66308 47832 66324
rect 48615 66358 48649 66374
rect 47866 66280 47882 66314
rect 48058 66280 48074 66314
rect 48364 66280 48380 66314
rect 48556 66280 48572 66314
rect 48615 66308 48649 66324
rect 47710 66210 47740 66262
rect 47650 66150 47740 66210
rect 47650 65910 47670 66150
rect 47710 66110 47740 66150
rect 47730 65952 47740 66110
rect 48710 66262 48718 66420
rect 48710 66230 48740 66262
rect 48780 66230 48800 66470
rect 48710 66150 48800 66230
rect 48710 66110 48740 66150
rect 47798 66048 47832 66064
rect 47866 66058 47882 66092
rect 48058 66058 48074 66092
rect 48364 66058 48380 66092
rect 48556 66058 48572 66092
rect 47798 65998 47832 66014
rect 48615 66048 48649 66064
rect 47866 65970 47882 66004
rect 48058 65970 48074 66004
rect 48364 65970 48380 66004
rect 48556 65970 48572 66004
rect 48615 65998 48649 66014
rect 47710 65910 47740 65952
rect 47650 65780 47740 65910
rect 48710 65952 48718 66110
rect 48710 65910 48740 65952
rect 48780 65910 48800 66150
rect 48710 65780 48800 65910
rect 52640 66470 52730 66590
rect 52640 66210 52660 66470
rect 52700 66420 52730 66470
rect 52720 66262 52730 66420
rect 53700 66470 53790 66590
rect 53700 66420 53730 66470
rect 52788 66358 52822 66374
rect 52856 66368 52872 66402
rect 53048 66368 53064 66402
rect 53354 66368 53370 66402
rect 53546 66368 53562 66402
rect 52788 66308 52822 66324
rect 53605 66358 53639 66374
rect 52856 66280 52872 66314
rect 53048 66280 53064 66314
rect 53354 66280 53370 66314
rect 53546 66280 53562 66314
rect 53605 66308 53639 66324
rect 52700 66210 52730 66262
rect 52640 66150 52730 66210
rect 52640 65910 52660 66150
rect 52700 66110 52730 66150
rect 52720 65952 52730 66110
rect 53700 66262 53708 66420
rect 53700 66230 53730 66262
rect 53770 66230 53790 66470
rect 53700 66150 53790 66230
rect 53700 66110 53730 66150
rect 52788 66048 52822 66064
rect 52856 66058 52872 66092
rect 53048 66058 53064 66092
rect 53354 66058 53370 66092
rect 53546 66058 53562 66092
rect 52788 65998 52822 66014
rect 53605 66048 53639 66064
rect 52856 65970 52872 66004
rect 53048 65970 53064 66004
rect 53354 65970 53370 66004
rect 53546 65970 53562 66004
rect 53605 65998 53639 66014
rect 52700 65910 52730 65952
rect 52640 65780 52730 65910
rect 53700 65952 53708 66110
rect 53700 65910 53730 65952
rect 53770 65910 53790 66150
rect 53700 65780 53790 65910
rect 57630 66470 57720 66590
rect 57630 66210 57650 66470
rect 57690 66420 57720 66470
rect 57710 66262 57720 66420
rect 58690 66470 58780 66590
rect 58690 66420 58720 66470
rect 57778 66358 57812 66374
rect 57846 66368 57862 66402
rect 58038 66368 58054 66402
rect 58344 66368 58360 66402
rect 58536 66368 58552 66402
rect 57778 66308 57812 66324
rect 58595 66358 58629 66374
rect 57846 66280 57862 66314
rect 58038 66280 58054 66314
rect 58344 66280 58360 66314
rect 58536 66280 58552 66314
rect 58595 66308 58629 66324
rect 57690 66210 57720 66262
rect 57630 66150 57720 66210
rect 57630 65910 57650 66150
rect 57690 66110 57720 66150
rect 57710 65952 57720 66110
rect 58690 66262 58698 66420
rect 58690 66230 58720 66262
rect 58760 66230 58780 66470
rect 58690 66150 58780 66230
rect 58690 66110 58720 66150
rect 57778 66048 57812 66064
rect 57846 66058 57862 66092
rect 58038 66058 58054 66092
rect 58344 66058 58360 66092
rect 58536 66058 58552 66092
rect 57778 65998 57812 66014
rect 58595 66048 58629 66064
rect 57846 65970 57862 66004
rect 58038 65970 58054 66004
rect 58344 65970 58360 66004
rect 58536 65970 58552 66004
rect 58595 65998 58629 66014
rect 57690 65910 57720 65952
rect 57630 65780 57720 65910
rect 58690 65952 58698 66110
rect 58690 65910 58720 65952
rect 58760 65910 58780 66150
rect 58690 65780 58780 65910
rect 62620 66470 62710 66590
rect 62620 66210 62640 66470
rect 62680 66420 62710 66470
rect 62700 66262 62710 66420
rect 63680 66470 63770 66590
rect 63680 66420 63710 66470
rect 62768 66358 62802 66374
rect 62836 66368 62852 66402
rect 63028 66368 63044 66402
rect 63334 66368 63350 66402
rect 63526 66368 63542 66402
rect 62768 66308 62802 66324
rect 63585 66358 63619 66374
rect 62836 66280 62852 66314
rect 63028 66280 63044 66314
rect 63334 66280 63350 66314
rect 63526 66280 63542 66314
rect 63585 66308 63619 66324
rect 62680 66210 62710 66262
rect 62620 66150 62710 66210
rect 62620 65910 62640 66150
rect 62680 66110 62710 66150
rect 62700 65952 62710 66110
rect 63680 66262 63688 66420
rect 63680 66230 63710 66262
rect 63750 66230 63770 66470
rect 63680 66150 63770 66230
rect 63680 66110 63710 66150
rect 62768 66048 62802 66064
rect 62836 66058 62852 66092
rect 63028 66058 63044 66092
rect 63334 66058 63350 66092
rect 63526 66058 63542 66092
rect 62768 65998 62802 66014
rect 63585 66048 63619 66064
rect 62836 65970 62852 66004
rect 63028 65970 63044 66004
rect 63334 65970 63350 66004
rect 63526 65970 63542 66004
rect 63585 65998 63619 66014
rect 62680 65910 62710 65952
rect 62620 65780 62710 65910
rect 63680 65952 63688 66110
rect 63680 65910 63710 65952
rect 63750 65910 63770 66150
rect 63680 65780 63770 65910
rect 67610 66470 67700 66590
rect 67610 66210 67630 66470
rect 67670 66420 67700 66470
rect 67690 66262 67700 66420
rect 68670 66470 68760 66590
rect 68670 66420 68700 66470
rect 67758 66358 67792 66374
rect 67826 66368 67842 66402
rect 68018 66368 68034 66402
rect 68324 66368 68340 66402
rect 68516 66368 68532 66402
rect 67758 66308 67792 66324
rect 68575 66358 68609 66374
rect 67826 66280 67842 66314
rect 68018 66280 68034 66314
rect 68324 66280 68340 66314
rect 68516 66280 68532 66314
rect 68575 66308 68609 66324
rect 67670 66210 67700 66262
rect 67610 66150 67700 66210
rect 67610 65910 67630 66150
rect 67670 66110 67700 66150
rect 67690 65952 67700 66110
rect 68670 66262 68678 66420
rect 68670 66230 68700 66262
rect 68740 66230 68760 66470
rect 68670 66150 68760 66230
rect 68670 66110 68700 66150
rect 67758 66048 67792 66064
rect 67826 66058 67842 66092
rect 68018 66058 68034 66092
rect 68324 66058 68340 66092
rect 68516 66058 68532 66092
rect 67758 65998 67792 66014
rect 68575 66048 68609 66064
rect 67826 65970 67842 66004
rect 68018 65970 68034 66004
rect 68324 65970 68340 66004
rect 68516 65970 68532 66004
rect 68575 65998 68609 66014
rect 67670 65910 67700 65952
rect 67610 65780 67700 65910
rect 68670 65952 68678 66110
rect 68670 65910 68700 65952
rect 68740 65910 68760 66150
rect 68670 65780 68760 65910
rect 72600 66470 72690 66590
rect 72600 66210 72620 66470
rect 72660 66420 72690 66470
rect 72680 66262 72690 66420
rect 73660 66470 73750 66590
rect 73660 66420 73690 66470
rect 72748 66358 72782 66374
rect 72816 66368 72832 66402
rect 73008 66368 73024 66402
rect 73314 66368 73330 66402
rect 73506 66368 73522 66402
rect 72748 66308 72782 66324
rect 73565 66358 73599 66374
rect 72816 66280 72832 66314
rect 73008 66280 73024 66314
rect 73314 66280 73330 66314
rect 73506 66280 73522 66314
rect 73565 66308 73599 66324
rect 72660 66210 72690 66262
rect 72600 66150 72690 66210
rect 72600 65910 72620 66150
rect 72660 66110 72690 66150
rect 72680 65952 72690 66110
rect 73660 66262 73668 66420
rect 73660 66230 73690 66262
rect 73730 66230 73750 66470
rect 73660 66150 73750 66230
rect 73660 66110 73690 66150
rect 72748 66048 72782 66064
rect 72816 66058 72832 66092
rect 73008 66058 73024 66092
rect 73314 66058 73330 66092
rect 73506 66058 73522 66092
rect 72748 65998 72782 66014
rect 73565 66048 73599 66064
rect 72816 65970 72832 66004
rect 73008 65970 73024 66004
rect 73314 65970 73330 66004
rect 73506 65970 73522 66004
rect 73565 65998 73599 66014
rect 72660 65910 72690 65952
rect 72600 65780 72690 65910
rect 73660 65952 73668 66110
rect 73660 65910 73690 65952
rect 73730 65910 73750 66150
rect 73660 65780 73750 65910
rect 77590 66470 77680 66590
rect 77590 66210 77610 66470
rect 77650 66420 77680 66470
rect 77670 66262 77680 66420
rect 78650 66470 78740 66590
rect 78650 66420 78680 66470
rect 77738 66358 77772 66374
rect 77806 66368 77822 66402
rect 77998 66368 78014 66402
rect 78304 66368 78320 66402
rect 78496 66368 78512 66402
rect 77738 66308 77772 66324
rect 78555 66358 78589 66374
rect 77806 66280 77822 66314
rect 77998 66280 78014 66314
rect 78304 66280 78320 66314
rect 78496 66280 78512 66314
rect 78555 66308 78589 66324
rect 77650 66210 77680 66262
rect 77590 66150 77680 66210
rect 77590 65910 77610 66150
rect 77650 66110 77680 66150
rect 77670 65952 77680 66110
rect 78650 66262 78658 66420
rect 78650 66230 78680 66262
rect 78720 66230 78740 66470
rect 78650 66150 78740 66230
rect 78650 66110 78680 66150
rect 77738 66048 77772 66064
rect 77806 66058 77822 66092
rect 77998 66058 78014 66092
rect 78304 66058 78320 66092
rect 78496 66058 78512 66092
rect 77738 65998 77772 66014
rect 78555 66048 78589 66064
rect 77806 65970 77822 66004
rect 77998 65970 78014 66004
rect 78304 65970 78320 66004
rect 78496 65970 78512 66004
rect 78555 65998 78589 66014
rect 77650 65910 77680 65952
rect 77590 65780 77680 65910
rect 78650 65952 78658 66110
rect 78650 65910 78680 65952
rect 78720 65910 78740 66150
rect 78650 65780 78740 65910
rect 2740 64760 2830 64880
rect 2740 64500 2760 64760
rect 2800 64710 2830 64760
rect 2820 64552 2830 64710
rect 3800 64760 3890 64880
rect 3800 64710 3830 64760
rect 2888 64648 2922 64664
rect 2956 64658 2972 64692
rect 3148 64658 3164 64692
rect 3454 64658 3470 64692
rect 3646 64658 3662 64692
rect 2888 64598 2922 64614
rect 3705 64648 3739 64664
rect 2956 64570 2972 64604
rect 3148 64570 3164 64604
rect 3454 64570 3470 64604
rect 3646 64570 3662 64604
rect 3705 64598 3739 64614
rect 2800 64500 2830 64552
rect 2740 64440 2830 64500
rect 2740 64200 2760 64440
rect 2800 64400 2830 64440
rect 2820 64242 2830 64400
rect 3800 64552 3808 64710
rect 3800 64520 3830 64552
rect 3870 64520 3890 64760
rect 3800 64440 3890 64520
rect 3800 64400 3830 64440
rect 2888 64338 2922 64354
rect 2956 64348 2972 64382
rect 3148 64348 3164 64382
rect 3454 64348 3470 64382
rect 3646 64348 3662 64382
rect 2888 64288 2922 64304
rect 3705 64338 3739 64354
rect 2956 64260 2972 64294
rect 3148 64260 3164 64294
rect 3454 64260 3470 64294
rect 3646 64260 3662 64294
rect 3705 64288 3739 64304
rect 2800 64200 2830 64242
rect 2740 64070 2830 64200
rect 3800 64242 3808 64400
rect 3800 64200 3830 64242
rect 3870 64200 3890 64440
rect 3800 64070 3890 64200
rect 7730 64760 7820 64880
rect 7730 64500 7750 64760
rect 7790 64710 7820 64760
rect 7810 64552 7820 64710
rect 8790 64760 8880 64880
rect 8790 64710 8820 64760
rect 7878 64648 7912 64664
rect 7946 64658 7962 64692
rect 8138 64658 8154 64692
rect 8444 64658 8460 64692
rect 8636 64658 8652 64692
rect 7878 64598 7912 64614
rect 8695 64648 8729 64664
rect 7946 64570 7962 64604
rect 8138 64570 8154 64604
rect 8444 64570 8460 64604
rect 8636 64570 8652 64604
rect 8695 64598 8729 64614
rect 7790 64500 7820 64552
rect 7730 64440 7820 64500
rect 7730 64200 7750 64440
rect 7790 64400 7820 64440
rect 7810 64242 7820 64400
rect 8790 64552 8798 64710
rect 8790 64520 8820 64552
rect 8860 64520 8880 64760
rect 8790 64440 8880 64520
rect 8790 64400 8820 64440
rect 7878 64338 7912 64354
rect 7946 64348 7962 64382
rect 8138 64348 8154 64382
rect 8444 64348 8460 64382
rect 8636 64348 8652 64382
rect 7878 64288 7912 64304
rect 8695 64338 8729 64354
rect 7946 64260 7962 64294
rect 8138 64260 8154 64294
rect 8444 64260 8460 64294
rect 8636 64260 8652 64294
rect 8695 64288 8729 64304
rect 7790 64200 7820 64242
rect 7730 64070 7820 64200
rect 8790 64242 8798 64400
rect 8790 64200 8820 64242
rect 8860 64200 8880 64440
rect 8790 64070 8880 64200
rect 12720 64760 12810 64880
rect 12720 64500 12740 64760
rect 12780 64710 12810 64760
rect 12800 64552 12810 64710
rect 13780 64760 13870 64880
rect 13780 64710 13810 64760
rect 12868 64648 12902 64664
rect 12936 64658 12952 64692
rect 13128 64658 13144 64692
rect 13434 64658 13450 64692
rect 13626 64658 13642 64692
rect 12868 64598 12902 64614
rect 13685 64648 13719 64664
rect 12936 64570 12952 64604
rect 13128 64570 13144 64604
rect 13434 64570 13450 64604
rect 13626 64570 13642 64604
rect 13685 64598 13719 64614
rect 12780 64500 12810 64552
rect 12720 64440 12810 64500
rect 12720 64200 12740 64440
rect 12780 64400 12810 64440
rect 12800 64242 12810 64400
rect 13780 64552 13788 64710
rect 13780 64520 13810 64552
rect 13850 64520 13870 64760
rect 13780 64440 13870 64520
rect 13780 64400 13810 64440
rect 12868 64338 12902 64354
rect 12936 64348 12952 64382
rect 13128 64348 13144 64382
rect 13434 64348 13450 64382
rect 13626 64348 13642 64382
rect 12868 64288 12902 64304
rect 13685 64338 13719 64354
rect 12936 64260 12952 64294
rect 13128 64260 13144 64294
rect 13434 64260 13450 64294
rect 13626 64260 13642 64294
rect 13685 64288 13719 64304
rect 12780 64200 12810 64242
rect 12720 64070 12810 64200
rect 13780 64242 13788 64400
rect 13780 64200 13810 64242
rect 13850 64200 13870 64440
rect 13780 64070 13870 64200
rect 17710 64760 17800 64880
rect 17710 64500 17730 64760
rect 17770 64710 17800 64760
rect 17790 64552 17800 64710
rect 18770 64760 18860 64880
rect 18770 64710 18800 64760
rect 17858 64648 17892 64664
rect 17926 64658 17942 64692
rect 18118 64658 18134 64692
rect 18424 64658 18440 64692
rect 18616 64658 18632 64692
rect 17858 64598 17892 64614
rect 18675 64648 18709 64664
rect 17926 64570 17942 64604
rect 18118 64570 18134 64604
rect 18424 64570 18440 64604
rect 18616 64570 18632 64604
rect 18675 64598 18709 64614
rect 17770 64500 17800 64552
rect 17710 64440 17800 64500
rect 17710 64200 17730 64440
rect 17770 64400 17800 64440
rect 17790 64242 17800 64400
rect 18770 64552 18778 64710
rect 18770 64520 18800 64552
rect 18840 64520 18860 64760
rect 18770 64440 18860 64520
rect 18770 64400 18800 64440
rect 17858 64338 17892 64354
rect 17926 64348 17942 64382
rect 18118 64348 18134 64382
rect 18424 64348 18440 64382
rect 18616 64348 18632 64382
rect 17858 64288 17892 64304
rect 18675 64338 18709 64354
rect 17926 64260 17942 64294
rect 18118 64260 18134 64294
rect 18424 64260 18440 64294
rect 18616 64260 18632 64294
rect 18675 64288 18709 64304
rect 17770 64200 17800 64242
rect 17710 64070 17800 64200
rect 18770 64242 18778 64400
rect 18770 64200 18800 64242
rect 18840 64200 18860 64440
rect 18770 64070 18860 64200
rect 22700 64760 22790 64880
rect 22700 64500 22720 64760
rect 22760 64710 22790 64760
rect 22780 64552 22790 64710
rect 23760 64760 23850 64880
rect 23760 64710 23790 64760
rect 22848 64648 22882 64664
rect 22916 64658 22932 64692
rect 23108 64658 23124 64692
rect 23414 64658 23430 64692
rect 23606 64658 23622 64692
rect 22848 64598 22882 64614
rect 23665 64648 23699 64664
rect 22916 64570 22932 64604
rect 23108 64570 23124 64604
rect 23414 64570 23430 64604
rect 23606 64570 23622 64604
rect 23665 64598 23699 64614
rect 22760 64500 22790 64552
rect 22700 64440 22790 64500
rect 22700 64200 22720 64440
rect 22760 64400 22790 64440
rect 22780 64242 22790 64400
rect 23760 64552 23768 64710
rect 23760 64520 23790 64552
rect 23830 64520 23850 64760
rect 23760 64440 23850 64520
rect 23760 64400 23790 64440
rect 22848 64338 22882 64354
rect 22916 64348 22932 64382
rect 23108 64348 23124 64382
rect 23414 64348 23430 64382
rect 23606 64348 23622 64382
rect 22848 64288 22882 64304
rect 23665 64338 23699 64354
rect 22916 64260 22932 64294
rect 23108 64260 23124 64294
rect 23414 64260 23430 64294
rect 23606 64260 23622 64294
rect 23665 64288 23699 64304
rect 22760 64200 22790 64242
rect 22700 64070 22790 64200
rect 23760 64242 23768 64400
rect 23760 64200 23790 64242
rect 23830 64200 23850 64440
rect 23760 64070 23850 64200
rect 27690 64760 27780 64880
rect 27690 64500 27710 64760
rect 27750 64710 27780 64760
rect 27770 64552 27780 64710
rect 28750 64760 28840 64880
rect 28750 64710 28780 64760
rect 27838 64648 27872 64664
rect 27906 64658 27922 64692
rect 28098 64658 28114 64692
rect 28404 64658 28420 64692
rect 28596 64658 28612 64692
rect 27838 64598 27872 64614
rect 28655 64648 28689 64664
rect 27906 64570 27922 64604
rect 28098 64570 28114 64604
rect 28404 64570 28420 64604
rect 28596 64570 28612 64604
rect 28655 64598 28689 64614
rect 27750 64500 27780 64552
rect 27690 64440 27780 64500
rect 27690 64200 27710 64440
rect 27750 64400 27780 64440
rect 27770 64242 27780 64400
rect 28750 64552 28758 64710
rect 28750 64520 28780 64552
rect 28820 64520 28840 64760
rect 28750 64440 28840 64520
rect 28750 64400 28780 64440
rect 27838 64338 27872 64354
rect 27906 64348 27922 64382
rect 28098 64348 28114 64382
rect 28404 64348 28420 64382
rect 28596 64348 28612 64382
rect 27838 64288 27872 64304
rect 28655 64338 28689 64354
rect 27906 64260 27922 64294
rect 28098 64260 28114 64294
rect 28404 64260 28420 64294
rect 28596 64260 28612 64294
rect 28655 64288 28689 64304
rect 27750 64200 27780 64242
rect 27690 64070 27780 64200
rect 28750 64242 28758 64400
rect 28750 64200 28780 64242
rect 28820 64200 28840 64440
rect 28750 64070 28840 64200
rect 32680 64760 32770 64880
rect 32680 64500 32700 64760
rect 32740 64710 32770 64760
rect 32760 64552 32770 64710
rect 33740 64760 33830 64880
rect 33740 64710 33770 64760
rect 32828 64648 32862 64664
rect 32896 64658 32912 64692
rect 33088 64658 33104 64692
rect 33394 64658 33410 64692
rect 33586 64658 33602 64692
rect 32828 64598 32862 64614
rect 33645 64648 33679 64664
rect 32896 64570 32912 64604
rect 33088 64570 33104 64604
rect 33394 64570 33410 64604
rect 33586 64570 33602 64604
rect 33645 64598 33679 64614
rect 32740 64500 32770 64552
rect 32680 64440 32770 64500
rect 32680 64200 32700 64440
rect 32740 64400 32770 64440
rect 32760 64242 32770 64400
rect 33740 64552 33748 64710
rect 33740 64520 33770 64552
rect 33810 64520 33830 64760
rect 33740 64440 33830 64520
rect 33740 64400 33770 64440
rect 32828 64338 32862 64354
rect 32896 64348 32912 64382
rect 33088 64348 33104 64382
rect 33394 64348 33410 64382
rect 33586 64348 33602 64382
rect 32828 64288 32862 64304
rect 33645 64338 33679 64354
rect 32896 64260 32912 64294
rect 33088 64260 33104 64294
rect 33394 64260 33410 64294
rect 33586 64260 33602 64294
rect 33645 64288 33679 64304
rect 32740 64200 32770 64242
rect 32680 64070 32770 64200
rect 33740 64242 33748 64400
rect 33740 64200 33770 64242
rect 33810 64200 33830 64440
rect 33740 64070 33830 64200
rect 37670 64760 37760 64880
rect 37670 64500 37690 64760
rect 37730 64710 37760 64760
rect 37750 64552 37760 64710
rect 38730 64760 38820 64880
rect 38730 64710 38760 64760
rect 37818 64648 37852 64664
rect 37886 64658 37902 64692
rect 38078 64658 38094 64692
rect 38384 64658 38400 64692
rect 38576 64658 38592 64692
rect 37818 64598 37852 64614
rect 38635 64648 38669 64664
rect 37886 64570 37902 64604
rect 38078 64570 38094 64604
rect 38384 64570 38400 64604
rect 38576 64570 38592 64604
rect 38635 64598 38669 64614
rect 37730 64500 37760 64552
rect 37670 64440 37760 64500
rect 37670 64200 37690 64440
rect 37730 64400 37760 64440
rect 37750 64242 37760 64400
rect 38730 64552 38738 64710
rect 38730 64520 38760 64552
rect 38800 64520 38820 64760
rect 38730 64440 38820 64520
rect 38730 64400 38760 64440
rect 37818 64338 37852 64354
rect 37886 64348 37902 64382
rect 38078 64348 38094 64382
rect 38384 64348 38400 64382
rect 38576 64348 38592 64382
rect 37818 64288 37852 64304
rect 38635 64338 38669 64354
rect 37886 64260 37902 64294
rect 38078 64260 38094 64294
rect 38384 64260 38400 64294
rect 38576 64260 38592 64294
rect 38635 64288 38669 64304
rect 37730 64200 37760 64242
rect 37670 64070 37760 64200
rect 38730 64242 38738 64400
rect 38730 64200 38760 64242
rect 38800 64200 38820 64440
rect 38730 64070 38820 64200
rect 42660 64760 42750 64880
rect 42660 64500 42680 64760
rect 42720 64710 42750 64760
rect 42740 64552 42750 64710
rect 43720 64760 43810 64880
rect 43720 64710 43750 64760
rect 42808 64648 42842 64664
rect 42876 64658 42892 64692
rect 43068 64658 43084 64692
rect 43374 64658 43390 64692
rect 43566 64658 43582 64692
rect 42808 64598 42842 64614
rect 43625 64648 43659 64664
rect 42876 64570 42892 64604
rect 43068 64570 43084 64604
rect 43374 64570 43390 64604
rect 43566 64570 43582 64604
rect 43625 64598 43659 64614
rect 42720 64500 42750 64552
rect 42660 64440 42750 64500
rect 42660 64200 42680 64440
rect 42720 64400 42750 64440
rect 42740 64242 42750 64400
rect 43720 64552 43728 64710
rect 43720 64520 43750 64552
rect 43790 64520 43810 64760
rect 43720 64440 43810 64520
rect 43720 64400 43750 64440
rect 42808 64338 42842 64354
rect 42876 64348 42892 64382
rect 43068 64348 43084 64382
rect 43374 64348 43390 64382
rect 43566 64348 43582 64382
rect 42808 64288 42842 64304
rect 43625 64338 43659 64354
rect 42876 64260 42892 64294
rect 43068 64260 43084 64294
rect 43374 64260 43390 64294
rect 43566 64260 43582 64294
rect 43625 64288 43659 64304
rect 42720 64200 42750 64242
rect 42660 64070 42750 64200
rect 43720 64242 43728 64400
rect 43720 64200 43750 64242
rect 43790 64200 43810 64440
rect 43720 64070 43810 64200
rect 47650 64760 47740 64880
rect 47650 64500 47670 64760
rect 47710 64710 47740 64760
rect 47730 64552 47740 64710
rect 48710 64760 48800 64880
rect 48710 64710 48740 64760
rect 47798 64648 47832 64664
rect 47866 64658 47882 64692
rect 48058 64658 48074 64692
rect 48364 64658 48380 64692
rect 48556 64658 48572 64692
rect 47798 64598 47832 64614
rect 48615 64648 48649 64664
rect 47866 64570 47882 64604
rect 48058 64570 48074 64604
rect 48364 64570 48380 64604
rect 48556 64570 48572 64604
rect 48615 64598 48649 64614
rect 47710 64500 47740 64552
rect 47650 64440 47740 64500
rect 47650 64200 47670 64440
rect 47710 64400 47740 64440
rect 47730 64242 47740 64400
rect 48710 64552 48718 64710
rect 48710 64520 48740 64552
rect 48780 64520 48800 64760
rect 48710 64440 48800 64520
rect 48710 64400 48740 64440
rect 47798 64338 47832 64354
rect 47866 64348 47882 64382
rect 48058 64348 48074 64382
rect 48364 64348 48380 64382
rect 48556 64348 48572 64382
rect 47798 64288 47832 64304
rect 48615 64338 48649 64354
rect 47866 64260 47882 64294
rect 48058 64260 48074 64294
rect 48364 64260 48380 64294
rect 48556 64260 48572 64294
rect 48615 64288 48649 64304
rect 47710 64200 47740 64242
rect 47650 64070 47740 64200
rect 48710 64242 48718 64400
rect 48710 64200 48740 64242
rect 48780 64200 48800 64440
rect 48710 64070 48800 64200
rect 52640 64760 52730 64880
rect 52640 64500 52660 64760
rect 52700 64710 52730 64760
rect 52720 64552 52730 64710
rect 53700 64760 53790 64880
rect 53700 64710 53730 64760
rect 52788 64648 52822 64664
rect 52856 64658 52872 64692
rect 53048 64658 53064 64692
rect 53354 64658 53370 64692
rect 53546 64658 53562 64692
rect 52788 64598 52822 64614
rect 53605 64648 53639 64664
rect 52856 64570 52872 64604
rect 53048 64570 53064 64604
rect 53354 64570 53370 64604
rect 53546 64570 53562 64604
rect 53605 64598 53639 64614
rect 52700 64500 52730 64552
rect 52640 64440 52730 64500
rect 52640 64200 52660 64440
rect 52700 64400 52730 64440
rect 52720 64242 52730 64400
rect 53700 64552 53708 64710
rect 53700 64520 53730 64552
rect 53770 64520 53790 64760
rect 53700 64440 53790 64520
rect 53700 64400 53730 64440
rect 52788 64338 52822 64354
rect 52856 64348 52872 64382
rect 53048 64348 53064 64382
rect 53354 64348 53370 64382
rect 53546 64348 53562 64382
rect 52788 64288 52822 64304
rect 53605 64338 53639 64354
rect 52856 64260 52872 64294
rect 53048 64260 53064 64294
rect 53354 64260 53370 64294
rect 53546 64260 53562 64294
rect 53605 64288 53639 64304
rect 52700 64200 52730 64242
rect 52640 64070 52730 64200
rect 53700 64242 53708 64400
rect 53700 64200 53730 64242
rect 53770 64200 53790 64440
rect 53700 64070 53790 64200
rect 57630 64760 57720 64880
rect 57630 64500 57650 64760
rect 57690 64710 57720 64760
rect 57710 64552 57720 64710
rect 58690 64760 58780 64880
rect 58690 64710 58720 64760
rect 57778 64648 57812 64664
rect 57846 64658 57862 64692
rect 58038 64658 58054 64692
rect 58344 64658 58360 64692
rect 58536 64658 58552 64692
rect 57778 64598 57812 64614
rect 58595 64648 58629 64664
rect 57846 64570 57862 64604
rect 58038 64570 58054 64604
rect 58344 64570 58360 64604
rect 58536 64570 58552 64604
rect 58595 64598 58629 64614
rect 57690 64500 57720 64552
rect 57630 64440 57720 64500
rect 57630 64200 57650 64440
rect 57690 64400 57720 64440
rect 57710 64242 57720 64400
rect 58690 64552 58698 64710
rect 58690 64520 58720 64552
rect 58760 64520 58780 64760
rect 58690 64440 58780 64520
rect 58690 64400 58720 64440
rect 57778 64338 57812 64354
rect 57846 64348 57862 64382
rect 58038 64348 58054 64382
rect 58344 64348 58360 64382
rect 58536 64348 58552 64382
rect 57778 64288 57812 64304
rect 58595 64338 58629 64354
rect 57846 64260 57862 64294
rect 58038 64260 58054 64294
rect 58344 64260 58360 64294
rect 58536 64260 58552 64294
rect 58595 64288 58629 64304
rect 57690 64200 57720 64242
rect 57630 64070 57720 64200
rect 58690 64242 58698 64400
rect 58690 64200 58720 64242
rect 58760 64200 58780 64440
rect 58690 64070 58780 64200
rect 62620 64760 62710 64880
rect 62620 64500 62640 64760
rect 62680 64710 62710 64760
rect 62700 64552 62710 64710
rect 63680 64760 63770 64880
rect 63680 64710 63710 64760
rect 62768 64648 62802 64664
rect 62836 64658 62852 64692
rect 63028 64658 63044 64692
rect 63334 64658 63350 64692
rect 63526 64658 63542 64692
rect 62768 64598 62802 64614
rect 63585 64648 63619 64664
rect 62836 64570 62852 64604
rect 63028 64570 63044 64604
rect 63334 64570 63350 64604
rect 63526 64570 63542 64604
rect 63585 64598 63619 64614
rect 62680 64500 62710 64552
rect 62620 64440 62710 64500
rect 62620 64200 62640 64440
rect 62680 64400 62710 64440
rect 62700 64242 62710 64400
rect 63680 64552 63688 64710
rect 63680 64520 63710 64552
rect 63750 64520 63770 64760
rect 63680 64440 63770 64520
rect 63680 64400 63710 64440
rect 62768 64338 62802 64354
rect 62836 64348 62852 64382
rect 63028 64348 63044 64382
rect 63334 64348 63350 64382
rect 63526 64348 63542 64382
rect 62768 64288 62802 64304
rect 63585 64338 63619 64354
rect 62836 64260 62852 64294
rect 63028 64260 63044 64294
rect 63334 64260 63350 64294
rect 63526 64260 63542 64294
rect 63585 64288 63619 64304
rect 62680 64200 62710 64242
rect 62620 64070 62710 64200
rect 63680 64242 63688 64400
rect 63680 64200 63710 64242
rect 63750 64200 63770 64440
rect 63680 64070 63770 64200
rect 67610 64760 67700 64880
rect 67610 64500 67630 64760
rect 67670 64710 67700 64760
rect 67690 64552 67700 64710
rect 68670 64760 68760 64880
rect 68670 64710 68700 64760
rect 67758 64648 67792 64664
rect 67826 64658 67842 64692
rect 68018 64658 68034 64692
rect 68324 64658 68340 64692
rect 68516 64658 68532 64692
rect 67758 64598 67792 64614
rect 68575 64648 68609 64664
rect 67826 64570 67842 64604
rect 68018 64570 68034 64604
rect 68324 64570 68340 64604
rect 68516 64570 68532 64604
rect 68575 64598 68609 64614
rect 67670 64500 67700 64552
rect 67610 64440 67700 64500
rect 67610 64200 67630 64440
rect 67670 64400 67700 64440
rect 67690 64242 67700 64400
rect 68670 64552 68678 64710
rect 68670 64520 68700 64552
rect 68740 64520 68760 64760
rect 68670 64440 68760 64520
rect 68670 64400 68700 64440
rect 67758 64338 67792 64354
rect 67826 64348 67842 64382
rect 68018 64348 68034 64382
rect 68324 64348 68340 64382
rect 68516 64348 68532 64382
rect 67758 64288 67792 64304
rect 68575 64338 68609 64354
rect 67826 64260 67842 64294
rect 68018 64260 68034 64294
rect 68324 64260 68340 64294
rect 68516 64260 68532 64294
rect 68575 64288 68609 64304
rect 67670 64200 67700 64242
rect 67610 64070 67700 64200
rect 68670 64242 68678 64400
rect 68670 64200 68700 64242
rect 68740 64200 68760 64440
rect 68670 64070 68760 64200
rect 72600 64760 72690 64880
rect 72600 64500 72620 64760
rect 72660 64710 72690 64760
rect 72680 64552 72690 64710
rect 73660 64760 73750 64880
rect 73660 64710 73690 64760
rect 72748 64648 72782 64664
rect 72816 64658 72832 64692
rect 73008 64658 73024 64692
rect 73314 64658 73330 64692
rect 73506 64658 73522 64692
rect 72748 64598 72782 64614
rect 73565 64648 73599 64664
rect 72816 64570 72832 64604
rect 73008 64570 73024 64604
rect 73314 64570 73330 64604
rect 73506 64570 73522 64604
rect 73565 64598 73599 64614
rect 72660 64500 72690 64552
rect 72600 64440 72690 64500
rect 72600 64200 72620 64440
rect 72660 64400 72690 64440
rect 72680 64242 72690 64400
rect 73660 64552 73668 64710
rect 73660 64520 73690 64552
rect 73730 64520 73750 64760
rect 73660 64440 73750 64520
rect 73660 64400 73690 64440
rect 72748 64338 72782 64354
rect 72816 64348 72832 64382
rect 73008 64348 73024 64382
rect 73314 64348 73330 64382
rect 73506 64348 73522 64382
rect 72748 64288 72782 64304
rect 73565 64338 73599 64354
rect 72816 64260 72832 64294
rect 73008 64260 73024 64294
rect 73314 64260 73330 64294
rect 73506 64260 73522 64294
rect 73565 64288 73599 64304
rect 72660 64200 72690 64242
rect 72600 64070 72690 64200
rect 73660 64242 73668 64400
rect 73660 64200 73690 64242
rect 73730 64200 73750 64440
rect 73660 64070 73750 64200
rect 77590 64760 77680 64880
rect 77590 64500 77610 64760
rect 77650 64710 77680 64760
rect 77670 64552 77680 64710
rect 78650 64760 78740 64880
rect 78650 64710 78680 64760
rect 77738 64648 77772 64664
rect 77806 64658 77822 64692
rect 77998 64658 78014 64692
rect 78304 64658 78320 64692
rect 78496 64658 78512 64692
rect 77738 64598 77772 64614
rect 78555 64648 78589 64664
rect 77806 64570 77822 64604
rect 77998 64570 78014 64604
rect 78304 64570 78320 64604
rect 78496 64570 78512 64604
rect 78555 64598 78589 64614
rect 77650 64500 77680 64552
rect 77590 64440 77680 64500
rect 77590 64200 77610 64440
rect 77650 64400 77680 64440
rect 77670 64242 77680 64400
rect 78650 64552 78658 64710
rect 78650 64520 78680 64552
rect 78720 64520 78740 64760
rect 78650 64440 78740 64520
rect 78650 64400 78680 64440
rect 77738 64338 77772 64354
rect 77806 64348 77822 64382
rect 77998 64348 78014 64382
rect 78304 64348 78320 64382
rect 78496 64348 78512 64382
rect 77738 64288 77772 64304
rect 78555 64338 78589 64354
rect 77806 64260 77822 64294
rect 77998 64260 78014 64294
rect 78304 64260 78320 64294
rect 78496 64260 78512 64294
rect 78555 64288 78589 64304
rect 77650 64200 77680 64242
rect 77590 64070 77680 64200
rect 78650 64242 78658 64400
rect 78650 64200 78680 64242
rect 78720 64200 78740 64440
rect 78650 64070 78740 64200
rect 2740 63050 2830 63170
rect 2740 62790 2760 63050
rect 2800 63000 2830 63050
rect 2820 62842 2830 63000
rect 3800 63050 3890 63170
rect 3800 63000 3830 63050
rect 2888 62938 2922 62954
rect 2956 62948 2972 62982
rect 3148 62948 3164 62982
rect 3454 62948 3470 62982
rect 3646 62948 3662 62982
rect 2888 62888 2922 62904
rect 3705 62938 3739 62954
rect 2956 62860 2972 62894
rect 3148 62860 3164 62894
rect 3454 62860 3470 62894
rect 3646 62860 3662 62894
rect 3705 62888 3739 62904
rect 2800 62790 2830 62842
rect 2740 62730 2830 62790
rect 2740 62490 2760 62730
rect 2800 62690 2830 62730
rect 2820 62532 2830 62690
rect 3800 62842 3808 63000
rect 3800 62810 3830 62842
rect 3870 62810 3890 63050
rect 3800 62730 3890 62810
rect 3800 62690 3830 62730
rect 2888 62628 2922 62644
rect 2956 62638 2972 62672
rect 3148 62638 3164 62672
rect 3454 62638 3470 62672
rect 3646 62638 3662 62672
rect 2888 62578 2922 62594
rect 3705 62628 3739 62644
rect 2956 62550 2972 62584
rect 3148 62550 3164 62584
rect 3454 62550 3470 62584
rect 3646 62550 3662 62584
rect 3705 62578 3739 62594
rect 2800 62490 2830 62532
rect 2740 62360 2830 62490
rect 3800 62532 3808 62690
rect 3800 62490 3830 62532
rect 3870 62490 3890 62730
rect 3800 62360 3890 62490
rect 7730 63050 7820 63170
rect 7730 62790 7750 63050
rect 7790 63000 7820 63050
rect 7810 62842 7820 63000
rect 8790 63050 8880 63170
rect 8790 63000 8820 63050
rect 7878 62938 7912 62954
rect 7946 62948 7962 62982
rect 8138 62948 8154 62982
rect 8444 62948 8460 62982
rect 8636 62948 8652 62982
rect 7878 62888 7912 62904
rect 8695 62938 8729 62954
rect 7946 62860 7962 62894
rect 8138 62860 8154 62894
rect 8444 62860 8460 62894
rect 8636 62860 8652 62894
rect 8695 62888 8729 62904
rect 7790 62790 7820 62842
rect 7730 62730 7820 62790
rect 7730 62490 7750 62730
rect 7790 62690 7820 62730
rect 7810 62532 7820 62690
rect 8790 62842 8798 63000
rect 8790 62810 8820 62842
rect 8860 62810 8880 63050
rect 8790 62730 8880 62810
rect 8790 62690 8820 62730
rect 7878 62628 7912 62644
rect 7946 62638 7962 62672
rect 8138 62638 8154 62672
rect 8444 62638 8460 62672
rect 8636 62638 8652 62672
rect 7878 62578 7912 62594
rect 8695 62628 8729 62644
rect 7946 62550 7962 62584
rect 8138 62550 8154 62584
rect 8444 62550 8460 62584
rect 8636 62550 8652 62584
rect 8695 62578 8729 62594
rect 7790 62490 7820 62532
rect 7730 62360 7820 62490
rect 8790 62532 8798 62690
rect 8790 62490 8820 62532
rect 8860 62490 8880 62730
rect 8790 62360 8880 62490
rect 12720 63050 12810 63170
rect 12720 62790 12740 63050
rect 12780 63000 12810 63050
rect 12800 62842 12810 63000
rect 13780 63050 13870 63170
rect 13780 63000 13810 63050
rect 12868 62938 12902 62954
rect 12936 62948 12952 62982
rect 13128 62948 13144 62982
rect 13434 62948 13450 62982
rect 13626 62948 13642 62982
rect 12868 62888 12902 62904
rect 13685 62938 13719 62954
rect 12936 62860 12952 62894
rect 13128 62860 13144 62894
rect 13434 62860 13450 62894
rect 13626 62860 13642 62894
rect 13685 62888 13719 62904
rect 12780 62790 12810 62842
rect 12720 62730 12810 62790
rect 12720 62490 12740 62730
rect 12780 62690 12810 62730
rect 12800 62532 12810 62690
rect 13780 62842 13788 63000
rect 13780 62810 13810 62842
rect 13850 62810 13870 63050
rect 13780 62730 13870 62810
rect 13780 62690 13810 62730
rect 12868 62628 12902 62644
rect 12936 62638 12952 62672
rect 13128 62638 13144 62672
rect 13434 62638 13450 62672
rect 13626 62638 13642 62672
rect 12868 62578 12902 62594
rect 13685 62628 13719 62644
rect 12936 62550 12952 62584
rect 13128 62550 13144 62584
rect 13434 62550 13450 62584
rect 13626 62550 13642 62584
rect 13685 62578 13719 62594
rect 12780 62490 12810 62532
rect 12720 62360 12810 62490
rect 13780 62532 13788 62690
rect 13780 62490 13810 62532
rect 13850 62490 13870 62730
rect 13780 62360 13870 62490
rect 17710 63050 17800 63170
rect 17710 62790 17730 63050
rect 17770 63000 17800 63050
rect 17790 62842 17800 63000
rect 18770 63050 18860 63170
rect 18770 63000 18800 63050
rect 17858 62938 17892 62954
rect 17926 62948 17942 62982
rect 18118 62948 18134 62982
rect 18424 62948 18440 62982
rect 18616 62948 18632 62982
rect 17858 62888 17892 62904
rect 18675 62938 18709 62954
rect 17926 62860 17942 62894
rect 18118 62860 18134 62894
rect 18424 62860 18440 62894
rect 18616 62860 18632 62894
rect 18675 62888 18709 62904
rect 17770 62790 17800 62842
rect 17710 62730 17800 62790
rect 17710 62490 17730 62730
rect 17770 62690 17800 62730
rect 17790 62532 17800 62690
rect 18770 62842 18778 63000
rect 18770 62810 18800 62842
rect 18840 62810 18860 63050
rect 18770 62730 18860 62810
rect 18770 62690 18800 62730
rect 17858 62628 17892 62644
rect 17926 62638 17942 62672
rect 18118 62638 18134 62672
rect 18424 62638 18440 62672
rect 18616 62638 18632 62672
rect 17858 62578 17892 62594
rect 18675 62628 18709 62644
rect 17926 62550 17942 62584
rect 18118 62550 18134 62584
rect 18424 62550 18440 62584
rect 18616 62550 18632 62584
rect 18675 62578 18709 62594
rect 17770 62490 17800 62532
rect 17710 62360 17800 62490
rect 18770 62532 18778 62690
rect 18770 62490 18800 62532
rect 18840 62490 18860 62730
rect 18770 62360 18860 62490
rect 22700 63050 22790 63170
rect 22700 62790 22720 63050
rect 22760 63000 22790 63050
rect 22780 62842 22790 63000
rect 23760 63050 23850 63170
rect 23760 63000 23790 63050
rect 22848 62938 22882 62954
rect 22916 62948 22932 62982
rect 23108 62948 23124 62982
rect 23414 62948 23430 62982
rect 23606 62948 23622 62982
rect 22848 62888 22882 62904
rect 23665 62938 23699 62954
rect 22916 62860 22932 62894
rect 23108 62860 23124 62894
rect 23414 62860 23430 62894
rect 23606 62860 23622 62894
rect 23665 62888 23699 62904
rect 22760 62790 22790 62842
rect 22700 62730 22790 62790
rect 22700 62490 22720 62730
rect 22760 62690 22790 62730
rect 22780 62532 22790 62690
rect 23760 62842 23768 63000
rect 23760 62810 23790 62842
rect 23830 62810 23850 63050
rect 23760 62730 23850 62810
rect 23760 62690 23790 62730
rect 22848 62628 22882 62644
rect 22916 62638 22932 62672
rect 23108 62638 23124 62672
rect 23414 62638 23430 62672
rect 23606 62638 23622 62672
rect 22848 62578 22882 62594
rect 23665 62628 23699 62644
rect 22916 62550 22932 62584
rect 23108 62550 23124 62584
rect 23414 62550 23430 62584
rect 23606 62550 23622 62584
rect 23665 62578 23699 62594
rect 22760 62490 22790 62532
rect 22700 62360 22790 62490
rect 23760 62532 23768 62690
rect 23760 62490 23790 62532
rect 23830 62490 23850 62730
rect 23760 62360 23850 62490
rect 27690 63050 27780 63170
rect 27690 62790 27710 63050
rect 27750 63000 27780 63050
rect 27770 62842 27780 63000
rect 28750 63050 28840 63170
rect 28750 63000 28780 63050
rect 27838 62938 27872 62954
rect 27906 62948 27922 62982
rect 28098 62948 28114 62982
rect 28404 62948 28420 62982
rect 28596 62948 28612 62982
rect 27838 62888 27872 62904
rect 28655 62938 28689 62954
rect 27906 62860 27922 62894
rect 28098 62860 28114 62894
rect 28404 62860 28420 62894
rect 28596 62860 28612 62894
rect 28655 62888 28689 62904
rect 27750 62790 27780 62842
rect 27690 62730 27780 62790
rect 27690 62490 27710 62730
rect 27750 62690 27780 62730
rect 27770 62532 27780 62690
rect 28750 62842 28758 63000
rect 28750 62810 28780 62842
rect 28820 62810 28840 63050
rect 28750 62730 28840 62810
rect 28750 62690 28780 62730
rect 27838 62628 27872 62644
rect 27906 62638 27922 62672
rect 28098 62638 28114 62672
rect 28404 62638 28420 62672
rect 28596 62638 28612 62672
rect 27838 62578 27872 62594
rect 28655 62628 28689 62644
rect 27906 62550 27922 62584
rect 28098 62550 28114 62584
rect 28404 62550 28420 62584
rect 28596 62550 28612 62584
rect 28655 62578 28689 62594
rect 27750 62490 27780 62532
rect 27690 62360 27780 62490
rect 28750 62532 28758 62690
rect 28750 62490 28780 62532
rect 28820 62490 28840 62730
rect 28750 62360 28840 62490
rect 32680 63050 32770 63170
rect 32680 62790 32700 63050
rect 32740 63000 32770 63050
rect 32760 62842 32770 63000
rect 33740 63050 33830 63170
rect 33740 63000 33770 63050
rect 32828 62938 32862 62954
rect 32896 62948 32912 62982
rect 33088 62948 33104 62982
rect 33394 62948 33410 62982
rect 33586 62948 33602 62982
rect 32828 62888 32862 62904
rect 33645 62938 33679 62954
rect 32896 62860 32912 62894
rect 33088 62860 33104 62894
rect 33394 62860 33410 62894
rect 33586 62860 33602 62894
rect 33645 62888 33679 62904
rect 32740 62790 32770 62842
rect 32680 62730 32770 62790
rect 32680 62490 32700 62730
rect 32740 62690 32770 62730
rect 32760 62532 32770 62690
rect 33740 62842 33748 63000
rect 33740 62810 33770 62842
rect 33810 62810 33830 63050
rect 33740 62730 33830 62810
rect 33740 62690 33770 62730
rect 32828 62628 32862 62644
rect 32896 62638 32912 62672
rect 33088 62638 33104 62672
rect 33394 62638 33410 62672
rect 33586 62638 33602 62672
rect 32828 62578 32862 62594
rect 33645 62628 33679 62644
rect 32896 62550 32912 62584
rect 33088 62550 33104 62584
rect 33394 62550 33410 62584
rect 33586 62550 33602 62584
rect 33645 62578 33679 62594
rect 32740 62490 32770 62532
rect 32680 62360 32770 62490
rect 33740 62532 33748 62690
rect 33740 62490 33770 62532
rect 33810 62490 33830 62730
rect 33740 62360 33830 62490
rect 37670 63050 37760 63170
rect 37670 62790 37690 63050
rect 37730 63000 37760 63050
rect 37750 62842 37760 63000
rect 38730 63050 38820 63170
rect 38730 63000 38760 63050
rect 37818 62938 37852 62954
rect 37886 62948 37902 62982
rect 38078 62948 38094 62982
rect 38384 62948 38400 62982
rect 38576 62948 38592 62982
rect 37818 62888 37852 62904
rect 38635 62938 38669 62954
rect 37886 62860 37902 62894
rect 38078 62860 38094 62894
rect 38384 62860 38400 62894
rect 38576 62860 38592 62894
rect 38635 62888 38669 62904
rect 37730 62790 37760 62842
rect 37670 62730 37760 62790
rect 37670 62490 37690 62730
rect 37730 62690 37760 62730
rect 37750 62532 37760 62690
rect 38730 62842 38738 63000
rect 38730 62810 38760 62842
rect 38800 62810 38820 63050
rect 38730 62730 38820 62810
rect 38730 62690 38760 62730
rect 37818 62628 37852 62644
rect 37886 62638 37902 62672
rect 38078 62638 38094 62672
rect 38384 62638 38400 62672
rect 38576 62638 38592 62672
rect 37818 62578 37852 62594
rect 38635 62628 38669 62644
rect 37886 62550 37902 62584
rect 38078 62550 38094 62584
rect 38384 62550 38400 62584
rect 38576 62550 38592 62584
rect 38635 62578 38669 62594
rect 37730 62490 37760 62532
rect 37670 62360 37760 62490
rect 38730 62532 38738 62690
rect 38730 62490 38760 62532
rect 38800 62490 38820 62730
rect 38730 62360 38820 62490
rect 42660 63050 42750 63170
rect 42660 62790 42680 63050
rect 42720 63000 42750 63050
rect 42740 62842 42750 63000
rect 43720 63050 43810 63170
rect 43720 63000 43750 63050
rect 42808 62938 42842 62954
rect 42876 62948 42892 62982
rect 43068 62948 43084 62982
rect 43374 62948 43390 62982
rect 43566 62948 43582 62982
rect 42808 62888 42842 62904
rect 43625 62938 43659 62954
rect 42876 62860 42892 62894
rect 43068 62860 43084 62894
rect 43374 62860 43390 62894
rect 43566 62860 43582 62894
rect 43625 62888 43659 62904
rect 42720 62790 42750 62842
rect 42660 62730 42750 62790
rect 42660 62490 42680 62730
rect 42720 62690 42750 62730
rect 42740 62532 42750 62690
rect 43720 62842 43728 63000
rect 43720 62810 43750 62842
rect 43790 62810 43810 63050
rect 43720 62730 43810 62810
rect 43720 62690 43750 62730
rect 42808 62628 42842 62644
rect 42876 62638 42892 62672
rect 43068 62638 43084 62672
rect 43374 62638 43390 62672
rect 43566 62638 43582 62672
rect 42808 62578 42842 62594
rect 43625 62628 43659 62644
rect 42876 62550 42892 62584
rect 43068 62550 43084 62584
rect 43374 62550 43390 62584
rect 43566 62550 43582 62584
rect 43625 62578 43659 62594
rect 42720 62490 42750 62532
rect 42660 62360 42750 62490
rect 43720 62532 43728 62690
rect 43720 62490 43750 62532
rect 43790 62490 43810 62730
rect 43720 62360 43810 62490
rect 47650 63050 47740 63170
rect 47650 62790 47670 63050
rect 47710 63000 47740 63050
rect 47730 62842 47740 63000
rect 48710 63050 48800 63170
rect 48710 63000 48740 63050
rect 47798 62938 47832 62954
rect 47866 62948 47882 62982
rect 48058 62948 48074 62982
rect 48364 62948 48380 62982
rect 48556 62948 48572 62982
rect 47798 62888 47832 62904
rect 48615 62938 48649 62954
rect 47866 62860 47882 62894
rect 48058 62860 48074 62894
rect 48364 62860 48380 62894
rect 48556 62860 48572 62894
rect 48615 62888 48649 62904
rect 47710 62790 47740 62842
rect 47650 62730 47740 62790
rect 47650 62490 47670 62730
rect 47710 62690 47740 62730
rect 47730 62532 47740 62690
rect 48710 62842 48718 63000
rect 48710 62810 48740 62842
rect 48780 62810 48800 63050
rect 48710 62730 48800 62810
rect 48710 62690 48740 62730
rect 47798 62628 47832 62644
rect 47866 62638 47882 62672
rect 48058 62638 48074 62672
rect 48364 62638 48380 62672
rect 48556 62638 48572 62672
rect 47798 62578 47832 62594
rect 48615 62628 48649 62644
rect 47866 62550 47882 62584
rect 48058 62550 48074 62584
rect 48364 62550 48380 62584
rect 48556 62550 48572 62584
rect 48615 62578 48649 62594
rect 47710 62490 47740 62532
rect 47650 62360 47740 62490
rect 48710 62532 48718 62690
rect 48710 62490 48740 62532
rect 48780 62490 48800 62730
rect 48710 62360 48800 62490
rect 52640 63050 52730 63170
rect 52640 62790 52660 63050
rect 52700 63000 52730 63050
rect 52720 62842 52730 63000
rect 53700 63050 53790 63170
rect 53700 63000 53730 63050
rect 52788 62938 52822 62954
rect 52856 62948 52872 62982
rect 53048 62948 53064 62982
rect 53354 62948 53370 62982
rect 53546 62948 53562 62982
rect 52788 62888 52822 62904
rect 53605 62938 53639 62954
rect 52856 62860 52872 62894
rect 53048 62860 53064 62894
rect 53354 62860 53370 62894
rect 53546 62860 53562 62894
rect 53605 62888 53639 62904
rect 52700 62790 52730 62842
rect 52640 62730 52730 62790
rect 52640 62490 52660 62730
rect 52700 62690 52730 62730
rect 52720 62532 52730 62690
rect 53700 62842 53708 63000
rect 53700 62810 53730 62842
rect 53770 62810 53790 63050
rect 53700 62730 53790 62810
rect 53700 62690 53730 62730
rect 52788 62628 52822 62644
rect 52856 62638 52872 62672
rect 53048 62638 53064 62672
rect 53354 62638 53370 62672
rect 53546 62638 53562 62672
rect 52788 62578 52822 62594
rect 53605 62628 53639 62644
rect 52856 62550 52872 62584
rect 53048 62550 53064 62584
rect 53354 62550 53370 62584
rect 53546 62550 53562 62584
rect 53605 62578 53639 62594
rect 52700 62490 52730 62532
rect 52640 62360 52730 62490
rect 53700 62532 53708 62690
rect 53700 62490 53730 62532
rect 53770 62490 53790 62730
rect 53700 62360 53790 62490
rect 57630 63050 57720 63170
rect 57630 62790 57650 63050
rect 57690 63000 57720 63050
rect 57710 62842 57720 63000
rect 58690 63050 58780 63170
rect 58690 63000 58720 63050
rect 57778 62938 57812 62954
rect 57846 62948 57862 62982
rect 58038 62948 58054 62982
rect 58344 62948 58360 62982
rect 58536 62948 58552 62982
rect 57778 62888 57812 62904
rect 58595 62938 58629 62954
rect 57846 62860 57862 62894
rect 58038 62860 58054 62894
rect 58344 62860 58360 62894
rect 58536 62860 58552 62894
rect 58595 62888 58629 62904
rect 57690 62790 57720 62842
rect 57630 62730 57720 62790
rect 57630 62490 57650 62730
rect 57690 62690 57720 62730
rect 57710 62532 57720 62690
rect 58690 62842 58698 63000
rect 58690 62810 58720 62842
rect 58760 62810 58780 63050
rect 58690 62730 58780 62810
rect 58690 62690 58720 62730
rect 57778 62628 57812 62644
rect 57846 62638 57862 62672
rect 58038 62638 58054 62672
rect 58344 62638 58360 62672
rect 58536 62638 58552 62672
rect 57778 62578 57812 62594
rect 58595 62628 58629 62644
rect 57846 62550 57862 62584
rect 58038 62550 58054 62584
rect 58344 62550 58360 62584
rect 58536 62550 58552 62584
rect 58595 62578 58629 62594
rect 57690 62490 57720 62532
rect 57630 62360 57720 62490
rect 58690 62532 58698 62690
rect 58690 62490 58720 62532
rect 58760 62490 58780 62730
rect 58690 62360 58780 62490
rect 62620 63050 62710 63170
rect 62620 62790 62640 63050
rect 62680 63000 62710 63050
rect 62700 62842 62710 63000
rect 63680 63050 63770 63170
rect 63680 63000 63710 63050
rect 62768 62938 62802 62954
rect 62836 62948 62852 62982
rect 63028 62948 63044 62982
rect 63334 62948 63350 62982
rect 63526 62948 63542 62982
rect 62768 62888 62802 62904
rect 63585 62938 63619 62954
rect 62836 62860 62852 62894
rect 63028 62860 63044 62894
rect 63334 62860 63350 62894
rect 63526 62860 63542 62894
rect 63585 62888 63619 62904
rect 62680 62790 62710 62842
rect 62620 62730 62710 62790
rect 62620 62490 62640 62730
rect 62680 62690 62710 62730
rect 62700 62532 62710 62690
rect 63680 62842 63688 63000
rect 63680 62810 63710 62842
rect 63750 62810 63770 63050
rect 63680 62730 63770 62810
rect 63680 62690 63710 62730
rect 62768 62628 62802 62644
rect 62836 62638 62852 62672
rect 63028 62638 63044 62672
rect 63334 62638 63350 62672
rect 63526 62638 63542 62672
rect 62768 62578 62802 62594
rect 63585 62628 63619 62644
rect 62836 62550 62852 62584
rect 63028 62550 63044 62584
rect 63334 62550 63350 62584
rect 63526 62550 63542 62584
rect 63585 62578 63619 62594
rect 62680 62490 62710 62532
rect 62620 62360 62710 62490
rect 63680 62532 63688 62690
rect 63680 62490 63710 62532
rect 63750 62490 63770 62730
rect 63680 62360 63770 62490
rect 67610 63050 67700 63170
rect 67610 62790 67630 63050
rect 67670 63000 67700 63050
rect 67690 62842 67700 63000
rect 68670 63050 68760 63170
rect 68670 63000 68700 63050
rect 67758 62938 67792 62954
rect 67826 62948 67842 62982
rect 68018 62948 68034 62982
rect 68324 62948 68340 62982
rect 68516 62948 68532 62982
rect 67758 62888 67792 62904
rect 68575 62938 68609 62954
rect 67826 62860 67842 62894
rect 68018 62860 68034 62894
rect 68324 62860 68340 62894
rect 68516 62860 68532 62894
rect 68575 62888 68609 62904
rect 67670 62790 67700 62842
rect 67610 62730 67700 62790
rect 67610 62490 67630 62730
rect 67670 62690 67700 62730
rect 67690 62532 67700 62690
rect 68670 62842 68678 63000
rect 68670 62810 68700 62842
rect 68740 62810 68760 63050
rect 68670 62730 68760 62810
rect 68670 62690 68700 62730
rect 67758 62628 67792 62644
rect 67826 62638 67842 62672
rect 68018 62638 68034 62672
rect 68324 62638 68340 62672
rect 68516 62638 68532 62672
rect 67758 62578 67792 62594
rect 68575 62628 68609 62644
rect 67826 62550 67842 62584
rect 68018 62550 68034 62584
rect 68324 62550 68340 62584
rect 68516 62550 68532 62584
rect 68575 62578 68609 62594
rect 67670 62490 67700 62532
rect 67610 62360 67700 62490
rect 68670 62532 68678 62690
rect 68670 62490 68700 62532
rect 68740 62490 68760 62730
rect 68670 62360 68760 62490
rect 72600 63050 72690 63170
rect 72600 62790 72620 63050
rect 72660 63000 72690 63050
rect 72680 62842 72690 63000
rect 73660 63050 73750 63170
rect 73660 63000 73690 63050
rect 72748 62938 72782 62954
rect 72816 62948 72832 62982
rect 73008 62948 73024 62982
rect 73314 62948 73330 62982
rect 73506 62948 73522 62982
rect 72748 62888 72782 62904
rect 73565 62938 73599 62954
rect 72816 62860 72832 62894
rect 73008 62860 73024 62894
rect 73314 62860 73330 62894
rect 73506 62860 73522 62894
rect 73565 62888 73599 62904
rect 72660 62790 72690 62842
rect 72600 62730 72690 62790
rect 72600 62490 72620 62730
rect 72660 62690 72690 62730
rect 72680 62532 72690 62690
rect 73660 62842 73668 63000
rect 73660 62810 73690 62842
rect 73730 62810 73750 63050
rect 73660 62730 73750 62810
rect 73660 62690 73690 62730
rect 72748 62628 72782 62644
rect 72816 62638 72832 62672
rect 73008 62638 73024 62672
rect 73314 62638 73330 62672
rect 73506 62638 73522 62672
rect 72748 62578 72782 62594
rect 73565 62628 73599 62644
rect 72816 62550 72832 62584
rect 73008 62550 73024 62584
rect 73314 62550 73330 62584
rect 73506 62550 73522 62584
rect 73565 62578 73599 62594
rect 72660 62490 72690 62532
rect 72600 62360 72690 62490
rect 73660 62532 73668 62690
rect 73660 62490 73690 62532
rect 73730 62490 73750 62730
rect 73660 62360 73750 62490
rect 77590 63050 77680 63170
rect 77590 62790 77610 63050
rect 77650 63000 77680 63050
rect 77670 62842 77680 63000
rect 78650 63050 78740 63170
rect 78650 63000 78680 63050
rect 77738 62938 77772 62954
rect 77806 62948 77822 62982
rect 77998 62948 78014 62982
rect 78304 62948 78320 62982
rect 78496 62948 78512 62982
rect 77738 62888 77772 62904
rect 78555 62938 78589 62954
rect 77806 62860 77822 62894
rect 77998 62860 78014 62894
rect 78304 62860 78320 62894
rect 78496 62860 78512 62894
rect 78555 62888 78589 62904
rect 77650 62790 77680 62842
rect 77590 62730 77680 62790
rect 77590 62490 77610 62730
rect 77650 62690 77680 62730
rect 77670 62532 77680 62690
rect 78650 62842 78658 63000
rect 78650 62810 78680 62842
rect 78720 62810 78740 63050
rect 78650 62730 78740 62810
rect 78650 62690 78680 62730
rect 77738 62628 77772 62644
rect 77806 62638 77822 62672
rect 77998 62638 78014 62672
rect 78304 62638 78320 62672
rect 78496 62638 78512 62672
rect 77738 62578 77772 62594
rect 78555 62628 78589 62644
rect 77806 62550 77822 62584
rect 77998 62550 78014 62584
rect 78304 62550 78320 62584
rect 78496 62550 78512 62584
rect 78555 62578 78589 62594
rect 77650 62490 77680 62532
rect 77590 62360 77680 62490
rect 78650 62532 78658 62690
rect 78650 62490 78680 62532
rect 78720 62490 78740 62730
rect 78650 62360 78740 62490
rect 2740 61340 2830 61460
rect 2740 61080 2760 61340
rect 2800 61290 2830 61340
rect 2820 61132 2830 61290
rect 3800 61340 3890 61460
rect 3800 61290 3830 61340
rect 2888 61228 2922 61244
rect 2956 61238 2972 61272
rect 3148 61238 3164 61272
rect 3454 61238 3470 61272
rect 3646 61238 3662 61272
rect 2888 61178 2922 61194
rect 3705 61228 3739 61244
rect 2956 61150 2972 61184
rect 3148 61150 3164 61184
rect 3454 61150 3470 61184
rect 3646 61150 3662 61184
rect 3705 61178 3739 61194
rect 2800 61080 2830 61132
rect 2740 61020 2830 61080
rect 2740 60780 2760 61020
rect 2800 60980 2830 61020
rect 2820 60822 2830 60980
rect 3800 61132 3808 61290
rect 3800 61100 3830 61132
rect 3870 61100 3890 61340
rect 3800 61020 3890 61100
rect 3800 60980 3830 61020
rect 2888 60918 2922 60934
rect 2956 60928 2972 60962
rect 3148 60928 3164 60962
rect 3454 60928 3470 60962
rect 3646 60928 3662 60962
rect 2888 60868 2922 60884
rect 3705 60918 3739 60934
rect 2956 60840 2972 60874
rect 3148 60840 3164 60874
rect 3454 60840 3470 60874
rect 3646 60840 3662 60874
rect 3705 60868 3739 60884
rect 2800 60780 2830 60822
rect 2740 60650 2830 60780
rect 3800 60822 3808 60980
rect 3800 60780 3830 60822
rect 3870 60780 3890 61020
rect 3800 60650 3890 60780
rect 7730 61340 7820 61460
rect 7730 61080 7750 61340
rect 7790 61290 7820 61340
rect 7810 61132 7820 61290
rect 8790 61340 8880 61460
rect 8790 61290 8820 61340
rect 7878 61228 7912 61244
rect 7946 61238 7962 61272
rect 8138 61238 8154 61272
rect 8444 61238 8460 61272
rect 8636 61238 8652 61272
rect 7878 61178 7912 61194
rect 8695 61228 8729 61244
rect 7946 61150 7962 61184
rect 8138 61150 8154 61184
rect 8444 61150 8460 61184
rect 8636 61150 8652 61184
rect 8695 61178 8729 61194
rect 7790 61080 7820 61132
rect 7730 61020 7820 61080
rect 7730 60780 7750 61020
rect 7790 60980 7820 61020
rect 7810 60822 7820 60980
rect 8790 61132 8798 61290
rect 8790 61100 8820 61132
rect 8860 61100 8880 61340
rect 8790 61020 8880 61100
rect 8790 60980 8820 61020
rect 7878 60918 7912 60934
rect 7946 60928 7962 60962
rect 8138 60928 8154 60962
rect 8444 60928 8460 60962
rect 8636 60928 8652 60962
rect 7878 60868 7912 60884
rect 8695 60918 8729 60934
rect 7946 60840 7962 60874
rect 8138 60840 8154 60874
rect 8444 60840 8460 60874
rect 8636 60840 8652 60874
rect 8695 60868 8729 60884
rect 7790 60780 7820 60822
rect 7730 60650 7820 60780
rect 8790 60822 8798 60980
rect 8790 60780 8820 60822
rect 8860 60780 8880 61020
rect 8790 60650 8880 60780
rect 12720 61340 12810 61460
rect 12720 61080 12740 61340
rect 12780 61290 12810 61340
rect 12800 61132 12810 61290
rect 13780 61340 13870 61460
rect 13780 61290 13810 61340
rect 12868 61228 12902 61244
rect 12936 61238 12952 61272
rect 13128 61238 13144 61272
rect 13434 61238 13450 61272
rect 13626 61238 13642 61272
rect 12868 61178 12902 61194
rect 13685 61228 13719 61244
rect 12936 61150 12952 61184
rect 13128 61150 13144 61184
rect 13434 61150 13450 61184
rect 13626 61150 13642 61184
rect 13685 61178 13719 61194
rect 12780 61080 12810 61132
rect 12720 61020 12810 61080
rect 12720 60780 12740 61020
rect 12780 60980 12810 61020
rect 12800 60822 12810 60980
rect 13780 61132 13788 61290
rect 13780 61100 13810 61132
rect 13850 61100 13870 61340
rect 13780 61020 13870 61100
rect 13780 60980 13810 61020
rect 12868 60918 12902 60934
rect 12936 60928 12952 60962
rect 13128 60928 13144 60962
rect 13434 60928 13450 60962
rect 13626 60928 13642 60962
rect 12868 60868 12902 60884
rect 13685 60918 13719 60934
rect 12936 60840 12952 60874
rect 13128 60840 13144 60874
rect 13434 60840 13450 60874
rect 13626 60840 13642 60874
rect 13685 60868 13719 60884
rect 12780 60780 12810 60822
rect 12720 60650 12810 60780
rect 13780 60822 13788 60980
rect 13780 60780 13810 60822
rect 13850 60780 13870 61020
rect 13780 60650 13870 60780
rect 17710 61340 17800 61460
rect 17710 61080 17730 61340
rect 17770 61290 17800 61340
rect 17790 61132 17800 61290
rect 18770 61340 18860 61460
rect 18770 61290 18800 61340
rect 17858 61228 17892 61244
rect 17926 61238 17942 61272
rect 18118 61238 18134 61272
rect 18424 61238 18440 61272
rect 18616 61238 18632 61272
rect 17858 61178 17892 61194
rect 18675 61228 18709 61244
rect 17926 61150 17942 61184
rect 18118 61150 18134 61184
rect 18424 61150 18440 61184
rect 18616 61150 18632 61184
rect 18675 61178 18709 61194
rect 17770 61080 17800 61132
rect 17710 61020 17800 61080
rect 17710 60780 17730 61020
rect 17770 60980 17800 61020
rect 17790 60822 17800 60980
rect 18770 61132 18778 61290
rect 18770 61100 18800 61132
rect 18840 61100 18860 61340
rect 18770 61020 18860 61100
rect 18770 60980 18800 61020
rect 17858 60918 17892 60934
rect 17926 60928 17942 60962
rect 18118 60928 18134 60962
rect 18424 60928 18440 60962
rect 18616 60928 18632 60962
rect 17858 60868 17892 60884
rect 18675 60918 18709 60934
rect 17926 60840 17942 60874
rect 18118 60840 18134 60874
rect 18424 60840 18440 60874
rect 18616 60840 18632 60874
rect 18675 60868 18709 60884
rect 17770 60780 17800 60822
rect 17710 60650 17800 60780
rect 18770 60822 18778 60980
rect 18770 60780 18800 60822
rect 18840 60780 18860 61020
rect 18770 60650 18860 60780
rect 22700 61340 22790 61460
rect 22700 61080 22720 61340
rect 22760 61290 22790 61340
rect 22780 61132 22790 61290
rect 23760 61340 23850 61460
rect 23760 61290 23790 61340
rect 22848 61228 22882 61244
rect 22916 61238 22932 61272
rect 23108 61238 23124 61272
rect 23414 61238 23430 61272
rect 23606 61238 23622 61272
rect 22848 61178 22882 61194
rect 23665 61228 23699 61244
rect 22916 61150 22932 61184
rect 23108 61150 23124 61184
rect 23414 61150 23430 61184
rect 23606 61150 23622 61184
rect 23665 61178 23699 61194
rect 22760 61080 22790 61132
rect 22700 61020 22790 61080
rect 22700 60780 22720 61020
rect 22760 60980 22790 61020
rect 22780 60822 22790 60980
rect 23760 61132 23768 61290
rect 23760 61100 23790 61132
rect 23830 61100 23850 61340
rect 23760 61020 23850 61100
rect 23760 60980 23790 61020
rect 22848 60918 22882 60934
rect 22916 60928 22932 60962
rect 23108 60928 23124 60962
rect 23414 60928 23430 60962
rect 23606 60928 23622 60962
rect 22848 60868 22882 60884
rect 23665 60918 23699 60934
rect 22916 60840 22932 60874
rect 23108 60840 23124 60874
rect 23414 60840 23430 60874
rect 23606 60840 23622 60874
rect 23665 60868 23699 60884
rect 22760 60780 22790 60822
rect 22700 60650 22790 60780
rect 23760 60822 23768 60980
rect 23760 60780 23790 60822
rect 23830 60780 23850 61020
rect 23760 60650 23850 60780
rect 27690 61340 27780 61460
rect 27690 61080 27710 61340
rect 27750 61290 27780 61340
rect 27770 61132 27780 61290
rect 28750 61340 28840 61460
rect 28750 61290 28780 61340
rect 27838 61228 27872 61244
rect 27906 61238 27922 61272
rect 28098 61238 28114 61272
rect 28404 61238 28420 61272
rect 28596 61238 28612 61272
rect 27838 61178 27872 61194
rect 28655 61228 28689 61244
rect 27906 61150 27922 61184
rect 28098 61150 28114 61184
rect 28404 61150 28420 61184
rect 28596 61150 28612 61184
rect 28655 61178 28689 61194
rect 27750 61080 27780 61132
rect 27690 61020 27780 61080
rect 27690 60780 27710 61020
rect 27750 60980 27780 61020
rect 27770 60822 27780 60980
rect 28750 61132 28758 61290
rect 28750 61100 28780 61132
rect 28820 61100 28840 61340
rect 28750 61020 28840 61100
rect 28750 60980 28780 61020
rect 27838 60918 27872 60934
rect 27906 60928 27922 60962
rect 28098 60928 28114 60962
rect 28404 60928 28420 60962
rect 28596 60928 28612 60962
rect 27838 60868 27872 60884
rect 28655 60918 28689 60934
rect 27906 60840 27922 60874
rect 28098 60840 28114 60874
rect 28404 60840 28420 60874
rect 28596 60840 28612 60874
rect 28655 60868 28689 60884
rect 27750 60780 27780 60822
rect 27690 60650 27780 60780
rect 28750 60822 28758 60980
rect 28750 60780 28780 60822
rect 28820 60780 28840 61020
rect 28750 60650 28840 60780
rect 32680 61340 32770 61460
rect 32680 61080 32700 61340
rect 32740 61290 32770 61340
rect 32760 61132 32770 61290
rect 33740 61340 33830 61460
rect 33740 61290 33770 61340
rect 32828 61228 32862 61244
rect 32896 61238 32912 61272
rect 33088 61238 33104 61272
rect 33394 61238 33410 61272
rect 33586 61238 33602 61272
rect 32828 61178 32862 61194
rect 33645 61228 33679 61244
rect 32896 61150 32912 61184
rect 33088 61150 33104 61184
rect 33394 61150 33410 61184
rect 33586 61150 33602 61184
rect 33645 61178 33679 61194
rect 32740 61080 32770 61132
rect 32680 61020 32770 61080
rect 32680 60780 32700 61020
rect 32740 60980 32770 61020
rect 32760 60822 32770 60980
rect 33740 61132 33748 61290
rect 33740 61100 33770 61132
rect 33810 61100 33830 61340
rect 33740 61020 33830 61100
rect 33740 60980 33770 61020
rect 32828 60918 32862 60934
rect 32896 60928 32912 60962
rect 33088 60928 33104 60962
rect 33394 60928 33410 60962
rect 33586 60928 33602 60962
rect 32828 60868 32862 60884
rect 33645 60918 33679 60934
rect 32896 60840 32912 60874
rect 33088 60840 33104 60874
rect 33394 60840 33410 60874
rect 33586 60840 33602 60874
rect 33645 60868 33679 60884
rect 32740 60780 32770 60822
rect 32680 60650 32770 60780
rect 33740 60822 33748 60980
rect 33740 60780 33770 60822
rect 33810 60780 33830 61020
rect 33740 60650 33830 60780
rect 37670 61340 37760 61460
rect 37670 61080 37690 61340
rect 37730 61290 37760 61340
rect 37750 61132 37760 61290
rect 38730 61340 38820 61460
rect 38730 61290 38760 61340
rect 37818 61228 37852 61244
rect 37886 61238 37902 61272
rect 38078 61238 38094 61272
rect 38384 61238 38400 61272
rect 38576 61238 38592 61272
rect 37818 61178 37852 61194
rect 38635 61228 38669 61244
rect 37886 61150 37902 61184
rect 38078 61150 38094 61184
rect 38384 61150 38400 61184
rect 38576 61150 38592 61184
rect 38635 61178 38669 61194
rect 37730 61080 37760 61132
rect 37670 61020 37760 61080
rect 37670 60780 37690 61020
rect 37730 60980 37760 61020
rect 37750 60822 37760 60980
rect 38730 61132 38738 61290
rect 38730 61100 38760 61132
rect 38800 61100 38820 61340
rect 38730 61020 38820 61100
rect 38730 60980 38760 61020
rect 37818 60918 37852 60934
rect 37886 60928 37902 60962
rect 38078 60928 38094 60962
rect 38384 60928 38400 60962
rect 38576 60928 38592 60962
rect 37818 60868 37852 60884
rect 38635 60918 38669 60934
rect 37886 60840 37902 60874
rect 38078 60840 38094 60874
rect 38384 60840 38400 60874
rect 38576 60840 38592 60874
rect 38635 60868 38669 60884
rect 37730 60780 37760 60822
rect 37670 60650 37760 60780
rect 38730 60822 38738 60980
rect 38730 60780 38760 60822
rect 38800 60780 38820 61020
rect 38730 60650 38820 60780
rect 42660 61340 42750 61460
rect 42660 61080 42680 61340
rect 42720 61290 42750 61340
rect 42740 61132 42750 61290
rect 43720 61340 43810 61460
rect 43720 61290 43750 61340
rect 42808 61228 42842 61244
rect 42876 61238 42892 61272
rect 43068 61238 43084 61272
rect 43374 61238 43390 61272
rect 43566 61238 43582 61272
rect 42808 61178 42842 61194
rect 43625 61228 43659 61244
rect 42876 61150 42892 61184
rect 43068 61150 43084 61184
rect 43374 61150 43390 61184
rect 43566 61150 43582 61184
rect 43625 61178 43659 61194
rect 42720 61080 42750 61132
rect 42660 61020 42750 61080
rect 42660 60780 42680 61020
rect 42720 60980 42750 61020
rect 42740 60822 42750 60980
rect 43720 61132 43728 61290
rect 43720 61100 43750 61132
rect 43790 61100 43810 61340
rect 43720 61020 43810 61100
rect 43720 60980 43750 61020
rect 42808 60918 42842 60934
rect 42876 60928 42892 60962
rect 43068 60928 43084 60962
rect 43374 60928 43390 60962
rect 43566 60928 43582 60962
rect 42808 60868 42842 60884
rect 43625 60918 43659 60934
rect 42876 60840 42892 60874
rect 43068 60840 43084 60874
rect 43374 60840 43390 60874
rect 43566 60840 43582 60874
rect 43625 60868 43659 60884
rect 42720 60780 42750 60822
rect 42660 60650 42750 60780
rect 43720 60822 43728 60980
rect 43720 60780 43750 60822
rect 43790 60780 43810 61020
rect 43720 60650 43810 60780
rect 47650 61340 47740 61460
rect 47650 61080 47670 61340
rect 47710 61290 47740 61340
rect 47730 61132 47740 61290
rect 48710 61340 48800 61460
rect 48710 61290 48740 61340
rect 47798 61228 47832 61244
rect 47866 61238 47882 61272
rect 48058 61238 48074 61272
rect 48364 61238 48380 61272
rect 48556 61238 48572 61272
rect 47798 61178 47832 61194
rect 48615 61228 48649 61244
rect 47866 61150 47882 61184
rect 48058 61150 48074 61184
rect 48364 61150 48380 61184
rect 48556 61150 48572 61184
rect 48615 61178 48649 61194
rect 47710 61080 47740 61132
rect 47650 61020 47740 61080
rect 47650 60780 47670 61020
rect 47710 60980 47740 61020
rect 47730 60822 47740 60980
rect 48710 61132 48718 61290
rect 48710 61100 48740 61132
rect 48780 61100 48800 61340
rect 48710 61020 48800 61100
rect 48710 60980 48740 61020
rect 47798 60918 47832 60934
rect 47866 60928 47882 60962
rect 48058 60928 48074 60962
rect 48364 60928 48380 60962
rect 48556 60928 48572 60962
rect 47798 60868 47832 60884
rect 48615 60918 48649 60934
rect 47866 60840 47882 60874
rect 48058 60840 48074 60874
rect 48364 60840 48380 60874
rect 48556 60840 48572 60874
rect 48615 60868 48649 60884
rect 47710 60780 47740 60822
rect 47650 60650 47740 60780
rect 48710 60822 48718 60980
rect 48710 60780 48740 60822
rect 48780 60780 48800 61020
rect 48710 60650 48800 60780
rect 52640 61340 52730 61460
rect 52640 61080 52660 61340
rect 52700 61290 52730 61340
rect 52720 61132 52730 61290
rect 53700 61340 53790 61460
rect 53700 61290 53730 61340
rect 52788 61228 52822 61244
rect 52856 61238 52872 61272
rect 53048 61238 53064 61272
rect 53354 61238 53370 61272
rect 53546 61238 53562 61272
rect 52788 61178 52822 61194
rect 53605 61228 53639 61244
rect 52856 61150 52872 61184
rect 53048 61150 53064 61184
rect 53354 61150 53370 61184
rect 53546 61150 53562 61184
rect 53605 61178 53639 61194
rect 52700 61080 52730 61132
rect 52640 61020 52730 61080
rect 52640 60780 52660 61020
rect 52700 60980 52730 61020
rect 52720 60822 52730 60980
rect 53700 61132 53708 61290
rect 53700 61100 53730 61132
rect 53770 61100 53790 61340
rect 53700 61020 53790 61100
rect 53700 60980 53730 61020
rect 52788 60918 52822 60934
rect 52856 60928 52872 60962
rect 53048 60928 53064 60962
rect 53354 60928 53370 60962
rect 53546 60928 53562 60962
rect 52788 60868 52822 60884
rect 53605 60918 53639 60934
rect 52856 60840 52872 60874
rect 53048 60840 53064 60874
rect 53354 60840 53370 60874
rect 53546 60840 53562 60874
rect 53605 60868 53639 60884
rect 52700 60780 52730 60822
rect 52640 60650 52730 60780
rect 53700 60822 53708 60980
rect 53700 60780 53730 60822
rect 53770 60780 53790 61020
rect 53700 60650 53790 60780
rect 57630 61340 57720 61460
rect 57630 61080 57650 61340
rect 57690 61290 57720 61340
rect 57710 61132 57720 61290
rect 58690 61340 58780 61460
rect 58690 61290 58720 61340
rect 57778 61228 57812 61244
rect 57846 61238 57862 61272
rect 58038 61238 58054 61272
rect 58344 61238 58360 61272
rect 58536 61238 58552 61272
rect 57778 61178 57812 61194
rect 58595 61228 58629 61244
rect 57846 61150 57862 61184
rect 58038 61150 58054 61184
rect 58344 61150 58360 61184
rect 58536 61150 58552 61184
rect 58595 61178 58629 61194
rect 57690 61080 57720 61132
rect 57630 61020 57720 61080
rect 57630 60780 57650 61020
rect 57690 60980 57720 61020
rect 57710 60822 57720 60980
rect 58690 61132 58698 61290
rect 58690 61100 58720 61132
rect 58760 61100 58780 61340
rect 58690 61020 58780 61100
rect 58690 60980 58720 61020
rect 57778 60918 57812 60934
rect 57846 60928 57862 60962
rect 58038 60928 58054 60962
rect 58344 60928 58360 60962
rect 58536 60928 58552 60962
rect 57778 60868 57812 60884
rect 58595 60918 58629 60934
rect 57846 60840 57862 60874
rect 58038 60840 58054 60874
rect 58344 60840 58360 60874
rect 58536 60840 58552 60874
rect 58595 60868 58629 60884
rect 57690 60780 57720 60822
rect 57630 60650 57720 60780
rect 58690 60822 58698 60980
rect 58690 60780 58720 60822
rect 58760 60780 58780 61020
rect 58690 60650 58780 60780
rect 62620 61340 62710 61460
rect 62620 61080 62640 61340
rect 62680 61290 62710 61340
rect 62700 61132 62710 61290
rect 63680 61340 63770 61460
rect 63680 61290 63710 61340
rect 62768 61228 62802 61244
rect 62836 61238 62852 61272
rect 63028 61238 63044 61272
rect 63334 61238 63350 61272
rect 63526 61238 63542 61272
rect 62768 61178 62802 61194
rect 63585 61228 63619 61244
rect 62836 61150 62852 61184
rect 63028 61150 63044 61184
rect 63334 61150 63350 61184
rect 63526 61150 63542 61184
rect 63585 61178 63619 61194
rect 62680 61080 62710 61132
rect 62620 61020 62710 61080
rect 62620 60780 62640 61020
rect 62680 60980 62710 61020
rect 62700 60822 62710 60980
rect 63680 61132 63688 61290
rect 63680 61100 63710 61132
rect 63750 61100 63770 61340
rect 63680 61020 63770 61100
rect 63680 60980 63710 61020
rect 62768 60918 62802 60934
rect 62836 60928 62852 60962
rect 63028 60928 63044 60962
rect 63334 60928 63350 60962
rect 63526 60928 63542 60962
rect 62768 60868 62802 60884
rect 63585 60918 63619 60934
rect 62836 60840 62852 60874
rect 63028 60840 63044 60874
rect 63334 60840 63350 60874
rect 63526 60840 63542 60874
rect 63585 60868 63619 60884
rect 62680 60780 62710 60822
rect 62620 60650 62710 60780
rect 63680 60822 63688 60980
rect 63680 60780 63710 60822
rect 63750 60780 63770 61020
rect 63680 60650 63770 60780
rect 67610 61340 67700 61460
rect 67610 61080 67630 61340
rect 67670 61290 67700 61340
rect 67690 61132 67700 61290
rect 68670 61340 68760 61460
rect 68670 61290 68700 61340
rect 67758 61228 67792 61244
rect 67826 61238 67842 61272
rect 68018 61238 68034 61272
rect 68324 61238 68340 61272
rect 68516 61238 68532 61272
rect 67758 61178 67792 61194
rect 68575 61228 68609 61244
rect 67826 61150 67842 61184
rect 68018 61150 68034 61184
rect 68324 61150 68340 61184
rect 68516 61150 68532 61184
rect 68575 61178 68609 61194
rect 67670 61080 67700 61132
rect 67610 61020 67700 61080
rect 67610 60780 67630 61020
rect 67670 60980 67700 61020
rect 67690 60822 67700 60980
rect 68670 61132 68678 61290
rect 68670 61100 68700 61132
rect 68740 61100 68760 61340
rect 68670 61020 68760 61100
rect 68670 60980 68700 61020
rect 67758 60918 67792 60934
rect 67826 60928 67842 60962
rect 68018 60928 68034 60962
rect 68324 60928 68340 60962
rect 68516 60928 68532 60962
rect 67758 60868 67792 60884
rect 68575 60918 68609 60934
rect 67826 60840 67842 60874
rect 68018 60840 68034 60874
rect 68324 60840 68340 60874
rect 68516 60840 68532 60874
rect 68575 60868 68609 60884
rect 67670 60780 67700 60822
rect 67610 60650 67700 60780
rect 68670 60822 68678 60980
rect 68670 60780 68700 60822
rect 68740 60780 68760 61020
rect 68670 60650 68760 60780
rect 72600 61340 72690 61460
rect 72600 61080 72620 61340
rect 72660 61290 72690 61340
rect 72680 61132 72690 61290
rect 73660 61340 73750 61460
rect 73660 61290 73690 61340
rect 72748 61228 72782 61244
rect 72816 61238 72832 61272
rect 73008 61238 73024 61272
rect 73314 61238 73330 61272
rect 73506 61238 73522 61272
rect 72748 61178 72782 61194
rect 73565 61228 73599 61244
rect 72816 61150 72832 61184
rect 73008 61150 73024 61184
rect 73314 61150 73330 61184
rect 73506 61150 73522 61184
rect 73565 61178 73599 61194
rect 72660 61080 72690 61132
rect 72600 61020 72690 61080
rect 72600 60780 72620 61020
rect 72660 60980 72690 61020
rect 72680 60822 72690 60980
rect 73660 61132 73668 61290
rect 73660 61100 73690 61132
rect 73730 61100 73750 61340
rect 73660 61020 73750 61100
rect 73660 60980 73690 61020
rect 72748 60918 72782 60934
rect 72816 60928 72832 60962
rect 73008 60928 73024 60962
rect 73314 60928 73330 60962
rect 73506 60928 73522 60962
rect 72748 60868 72782 60884
rect 73565 60918 73599 60934
rect 72816 60840 72832 60874
rect 73008 60840 73024 60874
rect 73314 60840 73330 60874
rect 73506 60840 73522 60874
rect 73565 60868 73599 60884
rect 72660 60780 72690 60822
rect 72600 60650 72690 60780
rect 73660 60822 73668 60980
rect 73660 60780 73690 60822
rect 73730 60780 73750 61020
rect 73660 60650 73750 60780
rect 77590 61340 77680 61460
rect 77590 61080 77610 61340
rect 77650 61290 77680 61340
rect 77670 61132 77680 61290
rect 78650 61340 78740 61460
rect 78650 61290 78680 61340
rect 77738 61228 77772 61244
rect 77806 61238 77822 61272
rect 77998 61238 78014 61272
rect 78304 61238 78320 61272
rect 78496 61238 78512 61272
rect 77738 61178 77772 61194
rect 78555 61228 78589 61244
rect 77806 61150 77822 61184
rect 77998 61150 78014 61184
rect 78304 61150 78320 61184
rect 78496 61150 78512 61184
rect 78555 61178 78589 61194
rect 77650 61080 77680 61132
rect 77590 61020 77680 61080
rect 77590 60780 77610 61020
rect 77650 60980 77680 61020
rect 77670 60822 77680 60980
rect 78650 61132 78658 61290
rect 78650 61100 78680 61132
rect 78720 61100 78740 61340
rect 78650 61020 78740 61100
rect 78650 60980 78680 61020
rect 77738 60918 77772 60934
rect 77806 60928 77822 60962
rect 77998 60928 78014 60962
rect 78304 60928 78320 60962
rect 78496 60928 78512 60962
rect 77738 60868 77772 60884
rect 78555 60918 78589 60934
rect 77806 60840 77822 60874
rect 77998 60840 78014 60874
rect 78304 60840 78320 60874
rect 78496 60840 78512 60874
rect 78555 60868 78589 60884
rect 77650 60780 77680 60822
rect 77590 60650 77680 60780
rect 78650 60822 78658 60980
rect 78650 60780 78680 60822
rect 78720 60780 78740 61020
rect 78650 60650 78740 60780
rect 2740 59630 2830 59750
rect 2740 59370 2760 59630
rect 2800 59580 2830 59630
rect 2820 59422 2830 59580
rect 3800 59630 3890 59750
rect 3800 59580 3830 59630
rect 2888 59518 2922 59534
rect 2956 59528 2972 59562
rect 3148 59528 3164 59562
rect 3454 59528 3470 59562
rect 3646 59528 3662 59562
rect 2888 59468 2922 59484
rect 3705 59518 3739 59534
rect 2956 59440 2972 59474
rect 3148 59440 3164 59474
rect 3454 59440 3470 59474
rect 3646 59440 3662 59474
rect 3705 59468 3739 59484
rect 2800 59370 2830 59422
rect 2740 59310 2830 59370
rect 2740 59070 2760 59310
rect 2800 59270 2830 59310
rect 2820 59112 2830 59270
rect 3800 59422 3808 59580
rect 3800 59390 3830 59422
rect 3870 59390 3890 59630
rect 3800 59310 3890 59390
rect 3800 59270 3830 59310
rect 2888 59208 2922 59224
rect 2956 59218 2972 59252
rect 3148 59218 3164 59252
rect 3454 59218 3470 59252
rect 3646 59218 3662 59252
rect 2888 59158 2922 59174
rect 3705 59208 3739 59224
rect 2956 59130 2972 59164
rect 3148 59130 3164 59164
rect 3454 59130 3470 59164
rect 3646 59130 3662 59164
rect 3705 59158 3739 59174
rect 2800 59070 2830 59112
rect 2740 58940 2830 59070
rect 3800 59112 3808 59270
rect 3800 59070 3830 59112
rect 3870 59070 3890 59310
rect 3800 58940 3890 59070
rect 7730 59630 7820 59750
rect 7730 59370 7750 59630
rect 7790 59580 7820 59630
rect 7810 59422 7820 59580
rect 8790 59630 8880 59750
rect 8790 59580 8820 59630
rect 7878 59518 7912 59534
rect 7946 59528 7962 59562
rect 8138 59528 8154 59562
rect 8444 59528 8460 59562
rect 8636 59528 8652 59562
rect 7878 59468 7912 59484
rect 8695 59518 8729 59534
rect 7946 59440 7962 59474
rect 8138 59440 8154 59474
rect 8444 59440 8460 59474
rect 8636 59440 8652 59474
rect 8695 59468 8729 59484
rect 7790 59370 7820 59422
rect 7730 59310 7820 59370
rect 7730 59070 7750 59310
rect 7790 59270 7820 59310
rect 7810 59112 7820 59270
rect 8790 59422 8798 59580
rect 8790 59390 8820 59422
rect 8860 59390 8880 59630
rect 8790 59310 8880 59390
rect 8790 59270 8820 59310
rect 7878 59208 7912 59224
rect 7946 59218 7962 59252
rect 8138 59218 8154 59252
rect 8444 59218 8460 59252
rect 8636 59218 8652 59252
rect 7878 59158 7912 59174
rect 8695 59208 8729 59224
rect 7946 59130 7962 59164
rect 8138 59130 8154 59164
rect 8444 59130 8460 59164
rect 8636 59130 8652 59164
rect 8695 59158 8729 59174
rect 7790 59070 7820 59112
rect 7730 58940 7820 59070
rect 8790 59112 8798 59270
rect 8790 59070 8820 59112
rect 8860 59070 8880 59310
rect 8790 58940 8880 59070
rect 12720 59630 12810 59750
rect 12720 59370 12740 59630
rect 12780 59580 12810 59630
rect 12800 59422 12810 59580
rect 13780 59630 13870 59750
rect 13780 59580 13810 59630
rect 12868 59518 12902 59534
rect 12936 59528 12952 59562
rect 13128 59528 13144 59562
rect 13434 59528 13450 59562
rect 13626 59528 13642 59562
rect 12868 59468 12902 59484
rect 13685 59518 13719 59534
rect 12936 59440 12952 59474
rect 13128 59440 13144 59474
rect 13434 59440 13450 59474
rect 13626 59440 13642 59474
rect 13685 59468 13719 59484
rect 12780 59370 12810 59422
rect 12720 59310 12810 59370
rect 12720 59070 12740 59310
rect 12780 59270 12810 59310
rect 12800 59112 12810 59270
rect 13780 59422 13788 59580
rect 13780 59390 13810 59422
rect 13850 59390 13870 59630
rect 13780 59310 13870 59390
rect 13780 59270 13810 59310
rect 12868 59208 12902 59224
rect 12936 59218 12952 59252
rect 13128 59218 13144 59252
rect 13434 59218 13450 59252
rect 13626 59218 13642 59252
rect 12868 59158 12902 59174
rect 13685 59208 13719 59224
rect 12936 59130 12952 59164
rect 13128 59130 13144 59164
rect 13434 59130 13450 59164
rect 13626 59130 13642 59164
rect 13685 59158 13719 59174
rect 12780 59070 12810 59112
rect 12720 58940 12810 59070
rect 13780 59112 13788 59270
rect 13780 59070 13810 59112
rect 13850 59070 13870 59310
rect 13780 58940 13870 59070
rect 17710 59630 17800 59750
rect 17710 59370 17730 59630
rect 17770 59580 17800 59630
rect 17790 59422 17800 59580
rect 18770 59630 18860 59750
rect 18770 59580 18800 59630
rect 17858 59518 17892 59534
rect 17926 59528 17942 59562
rect 18118 59528 18134 59562
rect 18424 59528 18440 59562
rect 18616 59528 18632 59562
rect 17858 59468 17892 59484
rect 18675 59518 18709 59534
rect 17926 59440 17942 59474
rect 18118 59440 18134 59474
rect 18424 59440 18440 59474
rect 18616 59440 18632 59474
rect 18675 59468 18709 59484
rect 17770 59370 17800 59422
rect 17710 59310 17800 59370
rect 17710 59070 17730 59310
rect 17770 59270 17800 59310
rect 17790 59112 17800 59270
rect 18770 59422 18778 59580
rect 18770 59390 18800 59422
rect 18840 59390 18860 59630
rect 18770 59310 18860 59390
rect 18770 59270 18800 59310
rect 17858 59208 17892 59224
rect 17926 59218 17942 59252
rect 18118 59218 18134 59252
rect 18424 59218 18440 59252
rect 18616 59218 18632 59252
rect 17858 59158 17892 59174
rect 18675 59208 18709 59224
rect 17926 59130 17942 59164
rect 18118 59130 18134 59164
rect 18424 59130 18440 59164
rect 18616 59130 18632 59164
rect 18675 59158 18709 59174
rect 17770 59070 17800 59112
rect 17710 58940 17800 59070
rect 18770 59112 18778 59270
rect 18770 59070 18800 59112
rect 18840 59070 18860 59310
rect 18770 58940 18860 59070
rect 22700 59630 22790 59750
rect 22700 59370 22720 59630
rect 22760 59580 22790 59630
rect 22780 59422 22790 59580
rect 23760 59630 23850 59750
rect 23760 59580 23790 59630
rect 22848 59518 22882 59534
rect 22916 59528 22932 59562
rect 23108 59528 23124 59562
rect 23414 59528 23430 59562
rect 23606 59528 23622 59562
rect 22848 59468 22882 59484
rect 23665 59518 23699 59534
rect 22916 59440 22932 59474
rect 23108 59440 23124 59474
rect 23414 59440 23430 59474
rect 23606 59440 23622 59474
rect 23665 59468 23699 59484
rect 22760 59370 22790 59422
rect 22700 59310 22790 59370
rect 22700 59070 22720 59310
rect 22760 59270 22790 59310
rect 22780 59112 22790 59270
rect 23760 59422 23768 59580
rect 23760 59390 23790 59422
rect 23830 59390 23850 59630
rect 23760 59310 23850 59390
rect 23760 59270 23790 59310
rect 22848 59208 22882 59224
rect 22916 59218 22932 59252
rect 23108 59218 23124 59252
rect 23414 59218 23430 59252
rect 23606 59218 23622 59252
rect 22848 59158 22882 59174
rect 23665 59208 23699 59224
rect 22916 59130 22932 59164
rect 23108 59130 23124 59164
rect 23414 59130 23430 59164
rect 23606 59130 23622 59164
rect 23665 59158 23699 59174
rect 22760 59070 22790 59112
rect 22700 58940 22790 59070
rect 23760 59112 23768 59270
rect 23760 59070 23790 59112
rect 23830 59070 23850 59310
rect 23760 58940 23850 59070
rect 27690 59630 27780 59750
rect 27690 59370 27710 59630
rect 27750 59580 27780 59630
rect 27770 59422 27780 59580
rect 28750 59630 28840 59750
rect 28750 59580 28780 59630
rect 27838 59518 27872 59534
rect 27906 59528 27922 59562
rect 28098 59528 28114 59562
rect 28404 59528 28420 59562
rect 28596 59528 28612 59562
rect 27838 59468 27872 59484
rect 28655 59518 28689 59534
rect 27906 59440 27922 59474
rect 28098 59440 28114 59474
rect 28404 59440 28420 59474
rect 28596 59440 28612 59474
rect 28655 59468 28689 59484
rect 27750 59370 27780 59422
rect 27690 59310 27780 59370
rect 27690 59070 27710 59310
rect 27750 59270 27780 59310
rect 27770 59112 27780 59270
rect 28750 59422 28758 59580
rect 28750 59390 28780 59422
rect 28820 59390 28840 59630
rect 28750 59310 28840 59390
rect 28750 59270 28780 59310
rect 27838 59208 27872 59224
rect 27906 59218 27922 59252
rect 28098 59218 28114 59252
rect 28404 59218 28420 59252
rect 28596 59218 28612 59252
rect 27838 59158 27872 59174
rect 28655 59208 28689 59224
rect 27906 59130 27922 59164
rect 28098 59130 28114 59164
rect 28404 59130 28420 59164
rect 28596 59130 28612 59164
rect 28655 59158 28689 59174
rect 27750 59070 27780 59112
rect 27690 58940 27780 59070
rect 28750 59112 28758 59270
rect 28750 59070 28780 59112
rect 28820 59070 28840 59310
rect 28750 58940 28840 59070
rect 32680 59630 32770 59750
rect 32680 59370 32700 59630
rect 32740 59580 32770 59630
rect 32760 59422 32770 59580
rect 33740 59630 33830 59750
rect 33740 59580 33770 59630
rect 32828 59518 32862 59534
rect 32896 59528 32912 59562
rect 33088 59528 33104 59562
rect 33394 59528 33410 59562
rect 33586 59528 33602 59562
rect 32828 59468 32862 59484
rect 33645 59518 33679 59534
rect 32896 59440 32912 59474
rect 33088 59440 33104 59474
rect 33394 59440 33410 59474
rect 33586 59440 33602 59474
rect 33645 59468 33679 59484
rect 32740 59370 32770 59422
rect 32680 59310 32770 59370
rect 32680 59070 32700 59310
rect 32740 59270 32770 59310
rect 32760 59112 32770 59270
rect 33740 59422 33748 59580
rect 33740 59390 33770 59422
rect 33810 59390 33830 59630
rect 33740 59310 33830 59390
rect 33740 59270 33770 59310
rect 32828 59208 32862 59224
rect 32896 59218 32912 59252
rect 33088 59218 33104 59252
rect 33394 59218 33410 59252
rect 33586 59218 33602 59252
rect 32828 59158 32862 59174
rect 33645 59208 33679 59224
rect 32896 59130 32912 59164
rect 33088 59130 33104 59164
rect 33394 59130 33410 59164
rect 33586 59130 33602 59164
rect 33645 59158 33679 59174
rect 32740 59070 32770 59112
rect 32680 58940 32770 59070
rect 33740 59112 33748 59270
rect 33740 59070 33770 59112
rect 33810 59070 33830 59310
rect 33740 58940 33830 59070
rect 37670 59630 37760 59750
rect 37670 59370 37690 59630
rect 37730 59580 37760 59630
rect 37750 59422 37760 59580
rect 38730 59630 38820 59750
rect 38730 59580 38760 59630
rect 37818 59518 37852 59534
rect 37886 59528 37902 59562
rect 38078 59528 38094 59562
rect 38384 59528 38400 59562
rect 38576 59528 38592 59562
rect 37818 59468 37852 59484
rect 38635 59518 38669 59534
rect 37886 59440 37902 59474
rect 38078 59440 38094 59474
rect 38384 59440 38400 59474
rect 38576 59440 38592 59474
rect 38635 59468 38669 59484
rect 37730 59370 37760 59422
rect 37670 59310 37760 59370
rect 37670 59070 37690 59310
rect 37730 59270 37760 59310
rect 37750 59112 37760 59270
rect 38730 59422 38738 59580
rect 38730 59390 38760 59422
rect 38800 59390 38820 59630
rect 38730 59310 38820 59390
rect 38730 59270 38760 59310
rect 37818 59208 37852 59224
rect 37886 59218 37902 59252
rect 38078 59218 38094 59252
rect 38384 59218 38400 59252
rect 38576 59218 38592 59252
rect 37818 59158 37852 59174
rect 38635 59208 38669 59224
rect 37886 59130 37902 59164
rect 38078 59130 38094 59164
rect 38384 59130 38400 59164
rect 38576 59130 38592 59164
rect 38635 59158 38669 59174
rect 37730 59070 37760 59112
rect 37670 58940 37760 59070
rect 38730 59112 38738 59270
rect 38730 59070 38760 59112
rect 38800 59070 38820 59310
rect 38730 58940 38820 59070
rect 42660 59630 42750 59750
rect 42660 59370 42680 59630
rect 42720 59580 42750 59630
rect 42740 59422 42750 59580
rect 43720 59630 43810 59750
rect 43720 59580 43750 59630
rect 42808 59518 42842 59534
rect 42876 59528 42892 59562
rect 43068 59528 43084 59562
rect 43374 59528 43390 59562
rect 43566 59528 43582 59562
rect 42808 59468 42842 59484
rect 43625 59518 43659 59534
rect 42876 59440 42892 59474
rect 43068 59440 43084 59474
rect 43374 59440 43390 59474
rect 43566 59440 43582 59474
rect 43625 59468 43659 59484
rect 42720 59370 42750 59422
rect 42660 59310 42750 59370
rect 42660 59070 42680 59310
rect 42720 59270 42750 59310
rect 42740 59112 42750 59270
rect 43720 59422 43728 59580
rect 43720 59390 43750 59422
rect 43790 59390 43810 59630
rect 43720 59310 43810 59390
rect 43720 59270 43750 59310
rect 42808 59208 42842 59224
rect 42876 59218 42892 59252
rect 43068 59218 43084 59252
rect 43374 59218 43390 59252
rect 43566 59218 43582 59252
rect 42808 59158 42842 59174
rect 43625 59208 43659 59224
rect 42876 59130 42892 59164
rect 43068 59130 43084 59164
rect 43374 59130 43390 59164
rect 43566 59130 43582 59164
rect 43625 59158 43659 59174
rect 42720 59070 42750 59112
rect 42660 58940 42750 59070
rect 43720 59112 43728 59270
rect 43720 59070 43750 59112
rect 43790 59070 43810 59310
rect 43720 58940 43810 59070
rect 47650 59630 47740 59750
rect 47650 59370 47670 59630
rect 47710 59580 47740 59630
rect 47730 59422 47740 59580
rect 48710 59630 48800 59750
rect 48710 59580 48740 59630
rect 47798 59518 47832 59534
rect 47866 59528 47882 59562
rect 48058 59528 48074 59562
rect 48364 59528 48380 59562
rect 48556 59528 48572 59562
rect 47798 59468 47832 59484
rect 48615 59518 48649 59534
rect 47866 59440 47882 59474
rect 48058 59440 48074 59474
rect 48364 59440 48380 59474
rect 48556 59440 48572 59474
rect 48615 59468 48649 59484
rect 47710 59370 47740 59422
rect 47650 59310 47740 59370
rect 47650 59070 47670 59310
rect 47710 59270 47740 59310
rect 47730 59112 47740 59270
rect 48710 59422 48718 59580
rect 48710 59390 48740 59422
rect 48780 59390 48800 59630
rect 48710 59310 48800 59390
rect 48710 59270 48740 59310
rect 47798 59208 47832 59224
rect 47866 59218 47882 59252
rect 48058 59218 48074 59252
rect 48364 59218 48380 59252
rect 48556 59218 48572 59252
rect 47798 59158 47832 59174
rect 48615 59208 48649 59224
rect 47866 59130 47882 59164
rect 48058 59130 48074 59164
rect 48364 59130 48380 59164
rect 48556 59130 48572 59164
rect 48615 59158 48649 59174
rect 47710 59070 47740 59112
rect 47650 58940 47740 59070
rect 48710 59112 48718 59270
rect 48710 59070 48740 59112
rect 48780 59070 48800 59310
rect 48710 58940 48800 59070
rect 52640 59630 52730 59750
rect 52640 59370 52660 59630
rect 52700 59580 52730 59630
rect 52720 59422 52730 59580
rect 53700 59630 53790 59750
rect 53700 59580 53730 59630
rect 52788 59518 52822 59534
rect 52856 59528 52872 59562
rect 53048 59528 53064 59562
rect 53354 59528 53370 59562
rect 53546 59528 53562 59562
rect 52788 59468 52822 59484
rect 53605 59518 53639 59534
rect 52856 59440 52872 59474
rect 53048 59440 53064 59474
rect 53354 59440 53370 59474
rect 53546 59440 53562 59474
rect 53605 59468 53639 59484
rect 52700 59370 52730 59422
rect 52640 59310 52730 59370
rect 52640 59070 52660 59310
rect 52700 59270 52730 59310
rect 52720 59112 52730 59270
rect 53700 59422 53708 59580
rect 53700 59390 53730 59422
rect 53770 59390 53790 59630
rect 53700 59310 53790 59390
rect 53700 59270 53730 59310
rect 52788 59208 52822 59224
rect 52856 59218 52872 59252
rect 53048 59218 53064 59252
rect 53354 59218 53370 59252
rect 53546 59218 53562 59252
rect 52788 59158 52822 59174
rect 53605 59208 53639 59224
rect 52856 59130 52872 59164
rect 53048 59130 53064 59164
rect 53354 59130 53370 59164
rect 53546 59130 53562 59164
rect 53605 59158 53639 59174
rect 52700 59070 52730 59112
rect 52640 58940 52730 59070
rect 53700 59112 53708 59270
rect 53700 59070 53730 59112
rect 53770 59070 53790 59310
rect 53700 58940 53790 59070
rect 57630 59630 57720 59750
rect 57630 59370 57650 59630
rect 57690 59580 57720 59630
rect 57710 59422 57720 59580
rect 58690 59630 58780 59750
rect 58690 59580 58720 59630
rect 57778 59518 57812 59534
rect 57846 59528 57862 59562
rect 58038 59528 58054 59562
rect 58344 59528 58360 59562
rect 58536 59528 58552 59562
rect 57778 59468 57812 59484
rect 58595 59518 58629 59534
rect 57846 59440 57862 59474
rect 58038 59440 58054 59474
rect 58344 59440 58360 59474
rect 58536 59440 58552 59474
rect 58595 59468 58629 59484
rect 57690 59370 57720 59422
rect 57630 59310 57720 59370
rect 57630 59070 57650 59310
rect 57690 59270 57720 59310
rect 57710 59112 57720 59270
rect 58690 59422 58698 59580
rect 58690 59390 58720 59422
rect 58760 59390 58780 59630
rect 58690 59310 58780 59390
rect 58690 59270 58720 59310
rect 57778 59208 57812 59224
rect 57846 59218 57862 59252
rect 58038 59218 58054 59252
rect 58344 59218 58360 59252
rect 58536 59218 58552 59252
rect 57778 59158 57812 59174
rect 58595 59208 58629 59224
rect 57846 59130 57862 59164
rect 58038 59130 58054 59164
rect 58344 59130 58360 59164
rect 58536 59130 58552 59164
rect 58595 59158 58629 59174
rect 57690 59070 57720 59112
rect 57630 58940 57720 59070
rect 58690 59112 58698 59270
rect 58690 59070 58720 59112
rect 58760 59070 58780 59310
rect 58690 58940 58780 59070
rect 62620 59630 62710 59750
rect 62620 59370 62640 59630
rect 62680 59580 62710 59630
rect 62700 59422 62710 59580
rect 63680 59630 63770 59750
rect 63680 59580 63710 59630
rect 62768 59518 62802 59534
rect 62836 59528 62852 59562
rect 63028 59528 63044 59562
rect 63334 59528 63350 59562
rect 63526 59528 63542 59562
rect 62768 59468 62802 59484
rect 63585 59518 63619 59534
rect 62836 59440 62852 59474
rect 63028 59440 63044 59474
rect 63334 59440 63350 59474
rect 63526 59440 63542 59474
rect 63585 59468 63619 59484
rect 62680 59370 62710 59422
rect 62620 59310 62710 59370
rect 62620 59070 62640 59310
rect 62680 59270 62710 59310
rect 62700 59112 62710 59270
rect 63680 59422 63688 59580
rect 63680 59390 63710 59422
rect 63750 59390 63770 59630
rect 63680 59310 63770 59390
rect 63680 59270 63710 59310
rect 62768 59208 62802 59224
rect 62836 59218 62852 59252
rect 63028 59218 63044 59252
rect 63334 59218 63350 59252
rect 63526 59218 63542 59252
rect 62768 59158 62802 59174
rect 63585 59208 63619 59224
rect 62836 59130 62852 59164
rect 63028 59130 63044 59164
rect 63334 59130 63350 59164
rect 63526 59130 63542 59164
rect 63585 59158 63619 59174
rect 62680 59070 62710 59112
rect 62620 58940 62710 59070
rect 63680 59112 63688 59270
rect 63680 59070 63710 59112
rect 63750 59070 63770 59310
rect 63680 58940 63770 59070
rect 67610 59630 67700 59750
rect 67610 59370 67630 59630
rect 67670 59580 67700 59630
rect 67690 59422 67700 59580
rect 68670 59630 68760 59750
rect 68670 59580 68700 59630
rect 67758 59518 67792 59534
rect 67826 59528 67842 59562
rect 68018 59528 68034 59562
rect 68324 59528 68340 59562
rect 68516 59528 68532 59562
rect 67758 59468 67792 59484
rect 68575 59518 68609 59534
rect 67826 59440 67842 59474
rect 68018 59440 68034 59474
rect 68324 59440 68340 59474
rect 68516 59440 68532 59474
rect 68575 59468 68609 59484
rect 67670 59370 67700 59422
rect 67610 59310 67700 59370
rect 67610 59070 67630 59310
rect 67670 59270 67700 59310
rect 67690 59112 67700 59270
rect 68670 59422 68678 59580
rect 68670 59390 68700 59422
rect 68740 59390 68760 59630
rect 68670 59310 68760 59390
rect 68670 59270 68700 59310
rect 67758 59208 67792 59224
rect 67826 59218 67842 59252
rect 68018 59218 68034 59252
rect 68324 59218 68340 59252
rect 68516 59218 68532 59252
rect 67758 59158 67792 59174
rect 68575 59208 68609 59224
rect 67826 59130 67842 59164
rect 68018 59130 68034 59164
rect 68324 59130 68340 59164
rect 68516 59130 68532 59164
rect 68575 59158 68609 59174
rect 67670 59070 67700 59112
rect 67610 58940 67700 59070
rect 68670 59112 68678 59270
rect 68670 59070 68700 59112
rect 68740 59070 68760 59310
rect 68670 58940 68760 59070
rect 72600 59630 72690 59750
rect 72600 59370 72620 59630
rect 72660 59580 72690 59630
rect 72680 59422 72690 59580
rect 73660 59630 73750 59750
rect 73660 59580 73690 59630
rect 72748 59518 72782 59534
rect 72816 59528 72832 59562
rect 73008 59528 73024 59562
rect 73314 59528 73330 59562
rect 73506 59528 73522 59562
rect 72748 59468 72782 59484
rect 73565 59518 73599 59534
rect 72816 59440 72832 59474
rect 73008 59440 73024 59474
rect 73314 59440 73330 59474
rect 73506 59440 73522 59474
rect 73565 59468 73599 59484
rect 72660 59370 72690 59422
rect 72600 59310 72690 59370
rect 72600 59070 72620 59310
rect 72660 59270 72690 59310
rect 72680 59112 72690 59270
rect 73660 59422 73668 59580
rect 73660 59390 73690 59422
rect 73730 59390 73750 59630
rect 73660 59310 73750 59390
rect 73660 59270 73690 59310
rect 72748 59208 72782 59224
rect 72816 59218 72832 59252
rect 73008 59218 73024 59252
rect 73314 59218 73330 59252
rect 73506 59218 73522 59252
rect 72748 59158 72782 59174
rect 73565 59208 73599 59224
rect 72816 59130 72832 59164
rect 73008 59130 73024 59164
rect 73314 59130 73330 59164
rect 73506 59130 73522 59164
rect 73565 59158 73599 59174
rect 72660 59070 72690 59112
rect 72600 58940 72690 59070
rect 73660 59112 73668 59270
rect 73660 59070 73690 59112
rect 73730 59070 73750 59310
rect 73660 58940 73750 59070
rect 77590 59630 77680 59750
rect 77590 59370 77610 59630
rect 77650 59580 77680 59630
rect 77670 59422 77680 59580
rect 78650 59630 78740 59750
rect 78650 59580 78680 59630
rect 77738 59518 77772 59534
rect 77806 59528 77822 59562
rect 77998 59528 78014 59562
rect 78304 59528 78320 59562
rect 78496 59528 78512 59562
rect 77738 59468 77772 59484
rect 78555 59518 78589 59534
rect 77806 59440 77822 59474
rect 77998 59440 78014 59474
rect 78304 59440 78320 59474
rect 78496 59440 78512 59474
rect 78555 59468 78589 59484
rect 77650 59370 77680 59422
rect 77590 59310 77680 59370
rect 77590 59070 77610 59310
rect 77650 59270 77680 59310
rect 77670 59112 77680 59270
rect 78650 59422 78658 59580
rect 78650 59390 78680 59422
rect 78720 59390 78740 59630
rect 78650 59310 78740 59390
rect 78650 59270 78680 59310
rect 77738 59208 77772 59224
rect 77806 59218 77822 59252
rect 77998 59218 78014 59252
rect 78304 59218 78320 59252
rect 78496 59218 78512 59252
rect 77738 59158 77772 59174
rect 78555 59208 78589 59224
rect 77806 59130 77822 59164
rect 77998 59130 78014 59164
rect 78304 59130 78320 59164
rect 78496 59130 78512 59164
rect 78555 59158 78589 59174
rect 77650 59070 77680 59112
rect 77590 58940 77680 59070
rect 78650 59112 78658 59270
rect 78650 59070 78680 59112
rect 78720 59070 78740 59310
rect 78650 58940 78740 59070
rect 2740 57920 2830 58040
rect 2740 57660 2760 57920
rect 2800 57870 2830 57920
rect 2820 57712 2830 57870
rect 3800 57920 3890 58040
rect 3800 57870 3830 57920
rect 2888 57808 2922 57824
rect 2956 57818 2972 57852
rect 3148 57818 3164 57852
rect 3454 57818 3470 57852
rect 3646 57818 3662 57852
rect 2888 57758 2922 57774
rect 3705 57808 3739 57824
rect 2956 57730 2972 57764
rect 3148 57730 3164 57764
rect 3454 57730 3470 57764
rect 3646 57730 3662 57764
rect 3705 57758 3739 57774
rect 2800 57660 2830 57712
rect 2740 57600 2830 57660
rect 2740 57360 2760 57600
rect 2800 57560 2830 57600
rect 2820 57402 2830 57560
rect 3800 57712 3808 57870
rect 3800 57680 3830 57712
rect 3870 57680 3890 57920
rect 3800 57600 3890 57680
rect 3800 57560 3830 57600
rect 2888 57498 2922 57514
rect 2956 57508 2972 57542
rect 3148 57508 3164 57542
rect 3454 57508 3470 57542
rect 3646 57508 3662 57542
rect 2888 57448 2922 57464
rect 3705 57498 3739 57514
rect 2956 57420 2972 57454
rect 3148 57420 3164 57454
rect 3454 57420 3470 57454
rect 3646 57420 3662 57454
rect 3705 57448 3739 57464
rect 2800 57360 2830 57402
rect 2740 57230 2830 57360
rect 3800 57402 3808 57560
rect 3800 57360 3830 57402
rect 3870 57360 3890 57600
rect 3800 57230 3890 57360
rect 7730 57920 7820 58040
rect 7730 57660 7750 57920
rect 7790 57870 7820 57920
rect 7810 57712 7820 57870
rect 8790 57920 8880 58040
rect 8790 57870 8820 57920
rect 7878 57808 7912 57824
rect 7946 57818 7962 57852
rect 8138 57818 8154 57852
rect 8444 57818 8460 57852
rect 8636 57818 8652 57852
rect 7878 57758 7912 57774
rect 8695 57808 8729 57824
rect 7946 57730 7962 57764
rect 8138 57730 8154 57764
rect 8444 57730 8460 57764
rect 8636 57730 8652 57764
rect 8695 57758 8729 57774
rect 7790 57660 7820 57712
rect 7730 57600 7820 57660
rect 7730 57360 7750 57600
rect 7790 57560 7820 57600
rect 7810 57402 7820 57560
rect 8790 57712 8798 57870
rect 8790 57680 8820 57712
rect 8860 57680 8880 57920
rect 8790 57600 8880 57680
rect 8790 57560 8820 57600
rect 7878 57498 7912 57514
rect 7946 57508 7962 57542
rect 8138 57508 8154 57542
rect 8444 57508 8460 57542
rect 8636 57508 8652 57542
rect 7878 57448 7912 57464
rect 8695 57498 8729 57514
rect 7946 57420 7962 57454
rect 8138 57420 8154 57454
rect 8444 57420 8460 57454
rect 8636 57420 8652 57454
rect 8695 57448 8729 57464
rect 7790 57360 7820 57402
rect 7730 57230 7820 57360
rect 8790 57402 8798 57560
rect 8790 57360 8820 57402
rect 8860 57360 8880 57600
rect 8790 57230 8880 57360
rect 12720 57920 12810 58040
rect 12720 57660 12740 57920
rect 12780 57870 12810 57920
rect 12800 57712 12810 57870
rect 13780 57920 13870 58040
rect 13780 57870 13810 57920
rect 12868 57808 12902 57824
rect 12936 57818 12952 57852
rect 13128 57818 13144 57852
rect 13434 57818 13450 57852
rect 13626 57818 13642 57852
rect 12868 57758 12902 57774
rect 13685 57808 13719 57824
rect 12936 57730 12952 57764
rect 13128 57730 13144 57764
rect 13434 57730 13450 57764
rect 13626 57730 13642 57764
rect 13685 57758 13719 57774
rect 12780 57660 12810 57712
rect 12720 57600 12810 57660
rect 12720 57360 12740 57600
rect 12780 57560 12810 57600
rect 12800 57402 12810 57560
rect 13780 57712 13788 57870
rect 13780 57680 13810 57712
rect 13850 57680 13870 57920
rect 13780 57600 13870 57680
rect 13780 57560 13810 57600
rect 12868 57498 12902 57514
rect 12936 57508 12952 57542
rect 13128 57508 13144 57542
rect 13434 57508 13450 57542
rect 13626 57508 13642 57542
rect 12868 57448 12902 57464
rect 13685 57498 13719 57514
rect 12936 57420 12952 57454
rect 13128 57420 13144 57454
rect 13434 57420 13450 57454
rect 13626 57420 13642 57454
rect 13685 57448 13719 57464
rect 12780 57360 12810 57402
rect 12720 57230 12810 57360
rect 13780 57402 13788 57560
rect 13780 57360 13810 57402
rect 13850 57360 13870 57600
rect 13780 57230 13870 57360
rect 17710 57920 17800 58040
rect 17710 57660 17730 57920
rect 17770 57870 17800 57920
rect 17790 57712 17800 57870
rect 18770 57920 18860 58040
rect 18770 57870 18800 57920
rect 17858 57808 17892 57824
rect 17926 57818 17942 57852
rect 18118 57818 18134 57852
rect 18424 57818 18440 57852
rect 18616 57818 18632 57852
rect 17858 57758 17892 57774
rect 18675 57808 18709 57824
rect 17926 57730 17942 57764
rect 18118 57730 18134 57764
rect 18424 57730 18440 57764
rect 18616 57730 18632 57764
rect 18675 57758 18709 57774
rect 17770 57660 17800 57712
rect 17710 57600 17800 57660
rect 17710 57360 17730 57600
rect 17770 57560 17800 57600
rect 17790 57402 17800 57560
rect 18770 57712 18778 57870
rect 18770 57680 18800 57712
rect 18840 57680 18860 57920
rect 18770 57600 18860 57680
rect 18770 57560 18800 57600
rect 17858 57498 17892 57514
rect 17926 57508 17942 57542
rect 18118 57508 18134 57542
rect 18424 57508 18440 57542
rect 18616 57508 18632 57542
rect 17858 57448 17892 57464
rect 18675 57498 18709 57514
rect 17926 57420 17942 57454
rect 18118 57420 18134 57454
rect 18424 57420 18440 57454
rect 18616 57420 18632 57454
rect 18675 57448 18709 57464
rect 17770 57360 17800 57402
rect 17710 57230 17800 57360
rect 18770 57402 18778 57560
rect 18770 57360 18800 57402
rect 18840 57360 18860 57600
rect 18770 57230 18860 57360
rect 22700 57920 22790 58040
rect 22700 57660 22720 57920
rect 22760 57870 22790 57920
rect 22780 57712 22790 57870
rect 23760 57920 23850 58040
rect 23760 57870 23790 57920
rect 22848 57808 22882 57824
rect 22916 57818 22932 57852
rect 23108 57818 23124 57852
rect 23414 57818 23430 57852
rect 23606 57818 23622 57852
rect 22848 57758 22882 57774
rect 23665 57808 23699 57824
rect 22916 57730 22932 57764
rect 23108 57730 23124 57764
rect 23414 57730 23430 57764
rect 23606 57730 23622 57764
rect 23665 57758 23699 57774
rect 22760 57660 22790 57712
rect 22700 57600 22790 57660
rect 22700 57360 22720 57600
rect 22760 57560 22790 57600
rect 22780 57402 22790 57560
rect 23760 57712 23768 57870
rect 23760 57680 23790 57712
rect 23830 57680 23850 57920
rect 23760 57600 23850 57680
rect 23760 57560 23790 57600
rect 22848 57498 22882 57514
rect 22916 57508 22932 57542
rect 23108 57508 23124 57542
rect 23414 57508 23430 57542
rect 23606 57508 23622 57542
rect 22848 57448 22882 57464
rect 23665 57498 23699 57514
rect 22916 57420 22932 57454
rect 23108 57420 23124 57454
rect 23414 57420 23430 57454
rect 23606 57420 23622 57454
rect 23665 57448 23699 57464
rect 22760 57360 22790 57402
rect 22700 57230 22790 57360
rect 23760 57402 23768 57560
rect 23760 57360 23790 57402
rect 23830 57360 23850 57600
rect 23760 57230 23850 57360
rect 27690 57920 27780 58040
rect 27690 57660 27710 57920
rect 27750 57870 27780 57920
rect 27770 57712 27780 57870
rect 28750 57920 28840 58040
rect 28750 57870 28780 57920
rect 27838 57808 27872 57824
rect 27906 57818 27922 57852
rect 28098 57818 28114 57852
rect 28404 57818 28420 57852
rect 28596 57818 28612 57852
rect 27838 57758 27872 57774
rect 28655 57808 28689 57824
rect 27906 57730 27922 57764
rect 28098 57730 28114 57764
rect 28404 57730 28420 57764
rect 28596 57730 28612 57764
rect 28655 57758 28689 57774
rect 27750 57660 27780 57712
rect 27690 57600 27780 57660
rect 27690 57360 27710 57600
rect 27750 57560 27780 57600
rect 27770 57402 27780 57560
rect 28750 57712 28758 57870
rect 28750 57680 28780 57712
rect 28820 57680 28840 57920
rect 28750 57600 28840 57680
rect 28750 57560 28780 57600
rect 27838 57498 27872 57514
rect 27906 57508 27922 57542
rect 28098 57508 28114 57542
rect 28404 57508 28420 57542
rect 28596 57508 28612 57542
rect 27838 57448 27872 57464
rect 28655 57498 28689 57514
rect 27906 57420 27922 57454
rect 28098 57420 28114 57454
rect 28404 57420 28420 57454
rect 28596 57420 28612 57454
rect 28655 57448 28689 57464
rect 27750 57360 27780 57402
rect 27690 57230 27780 57360
rect 28750 57402 28758 57560
rect 28750 57360 28780 57402
rect 28820 57360 28840 57600
rect 28750 57230 28840 57360
rect 32680 57920 32770 58040
rect 32680 57660 32700 57920
rect 32740 57870 32770 57920
rect 32760 57712 32770 57870
rect 33740 57920 33830 58040
rect 33740 57870 33770 57920
rect 32828 57808 32862 57824
rect 32896 57818 32912 57852
rect 33088 57818 33104 57852
rect 33394 57818 33410 57852
rect 33586 57818 33602 57852
rect 32828 57758 32862 57774
rect 33645 57808 33679 57824
rect 32896 57730 32912 57764
rect 33088 57730 33104 57764
rect 33394 57730 33410 57764
rect 33586 57730 33602 57764
rect 33645 57758 33679 57774
rect 32740 57660 32770 57712
rect 32680 57600 32770 57660
rect 32680 57360 32700 57600
rect 32740 57560 32770 57600
rect 32760 57402 32770 57560
rect 33740 57712 33748 57870
rect 33740 57680 33770 57712
rect 33810 57680 33830 57920
rect 33740 57600 33830 57680
rect 33740 57560 33770 57600
rect 32828 57498 32862 57514
rect 32896 57508 32912 57542
rect 33088 57508 33104 57542
rect 33394 57508 33410 57542
rect 33586 57508 33602 57542
rect 32828 57448 32862 57464
rect 33645 57498 33679 57514
rect 32896 57420 32912 57454
rect 33088 57420 33104 57454
rect 33394 57420 33410 57454
rect 33586 57420 33602 57454
rect 33645 57448 33679 57464
rect 32740 57360 32770 57402
rect 32680 57230 32770 57360
rect 33740 57402 33748 57560
rect 33740 57360 33770 57402
rect 33810 57360 33830 57600
rect 33740 57230 33830 57360
rect 37670 57920 37760 58040
rect 37670 57660 37690 57920
rect 37730 57870 37760 57920
rect 37750 57712 37760 57870
rect 38730 57920 38820 58040
rect 38730 57870 38760 57920
rect 37818 57808 37852 57824
rect 37886 57818 37902 57852
rect 38078 57818 38094 57852
rect 38384 57818 38400 57852
rect 38576 57818 38592 57852
rect 37818 57758 37852 57774
rect 38635 57808 38669 57824
rect 37886 57730 37902 57764
rect 38078 57730 38094 57764
rect 38384 57730 38400 57764
rect 38576 57730 38592 57764
rect 38635 57758 38669 57774
rect 37730 57660 37760 57712
rect 37670 57600 37760 57660
rect 37670 57360 37690 57600
rect 37730 57560 37760 57600
rect 37750 57402 37760 57560
rect 38730 57712 38738 57870
rect 38730 57680 38760 57712
rect 38800 57680 38820 57920
rect 38730 57600 38820 57680
rect 38730 57560 38760 57600
rect 37818 57498 37852 57514
rect 37886 57508 37902 57542
rect 38078 57508 38094 57542
rect 38384 57508 38400 57542
rect 38576 57508 38592 57542
rect 37818 57448 37852 57464
rect 38635 57498 38669 57514
rect 37886 57420 37902 57454
rect 38078 57420 38094 57454
rect 38384 57420 38400 57454
rect 38576 57420 38592 57454
rect 38635 57448 38669 57464
rect 37730 57360 37760 57402
rect 37670 57230 37760 57360
rect 38730 57402 38738 57560
rect 38730 57360 38760 57402
rect 38800 57360 38820 57600
rect 38730 57230 38820 57360
rect 42660 57920 42750 58040
rect 42660 57660 42680 57920
rect 42720 57870 42750 57920
rect 42740 57712 42750 57870
rect 43720 57920 43810 58040
rect 43720 57870 43750 57920
rect 42808 57808 42842 57824
rect 42876 57818 42892 57852
rect 43068 57818 43084 57852
rect 43374 57818 43390 57852
rect 43566 57818 43582 57852
rect 42808 57758 42842 57774
rect 43625 57808 43659 57824
rect 42876 57730 42892 57764
rect 43068 57730 43084 57764
rect 43374 57730 43390 57764
rect 43566 57730 43582 57764
rect 43625 57758 43659 57774
rect 42720 57660 42750 57712
rect 42660 57600 42750 57660
rect 42660 57360 42680 57600
rect 42720 57560 42750 57600
rect 42740 57402 42750 57560
rect 43720 57712 43728 57870
rect 43720 57680 43750 57712
rect 43790 57680 43810 57920
rect 43720 57600 43810 57680
rect 43720 57560 43750 57600
rect 42808 57498 42842 57514
rect 42876 57508 42892 57542
rect 43068 57508 43084 57542
rect 43374 57508 43390 57542
rect 43566 57508 43582 57542
rect 42808 57448 42842 57464
rect 43625 57498 43659 57514
rect 42876 57420 42892 57454
rect 43068 57420 43084 57454
rect 43374 57420 43390 57454
rect 43566 57420 43582 57454
rect 43625 57448 43659 57464
rect 42720 57360 42750 57402
rect 42660 57230 42750 57360
rect 43720 57402 43728 57560
rect 43720 57360 43750 57402
rect 43790 57360 43810 57600
rect 43720 57230 43810 57360
rect 47650 57920 47740 58040
rect 47650 57660 47670 57920
rect 47710 57870 47740 57920
rect 47730 57712 47740 57870
rect 48710 57920 48800 58040
rect 48710 57870 48740 57920
rect 47798 57808 47832 57824
rect 47866 57818 47882 57852
rect 48058 57818 48074 57852
rect 48364 57818 48380 57852
rect 48556 57818 48572 57852
rect 47798 57758 47832 57774
rect 48615 57808 48649 57824
rect 47866 57730 47882 57764
rect 48058 57730 48074 57764
rect 48364 57730 48380 57764
rect 48556 57730 48572 57764
rect 48615 57758 48649 57774
rect 47710 57660 47740 57712
rect 47650 57600 47740 57660
rect 47650 57360 47670 57600
rect 47710 57560 47740 57600
rect 47730 57402 47740 57560
rect 48710 57712 48718 57870
rect 48710 57680 48740 57712
rect 48780 57680 48800 57920
rect 48710 57600 48800 57680
rect 48710 57560 48740 57600
rect 47798 57498 47832 57514
rect 47866 57508 47882 57542
rect 48058 57508 48074 57542
rect 48364 57508 48380 57542
rect 48556 57508 48572 57542
rect 47798 57448 47832 57464
rect 48615 57498 48649 57514
rect 47866 57420 47882 57454
rect 48058 57420 48074 57454
rect 48364 57420 48380 57454
rect 48556 57420 48572 57454
rect 48615 57448 48649 57464
rect 47710 57360 47740 57402
rect 47650 57230 47740 57360
rect 48710 57402 48718 57560
rect 48710 57360 48740 57402
rect 48780 57360 48800 57600
rect 48710 57230 48800 57360
rect 52640 57920 52730 58040
rect 52640 57660 52660 57920
rect 52700 57870 52730 57920
rect 52720 57712 52730 57870
rect 53700 57920 53790 58040
rect 53700 57870 53730 57920
rect 52788 57808 52822 57824
rect 52856 57818 52872 57852
rect 53048 57818 53064 57852
rect 53354 57818 53370 57852
rect 53546 57818 53562 57852
rect 52788 57758 52822 57774
rect 53605 57808 53639 57824
rect 52856 57730 52872 57764
rect 53048 57730 53064 57764
rect 53354 57730 53370 57764
rect 53546 57730 53562 57764
rect 53605 57758 53639 57774
rect 52700 57660 52730 57712
rect 52640 57600 52730 57660
rect 52640 57360 52660 57600
rect 52700 57560 52730 57600
rect 52720 57402 52730 57560
rect 53700 57712 53708 57870
rect 53700 57680 53730 57712
rect 53770 57680 53790 57920
rect 53700 57600 53790 57680
rect 53700 57560 53730 57600
rect 52788 57498 52822 57514
rect 52856 57508 52872 57542
rect 53048 57508 53064 57542
rect 53354 57508 53370 57542
rect 53546 57508 53562 57542
rect 52788 57448 52822 57464
rect 53605 57498 53639 57514
rect 52856 57420 52872 57454
rect 53048 57420 53064 57454
rect 53354 57420 53370 57454
rect 53546 57420 53562 57454
rect 53605 57448 53639 57464
rect 52700 57360 52730 57402
rect 52640 57230 52730 57360
rect 53700 57402 53708 57560
rect 53700 57360 53730 57402
rect 53770 57360 53790 57600
rect 53700 57230 53790 57360
rect 57630 57920 57720 58040
rect 57630 57660 57650 57920
rect 57690 57870 57720 57920
rect 57710 57712 57720 57870
rect 58690 57920 58780 58040
rect 58690 57870 58720 57920
rect 57778 57808 57812 57824
rect 57846 57818 57862 57852
rect 58038 57818 58054 57852
rect 58344 57818 58360 57852
rect 58536 57818 58552 57852
rect 57778 57758 57812 57774
rect 58595 57808 58629 57824
rect 57846 57730 57862 57764
rect 58038 57730 58054 57764
rect 58344 57730 58360 57764
rect 58536 57730 58552 57764
rect 58595 57758 58629 57774
rect 57690 57660 57720 57712
rect 57630 57600 57720 57660
rect 57630 57360 57650 57600
rect 57690 57560 57720 57600
rect 57710 57402 57720 57560
rect 58690 57712 58698 57870
rect 58690 57680 58720 57712
rect 58760 57680 58780 57920
rect 58690 57600 58780 57680
rect 58690 57560 58720 57600
rect 57778 57498 57812 57514
rect 57846 57508 57862 57542
rect 58038 57508 58054 57542
rect 58344 57508 58360 57542
rect 58536 57508 58552 57542
rect 57778 57448 57812 57464
rect 58595 57498 58629 57514
rect 57846 57420 57862 57454
rect 58038 57420 58054 57454
rect 58344 57420 58360 57454
rect 58536 57420 58552 57454
rect 58595 57448 58629 57464
rect 57690 57360 57720 57402
rect 57630 57230 57720 57360
rect 58690 57402 58698 57560
rect 58690 57360 58720 57402
rect 58760 57360 58780 57600
rect 58690 57230 58780 57360
rect 62620 57920 62710 58040
rect 62620 57660 62640 57920
rect 62680 57870 62710 57920
rect 62700 57712 62710 57870
rect 63680 57920 63770 58040
rect 63680 57870 63710 57920
rect 62768 57808 62802 57824
rect 62836 57818 62852 57852
rect 63028 57818 63044 57852
rect 63334 57818 63350 57852
rect 63526 57818 63542 57852
rect 62768 57758 62802 57774
rect 63585 57808 63619 57824
rect 62836 57730 62852 57764
rect 63028 57730 63044 57764
rect 63334 57730 63350 57764
rect 63526 57730 63542 57764
rect 63585 57758 63619 57774
rect 62680 57660 62710 57712
rect 62620 57600 62710 57660
rect 62620 57360 62640 57600
rect 62680 57560 62710 57600
rect 62700 57402 62710 57560
rect 63680 57712 63688 57870
rect 63680 57680 63710 57712
rect 63750 57680 63770 57920
rect 63680 57600 63770 57680
rect 63680 57560 63710 57600
rect 62768 57498 62802 57514
rect 62836 57508 62852 57542
rect 63028 57508 63044 57542
rect 63334 57508 63350 57542
rect 63526 57508 63542 57542
rect 62768 57448 62802 57464
rect 63585 57498 63619 57514
rect 62836 57420 62852 57454
rect 63028 57420 63044 57454
rect 63334 57420 63350 57454
rect 63526 57420 63542 57454
rect 63585 57448 63619 57464
rect 62680 57360 62710 57402
rect 62620 57230 62710 57360
rect 63680 57402 63688 57560
rect 63680 57360 63710 57402
rect 63750 57360 63770 57600
rect 63680 57230 63770 57360
rect 67610 57920 67700 58040
rect 67610 57660 67630 57920
rect 67670 57870 67700 57920
rect 67690 57712 67700 57870
rect 68670 57920 68760 58040
rect 68670 57870 68700 57920
rect 67758 57808 67792 57824
rect 67826 57818 67842 57852
rect 68018 57818 68034 57852
rect 68324 57818 68340 57852
rect 68516 57818 68532 57852
rect 67758 57758 67792 57774
rect 68575 57808 68609 57824
rect 67826 57730 67842 57764
rect 68018 57730 68034 57764
rect 68324 57730 68340 57764
rect 68516 57730 68532 57764
rect 68575 57758 68609 57774
rect 67670 57660 67700 57712
rect 67610 57600 67700 57660
rect 67610 57360 67630 57600
rect 67670 57560 67700 57600
rect 67690 57402 67700 57560
rect 68670 57712 68678 57870
rect 68670 57680 68700 57712
rect 68740 57680 68760 57920
rect 68670 57600 68760 57680
rect 68670 57560 68700 57600
rect 67758 57498 67792 57514
rect 67826 57508 67842 57542
rect 68018 57508 68034 57542
rect 68324 57508 68340 57542
rect 68516 57508 68532 57542
rect 67758 57448 67792 57464
rect 68575 57498 68609 57514
rect 67826 57420 67842 57454
rect 68018 57420 68034 57454
rect 68324 57420 68340 57454
rect 68516 57420 68532 57454
rect 68575 57448 68609 57464
rect 67670 57360 67700 57402
rect 67610 57230 67700 57360
rect 68670 57402 68678 57560
rect 68670 57360 68700 57402
rect 68740 57360 68760 57600
rect 68670 57230 68760 57360
rect 72600 57920 72690 58040
rect 72600 57660 72620 57920
rect 72660 57870 72690 57920
rect 72680 57712 72690 57870
rect 73660 57920 73750 58040
rect 73660 57870 73690 57920
rect 72748 57808 72782 57824
rect 72816 57818 72832 57852
rect 73008 57818 73024 57852
rect 73314 57818 73330 57852
rect 73506 57818 73522 57852
rect 72748 57758 72782 57774
rect 73565 57808 73599 57824
rect 72816 57730 72832 57764
rect 73008 57730 73024 57764
rect 73314 57730 73330 57764
rect 73506 57730 73522 57764
rect 73565 57758 73599 57774
rect 72660 57660 72690 57712
rect 72600 57600 72690 57660
rect 72600 57360 72620 57600
rect 72660 57560 72690 57600
rect 72680 57402 72690 57560
rect 73660 57712 73668 57870
rect 73660 57680 73690 57712
rect 73730 57680 73750 57920
rect 73660 57600 73750 57680
rect 73660 57560 73690 57600
rect 72748 57498 72782 57514
rect 72816 57508 72832 57542
rect 73008 57508 73024 57542
rect 73314 57508 73330 57542
rect 73506 57508 73522 57542
rect 72748 57448 72782 57464
rect 73565 57498 73599 57514
rect 72816 57420 72832 57454
rect 73008 57420 73024 57454
rect 73314 57420 73330 57454
rect 73506 57420 73522 57454
rect 73565 57448 73599 57464
rect 72660 57360 72690 57402
rect 72600 57230 72690 57360
rect 73660 57402 73668 57560
rect 73660 57360 73690 57402
rect 73730 57360 73750 57600
rect 73660 57230 73750 57360
rect 77590 57920 77680 58040
rect 77590 57660 77610 57920
rect 77650 57870 77680 57920
rect 77670 57712 77680 57870
rect 78650 57920 78740 58040
rect 78650 57870 78680 57920
rect 77738 57808 77772 57824
rect 77806 57818 77822 57852
rect 77998 57818 78014 57852
rect 78304 57818 78320 57852
rect 78496 57818 78512 57852
rect 77738 57758 77772 57774
rect 78555 57808 78589 57824
rect 77806 57730 77822 57764
rect 77998 57730 78014 57764
rect 78304 57730 78320 57764
rect 78496 57730 78512 57764
rect 78555 57758 78589 57774
rect 77650 57660 77680 57712
rect 77590 57600 77680 57660
rect 77590 57360 77610 57600
rect 77650 57560 77680 57600
rect 77670 57402 77680 57560
rect 78650 57712 78658 57870
rect 78650 57680 78680 57712
rect 78720 57680 78740 57920
rect 78650 57600 78740 57680
rect 78650 57560 78680 57600
rect 77738 57498 77772 57514
rect 77806 57508 77822 57542
rect 77998 57508 78014 57542
rect 78304 57508 78320 57542
rect 78496 57508 78512 57542
rect 77738 57448 77772 57464
rect 78555 57498 78589 57514
rect 77806 57420 77822 57454
rect 77998 57420 78014 57454
rect 78304 57420 78320 57454
rect 78496 57420 78512 57454
rect 78555 57448 78589 57464
rect 77650 57360 77680 57402
rect 77590 57230 77680 57360
rect 78650 57402 78658 57560
rect 78650 57360 78680 57402
rect 78720 57360 78740 57600
rect 78650 57230 78740 57360
rect 2740 56210 2830 56330
rect 2740 55950 2760 56210
rect 2800 56160 2830 56210
rect 2820 56002 2830 56160
rect 3800 56210 3890 56330
rect 3800 56160 3830 56210
rect 2888 56098 2922 56114
rect 2956 56108 2972 56142
rect 3148 56108 3164 56142
rect 3454 56108 3470 56142
rect 3646 56108 3662 56142
rect 2888 56048 2922 56064
rect 3705 56098 3739 56114
rect 2956 56020 2972 56054
rect 3148 56020 3164 56054
rect 3454 56020 3470 56054
rect 3646 56020 3662 56054
rect 3705 56048 3739 56064
rect 2800 55950 2830 56002
rect 2740 55890 2830 55950
rect 2740 55650 2760 55890
rect 2800 55850 2830 55890
rect 2820 55692 2830 55850
rect 3800 56002 3808 56160
rect 3800 55970 3830 56002
rect 3870 55970 3890 56210
rect 3800 55890 3890 55970
rect 3800 55850 3830 55890
rect 2888 55788 2922 55804
rect 2956 55798 2972 55832
rect 3148 55798 3164 55832
rect 3454 55798 3470 55832
rect 3646 55798 3662 55832
rect 2888 55738 2922 55754
rect 3705 55788 3739 55804
rect 2956 55710 2972 55744
rect 3148 55710 3164 55744
rect 3454 55710 3470 55744
rect 3646 55710 3662 55744
rect 3705 55738 3739 55754
rect 2800 55650 2830 55692
rect 2740 55520 2830 55650
rect 3800 55692 3808 55850
rect 3800 55650 3830 55692
rect 3870 55650 3890 55890
rect 3800 55520 3890 55650
rect 7730 56210 7820 56330
rect 7730 55950 7750 56210
rect 7790 56160 7820 56210
rect 7810 56002 7820 56160
rect 8790 56210 8880 56330
rect 8790 56160 8820 56210
rect 7878 56098 7912 56114
rect 7946 56108 7962 56142
rect 8138 56108 8154 56142
rect 8444 56108 8460 56142
rect 8636 56108 8652 56142
rect 7878 56048 7912 56064
rect 8695 56098 8729 56114
rect 7946 56020 7962 56054
rect 8138 56020 8154 56054
rect 8444 56020 8460 56054
rect 8636 56020 8652 56054
rect 8695 56048 8729 56064
rect 7790 55950 7820 56002
rect 7730 55890 7820 55950
rect 7730 55650 7750 55890
rect 7790 55850 7820 55890
rect 7810 55692 7820 55850
rect 8790 56002 8798 56160
rect 8790 55970 8820 56002
rect 8860 55970 8880 56210
rect 8790 55890 8880 55970
rect 8790 55850 8820 55890
rect 7878 55788 7912 55804
rect 7946 55798 7962 55832
rect 8138 55798 8154 55832
rect 8444 55798 8460 55832
rect 8636 55798 8652 55832
rect 7878 55738 7912 55754
rect 8695 55788 8729 55804
rect 7946 55710 7962 55744
rect 8138 55710 8154 55744
rect 8444 55710 8460 55744
rect 8636 55710 8652 55744
rect 8695 55738 8729 55754
rect 7790 55650 7820 55692
rect 7730 55520 7820 55650
rect 8790 55692 8798 55850
rect 8790 55650 8820 55692
rect 8860 55650 8880 55890
rect 8790 55520 8880 55650
rect 12720 56210 12810 56330
rect 12720 55950 12740 56210
rect 12780 56160 12810 56210
rect 12800 56002 12810 56160
rect 13780 56210 13870 56330
rect 13780 56160 13810 56210
rect 12868 56098 12902 56114
rect 12936 56108 12952 56142
rect 13128 56108 13144 56142
rect 13434 56108 13450 56142
rect 13626 56108 13642 56142
rect 12868 56048 12902 56064
rect 13685 56098 13719 56114
rect 12936 56020 12952 56054
rect 13128 56020 13144 56054
rect 13434 56020 13450 56054
rect 13626 56020 13642 56054
rect 13685 56048 13719 56064
rect 12780 55950 12810 56002
rect 12720 55890 12810 55950
rect 12720 55650 12740 55890
rect 12780 55850 12810 55890
rect 12800 55692 12810 55850
rect 13780 56002 13788 56160
rect 13780 55970 13810 56002
rect 13850 55970 13870 56210
rect 13780 55890 13870 55970
rect 13780 55850 13810 55890
rect 12868 55788 12902 55804
rect 12936 55798 12952 55832
rect 13128 55798 13144 55832
rect 13434 55798 13450 55832
rect 13626 55798 13642 55832
rect 12868 55738 12902 55754
rect 13685 55788 13719 55804
rect 12936 55710 12952 55744
rect 13128 55710 13144 55744
rect 13434 55710 13450 55744
rect 13626 55710 13642 55744
rect 13685 55738 13719 55754
rect 12780 55650 12810 55692
rect 12720 55520 12810 55650
rect 13780 55692 13788 55850
rect 13780 55650 13810 55692
rect 13850 55650 13870 55890
rect 13780 55520 13870 55650
rect 17710 56210 17800 56330
rect 17710 55950 17730 56210
rect 17770 56160 17800 56210
rect 17790 56002 17800 56160
rect 18770 56210 18860 56330
rect 18770 56160 18800 56210
rect 17858 56098 17892 56114
rect 17926 56108 17942 56142
rect 18118 56108 18134 56142
rect 18424 56108 18440 56142
rect 18616 56108 18632 56142
rect 17858 56048 17892 56064
rect 18675 56098 18709 56114
rect 17926 56020 17942 56054
rect 18118 56020 18134 56054
rect 18424 56020 18440 56054
rect 18616 56020 18632 56054
rect 18675 56048 18709 56064
rect 17770 55950 17800 56002
rect 17710 55890 17800 55950
rect 17710 55650 17730 55890
rect 17770 55850 17800 55890
rect 17790 55692 17800 55850
rect 18770 56002 18778 56160
rect 18770 55970 18800 56002
rect 18840 55970 18860 56210
rect 18770 55890 18860 55970
rect 18770 55850 18800 55890
rect 17858 55788 17892 55804
rect 17926 55798 17942 55832
rect 18118 55798 18134 55832
rect 18424 55798 18440 55832
rect 18616 55798 18632 55832
rect 17858 55738 17892 55754
rect 18675 55788 18709 55804
rect 17926 55710 17942 55744
rect 18118 55710 18134 55744
rect 18424 55710 18440 55744
rect 18616 55710 18632 55744
rect 18675 55738 18709 55754
rect 17770 55650 17800 55692
rect 17710 55520 17800 55650
rect 18770 55692 18778 55850
rect 18770 55650 18800 55692
rect 18840 55650 18860 55890
rect 18770 55520 18860 55650
rect 22700 56210 22790 56330
rect 22700 55950 22720 56210
rect 22760 56160 22790 56210
rect 22780 56002 22790 56160
rect 23760 56210 23850 56330
rect 23760 56160 23790 56210
rect 22848 56098 22882 56114
rect 22916 56108 22932 56142
rect 23108 56108 23124 56142
rect 23414 56108 23430 56142
rect 23606 56108 23622 56142
rect 22848 56048 22882 56064
rect 23665 56098 23699 56114
rect 22916 56020 22932 56054
rect 23108 56020 23124 56054
rect 23414 56020 23430 56054
rect 23606 56020 23622 56054
rect 23665 56048 23699 56064
rect 22760 55950 22790 56002
rect 22700 55890 22790 55950
rect 22700 55650 22720 55890
rect 22760 55850 22790 55890
rect 22780 55692 22790 55850
rect 23760 56002 23768 56160
rect 23760 55970 23790 56002
rect 23830 55970 23850 56210
rect 23760 55890 23850 55970
rect 23760 55850 23790 55890
rect 22848 55788 22882 55804
rect 22916 55798 22932 55832
rect 23108 55798 23124 55832
rect 23414 55798 23430 55832
rect 23606 55798 23622 55832
rect 22848 55738 22882 55754
rect 23665 55788 23699 55804
rect 22916 55710 22932 55744
rect 23108 55710 23124 55744
rect 23414 55710 23430 55744
rect 23606 55710 23622 55744
rect 23665 55738 23699 55754
rect 22760 55650 22790 55692
rect 22700 55520 22790 55650
rect 23760 55692 23768 55850
rect 23760 55650 23790 55692
rect 23830 55650 23850 55890
rect 23760 55520 23850 55650
rect 27690 56210 27780 56330
rect 27690 55950 27710 56210
rect 27750 56160 27780 56210
rect 27770 56002 27780 56160
rect 28750 56210 28840 56330
rect 28750 56160 28780 56210
rect 27838 56098 27872 56114
rect 27906 56108 27922 56142
rect 28098 56108 28114 56142
rect 28404 56108 28420 56142
rect 28596 56108 28612 56142
rect 27838 56048 27872 56064
rect 28655 56098 28689 56114
rect 27906 56020 27922 56054
rect 28098 56020 28114 56054
rect 28404 56020 28420 56054
rect 28596 56020 28612 56054
rect 28655 56048 28689 56064
rect 27750 55950 27780 56002
rect 27690 55890 27780 55950
rect 27690 55650 27710 55890
rect 27750 55850 27780 55890
rect 27770 55692 27780 55850
rect 28750 56002 28758 56160
rect 28750 55970 28780 56002
rect 28820 55970 28840 56210
rect 28750 55890 28840 55970
rect 28750 55850 28780 55890
rect 27838 55788 27872 55804
rect 27906 55798 27922 55832
rect 28098 55798 28114 55832
rect 28404 55798 28420 55832
rect 28596 55798 28612 55832
rect 27838 55738 27872 55754
rect 28655 55788 28689 55804
rect 27906 55710 27922 55744
rect 28098 55710 28114 55744
rect 28404 55710 28420 55744
rect 28596 55710 28612 55744
rect 28655 55738 28689 55754
rect 27750 55650 27780 55692
rect 27690 55520 27780 55650
rect 28750 55692 28758 55850
rect 28750 55650 28780 55692
rect 28820 55650 28840 55890
rect 28750 55520 28840 55650
rect 32680 56210 32770 56330
rect 32680 55950 32700 56210
rect 32740 56160 32770 56210
rect 32760 56002 32770 56160
rect 33740 56210 33830 56330
rect 33740 56160 33770 56210
rect 32828 56098 32862 56114
rect 32896 56108 32912 56142
rect 33088 56108 33104 56142
rect 33394 56108 33410 56142
rect 33586 56108 33602 56142
rect 32828 56048 32862 56064
rect 33645 56098 33679 56114
rect 32896 56020 32912 56054
rect 33088 56020 33104 56054
rect 33394 56020 33410 56054
rect 33586 56020 33602 56054
rect 33645 56048 33679 56064
rect 32740 55950 32770 56002
rect 32680 55890 32770 55950
rect 32680 55650 32700 55890
rect 32740 55850 32770 55890
rect 32760 55692 32770 55850
rect 33740 56002 33748 56160
rect 33740 55970 33770 56002
rect 33810 55970 33830 56210
rect 33740 55890 33830 55970
rect 33740 55850 33770 55890
rect 32828 55788 32862 55804
rect 32896 55798 32912 55832
rect 33088 55798 33104 55832
rect 33394 55798 33410 55832
rect 33586 55798 33602 55832
rect 32828 55738 32862 55754
rect 33645 55788 33679 55804
rect 32896 55710 32912 55744
rect 33088 55710 33104 55744
rect 33394 55710 33410 55744
rect 33586 55710 33602 55744
rect 33645 55738 33679 55754
rect 32740 55650 32770 55692
rect 32680 55520 32770 55650
rect 33740 55692 33748 55850
rect 33740 55650 33770 55692
rect 33810 55650 33830 55890
rect 33740 55520 33830 55650
rect 37670 56210 37760 56330
rect 37670 55950 37690 56210
rect 37730 56160 37760 56210
rect 37750 56002 37760 56160
rect 38730 56210 38820 56330
rect 38730 56160 38760 56210
rect 37818 56098 37852 56114
rect 37886 56108 37902 56142
rect 38078 56108 38094 56142
rect 38384 56108 38400 56142
rect 38576 56108 38592 56142
rect 37818 56048 37852 56064
rect 38635 56098 38669 56114
rect 37886 56020 37902 56054
rect 38078 56020 38094 56054
rect 38384 56020 38400 56054
rect 38576 56020 38592 56054
rect 38635 56048 38669 56064
rect 37730 55950 37760 56002
rect 37670 55890 37760 55950
rect 37670 55650 37690 55890
rect 37730 55850 37760 55890
rect 37750 55692 37760 55850
rect 38730 56002 38738 56160
rect 38730 55970 38760 56002
rect 38800 55970 38820 56210
rect 38730 55890 38820 55970
rect 38730 55850 38760 55890
rect 37818 55788 37852 55804
rect 37886 55798 37902 55832
rect 38078 55798 38094 55832
rect 38384 55798 38400 55832
rect 38576 55798 38592 55832
rect 37818 55738 37852 55754
rect 38635 55788 38669 55804
rect 37886 55710 37902 55744
rect 38078 55710 38094 55744
rect 38384 55710 38400 55744
rect 38576 55710 38592 55744
rect 38635 55738 38669 55754
rect 37730 55650 37760 55692
rect 37670 55520 37760 55650
rect 38730 55692 38738 55850
rect 38730 55650 38760 55692
rect 38800 55650 38820 55890
rect 38730 55520 38820 55650
rect 42660 56210 42750 56330
rect 42660 55950 42680 56210
rect 42720 56160 42750 56210
rect 42740 56002 42750 56160
rect 43720 56210 43810 56330
rect 43720 56160 43750 56210
rect 42808 56098 42842 56114
rect 42876 56108 42892 56142
rect 43068 56108 43084 56142
rect 43374 56108 43390 56142
rect 43566 56108 43582 56142
rect 42808 56048 42842 56064
rect 43625 56098 43659 56114
rect 42876 56020 42892 56054
rect 43068 56020 43084 56054
rect 43374 56020 43390 56054
rect 43566 56020 43582 56054
rect 43625 56048 43659 56064
rect 42720 55950 42750 56002
rect 42660 55890 42750 55950
rect 42660 55650 42680 55890
rect 42720 55850 42750 55890
rect 42740 55692 42750 55850
rect 43720 56002 43728 56160
rect 43720 55970 43750 56002
rect 43790 55970 43810 56210
rect 43720 55890 43810 55970
rect 43720 55850 43750 55890
rect 42808 55788 42842 55804
rect 42876 55798 42892 55832
rect 43068 55798 43084 55832
rect 43374 55798 43390 55832
rect 43566 55798 43582 55832
rect 42808 55738 42842 55754
rect 43625 55788 43659 55804
rect 42876 55710 42892 55744
rect 43068 55710 43084 55744
rect 43374 55710 43390 55744
rect 43566 55710 43582 55744
rect 43625 55738 43659 55754
rect 42720 55650 42750 55692
rect 42660 55520 42750 55650
rect 43720 55692 43728 55850
rect 43720 55650 43750 55692
rect 43790 55650 43810 55890
rect 43720 55520 43810 55650
rect 47650 56210 47740 56330
rect 47650 55950 47670 56210
rect 47710 56160 47740 56210
rect 47730 56002 47740 56160
rect 48710 56210 48800 56330
rect 48710 56160 48740 56210
rect 47798 56098 47832 56114
rect 47866 56108 47882 56142
rect 48058 56108 48074 56142
rect 48364 56108 48380 56142
rect 48556 56108 48572 56142
rect 47798 56048 47832 56064
rect 48615 56098 48649 56114
rect 47866 56020 47882 56054
rect 48058 56020 48074 56054
rect 48364 56020 48380 56054
rect 48556 56020 48572 56054
rect 48615 56048 48649 56064
rect 47710 55950 47740 56002
rect 47650 55890 47740 55950
rect 47650 55650 47670 55890
rect 47710 55850 47740 55890
rect 47730 55692 47740 55850
rect 48710 56002 48718 56160
rect 48710 55970 48740 56002
rect 48780 55970 48800 56210
rect 48710 55890 48800 55970
rect 48710 55850 48740 55890
rect 47798 55788 47832 55804
rect 47866 55798 47882 55832
rect 48058 55798 48074 55832
rect 48364 55798 48380 55832
rect 48556 55798 48572 55832
rect 47798 55738 47832 55754
rect 48615 55788 48649 55804
rect 47866 55710 47882 55744
rect 48058 55710 48074 55744
rect 48364 55710 48380 55744
rect 48556 55710 48572 55744
rect 48615 55738 48649 55754
rect 47710 55650 47740 55692
rect 47650 55520 47740 55650
rect 48710 55692 48718 55850
rect 48710 55650 48740 55692
rect 48780 55650 48800 55890
rect 48710 55520 48800 55650
rect 52640 56210 52730 56330
rect 52640 55950 52660 56210
rect 52700 56160 52730 56210
rect 52720 56002 52730 56160
rect 53700 56210 53790 56330
rect 53700 56160 53730 56210
rect 52788 56098 52822 56114
rect 52856 56108 52872 56142
rect 53048 56108 53064 56142
rect 53354 56108 53370 56142
rect 53546 56108 53562 56142
rect 52788 56048 52822 56064
rect 53605 56098 53639 56114
rect 52856 56020 52872 56054
rect 53048 56020 53064 56054
rect 53354 56020 53370 56054
rect 53546 56020 53562 56054
rect 53605 56048 53639 56064
rect 52700 55950 52730 56002
rect 52640 55890 52730 55950
rect 52640 55650 52660 55890
rect 52700 55850 52730 55890
rect 52720 55692 52730 55850
rect 53700 56002 53708 56160
rect 53700 55970 53730 56002
rect 53770 55970 53790 56210
rect 53700 55890 53790 55970
rect 53700 55850 53730 55890
rect 52788 55788 52822 55804
rect 52856 55798 52872 55832
rect 53048 55798 53064 55832
rect 53354 55798 53370 55832
rect 53546 55798 53562 55832
rect 52788 55738 52822 55754
rect 53605 55788 53639 55804
rect 52856 55710 52872 55744
rect 53048 55710 53064 55744
rect 53354 55710 53370 55744
rect 53546 55710 53562 55744
rect 53605 55738 53639 55754
rect 52700 55650 52730 55692
rect 52640 55520 52730 55650
rect 53700 55692 53708 55850
rect 53700 55650 53730 55692
rect 53770 55650 53790 55890
rect 53700 55520 53790 55650
rect 57630 56210 57720 56330
rect 57630 55950 57650 56210
rect 57690 56160 57720 56210
rect 57710 56002 57720 56160
rect 58690 56210 58780 56330
rect 58690 56160 58720 56210
rect 57778 56098 57812 56114
rect 57846 56108 57862 56142
rect 58038 56108 58054 56142
rect 58344 56108 58360 56142
rect 58536 56108 58552 56142
rect 57778 56048 57812 56064
rect 58595 56098 58629 56114
rect 57846 56020 57862 56054
rect 58038 56020 58054 56054
rect 58344 56020 58360 56054
rect 58536 56020 58552 56054
rect 58595 56048 58629 56064
rect 57690 55950 57720 56002
rect 57630 55890 57720 55950
rect 57630 55650 57650 55890
rect 57690 55850 57720 55890
rect 57710 55692 57720 55850
rect 58690 56002 58698 56160
rect 58690 55970 58720 56002
rect 58760 55970 58780 56210
rect 58690 55890 58780 55970
rect 58690 55850 58720 55890
rect 57778 55788 57812 55804
rect 57846 55798 57862 55832
rect 58038 55798 58054 55832
rect 58344 55798 58360 55832
rect 58536 55798 58552 55832
rect 57778 55738 57812 55754
rect 58595 55788 58629 55804
rect 57846 55710 57862 55744
rect 58038 55710 58054 55744
rect 58344 55710 58360 55744
rect 58536 55710 58552 55744
rect 58595 55738 58629 55754
rect 57690 55650 57720 55692
rect 57630 55520 57720 55650
rect 58690 55692 58698 55850
rect 58690 55650 58720 55692
rect 58760 55650 58780 55890
rect 58690 55520 58780 55650
rect 62620 56210 62710 56330
rect 62620 55950 62640 56210
rect 62680 56160 62710 56210
rect 62700 56002 62710 56160
rect 63680 56210 63770 56330
rect 63680 56160 63710 56210
rect 62768 56098 62802 56114
rect 62836 56108 62852 56142
rect 63028 56108 63044 56142
rect 63334 56108 63350 56142
rect 63526 56108 63542 56142
rect 62768 56048 62802 56064
rect 63585 56098 63619 56114
rect 62836 56020 62852 56054
rect 63028 56020 63044 56054
rect 63334 56020 63350 56054
rect 63526 56020 63542 56054
rect 63585 56048 63619 56064
rect 62680 55950 62710 56002
rect 62620 55890 62710 55950
rect 62620 55650 62640 55890
rect 62680 55850 62710 55890
rect 62700 55692 62710 55850
rect 63680 56002 63688 56160
rect 63680 55970 63710 56002
rect 63750 55970 63770 56210
rect 63680 55890 63770 55970
rect 63680 55850 63710 55890
rect 62768 55788 62802 55804
rect 62836 55798 62852 55832
rect 63028 55798 63044 55832
rect 63334 55798 63350 55832
rect 63526 55798 63542 55832
rect 62768 55738 62802 55754
rect 63585 55788 63619 55804
rect 62836 55710 62852 55744
rect 63028 55710 63044 55744
rect 63334 55710 63350 55744
rect 63526 55710 63542 55744
rect 63585 55738 63619 55754
rect 62680 55650 62710 55692
rect 62620 55520 62710 55650
rect 63680 55692 63688 55850
rect 63680 55650 63710 55692
rect 63750 55650 63770 55890
rect 63680 55520 63770 55650
rect 67610 56210 67700 56330
rect 67610 55950 67630 56210
rect 67670 56160 67700 56210
rect 67690 56002 67700 56160
rect 68670 56210 68760 56330
rect 68670 56160 68700 56210
rect 67758 56098 67792 56114
rect 67826 56108 67842 56142
rect 68018 56108 68034 56142
rect 68324 56108 68340 56142
rect 68516 56108 68532 56142
rect 67758 56048 67792 56064
rect 68575 56098 68609 56114
rect 67826 56020 67842 56054
rect 68018 56020 68034 56054
rect 68324 56020 68340 56054
rect 68516 56020 68532 56054
rect 68575 56048 68609 56064
rect 67670 55950 67700 56002
rect 67610 55890 67700 55950
rect 67610 55650 67630 55890
rect 67670 55850 67700 55890
rect 67690 55692 67700 55850
rect 68670 56002 68678 56160
rect 68670 55970 68700 56002
rect 68740 55970 68760 56210
rect 68670 55890 68760 55970
rect 68670 55850 68700 55890
rect 67758 55788 67792 55804
rect 67826 55798 67842 55832
rect 68018 55798 68034 55832
rect 68324 55798 68340 55832
rect 68516 55798 68532 55832
rect 67758 55738 67792 55754
rect 68575 55788 68609 55804
rect 67826 55710 67842 55744
rect 68018 55710 68034 55744
rect 68324 55710 68340 55744
rect 68516 55710 68532 55744
rect 68575 55738 68609 55754
rect 67670 55650 67700 55692
rect 67610 55520 67700 55650
rect 68670 55692 68678 55850
rect 68670 55650 68700 55692
rect 68740 55650 68760 55890
rect 68670 55520 68760 55650
rect 72600 56210 72690 56330
rect 72600 55950 72620 56210
rect 72660 56160 72690 56210
rect 72680 56002 72690 56160
rect 73660 56210 73750 56330
rect 73660 56160 73690 56210
rect 72748 56098 72782 56114
rect 72816 56108 72832 56142
rect 73008 56108 73024 56142
rect 73314 56108 73330 56142
rect 73506 56108 73522 56142
rect 72748 56048 72782 56064
rect 73565 56098 73599 56114
rect 72816 56020 72832 56054
rect 73008 56020 73024 56054
rect 73314 56020 73330 56054
rect 73506 56020 73522 56054
rect 73565 56048 73599 56064
rect 72660 55950 72690 56002
rect 72600 55890 72690 55950
rect 72600 55650 72620 55890
rect 72660 55850 72690 55890
rect 72680 55692 72690 55850
rect 73660 56002 73668 56160
rect 73660 55970 73690 56002
rect 73730 55970 73750 56210
rect 73660 55890 73750 55970
rect 73660 55850 73690 55890
rect 72748 55788 72782 55804
rect 72816 55798 72832 55832
rect 73008 55798 73024 55832
rect 73314 55798 73330 55832
rect 73506 55798 73522 55832
rect 72748 55738 72782 55754
rect 73565 55788 73599 55804
rect 72816 55710 72832 55744
rect 73008 55710 73024 55744
rect 73314 55710 73330 55744
rect 73506 55710 73522 55744
rect 73565 55738 73599 55754
rect 72660 55650 72690 55692
rect 72600 55520 72690 55650
rect 73660 55692 73668 55850
rect 73660 55650 73690 55692
rect 73730 55650 73750 55890
rect 73660 55520 73750 55650
rect 77590 56210 77680 56330
rect 77590 55950 77610 56210
rect 77650 56160 77680 56210
rect 77670 56002 77680 56160
rect 78650 56210 78740 56330
rect 78650 56160 78680 56210
rect 77738 56098 77772 56114
rect 77806 56108 77822 56142
rect 77998 56108 78014 56142
rect 78304 56108 78320 56142
rect 78496 56108 78512 56142
rect 77738 56048 77772 56064
rect 78555 56098 78589 56114
rect 77806 56020 77822 56054
rect 77998 56020 78014 56054
rect 78304 56020 78320 56054
rect 78496 56020 78512 56054
rect 78555 56048 78589 56064
rect 77650 55950 77680 56002
rect 77590 55890 77680 55950
rect 77590 55650 77610 55890
rect 77650 55850 77680 55890
rect 77670 55692 77680 55850
rect 78650 56002 78658 56160
rect 78650 55970 78680 56002
rect 78720 55970 78740 56210
rect 78650 55890 78740 55970
rect 78650 55850 78680 55890
rect 77738 55788 77772 55804
rect 77806 55798 77822 55832
rect 77998 55798 78014 55832
rect 78304 55798 78320 55832
rect 78496 55798 78512 55832
rect 77738 55738 77772 55754
rect 78555 55788 78589 55804
rect 77806 55710 77822 55744
rect 77998 55710 78014 55744
rect 78304 55710 78320 55744
rect 78496 55710 78512 55744
rect 78555 55738 78589 55754
rect 77650 55650 77680 55692
rect 77590 55520 77680 55650
rect 78650 55692 78658 55850
rect 78650 55650 78680 55692
rect 78720 55650 78740 55890
rect 78650 55520 78740 55650
rect 2740 54500 2830 54620
rect 2740 54240 2760 54500
rect 2800 54450 2830 54500
rect 2820 54292 2830 54450
rect 3800 54500 3890 54620
rect 3800 54450 3830 54500
rect 2888 54388 2922 54404
rect 2956 54398 2972 54432
rect 3148 54398 3164 54432
rect 3454 54398 3470 54432
rect 3646 54398 3662 54432
rect 2888 54338 2922 54354
rect 3705 54388 3739 54404
rect 2956 54310 2972 54344
rect 3148 54310 3164 54344
rect 3454 54310 3470 54344
rect 3646 54310 3662 54344
rect 3705 54338 3739 54354
rect 2800 54240 2830 54292
rect 2740 54180 2830 54240
rect 2740 53940 2760 54180
rect 2800 54140 2830 54180
rect 2820 53982 2830 54140
rect 3800 54292 3808 54450
rect 3800 54260 3830 54292
rect 3870 54260 3890 54500
rect 3800 54180 3890 54260
rect 3800 54140 3830 54180
rect 2888 54078 2922 54094
rect 2956 54088 2972 54122
rect 3148 54088 3164 54122
rect 3454 54088 3470 54122
rect 3646 54088 3662 54122
rect 2888 54028 2922 54044
rect 3705 54078 3739 54094
rect 2956 54000 2972 54034
rect 3148 54000 3164 54034
rect 3454 54000 3470 54034
rect 3646 54000 3662 54034
rect 3705 54028 3739 54044
rect 2800 53940 2830 53982
rect 2740 53810 2830 53940
rect 3800 53982 3808 54140
rect 3800 53940 3830 53982
rect 3870 53940 3890 54180
rect 3800 53810 3890 53940
rect 7730 54500 7820 54620
rect 7730 54240 7750 54500
rect 7790 54450 7820 54500
rect 7810 54292 7820 54450
rect 8790 54500 8880 54620
rect 8790 54450 8820 54500
rect 7878 54388 7912 54404
rect 7946 54398 7962 54432
rect 8138 54398 8154 54432
rect 8444 54398 8460 54432
rect 8636 54398 8652 54432
rect 7878 54338 7912 54354
rect 8695 54388 8729 54404
rect 7946 54310 7962 54344
rect 8138 54310 8154 54344
rect 8444 54310 8460 54344
rect 8636 54310 8652 54344
rect 8695 54338 8729 54354
rect 7790 54240 7820 54292
rect 7730 54180 7820 54240
rect 7730 53940 7750 54180
rect 7790 54140 7820 54180
rect 7810 53982 7820 54140
rect 8790 54292 8798 54450
rect 8790 54260 8820 54292
rect 8860 54260 8880 54500
rect 8790 54180 8880 54260
rect 8790 54140 8820 54180
rect 7878 54078 7912 54094
rect 7946 54088 7962 54122
rect 8138 54088 8154 54122
rect 8444 54088 8460 54122
rect 8636 54088 8652 54122
rect 7878 54028 7912 54044
rect 8695 54078 8729 54094
rect 7946 54000 7962 54034
rect 8138 54000 8154 54034
rect 8444 54000 8460 54034
rect 8636 54000 8652 54034
rect 8695 54028 8729 54044
rect 7790 53940 7820 53982
rect 7730 53810 7820 53940
rect 8790 53982 8798 54140
rect 8790 53940 8820 53982
rect 8860 53940 8880 54180
rect 8790 53810 8880 53940
rect 12720 54500 12810 54620
rect 12720 54240 12740 54500
rect 12780 54450 12810 54500
rect 12800 54292 12810 54450
rect 13780 54500 13870 54620
rect 13780 54450 13810 54500
rect 12868 54388 12902 54404
rect 12936 54398 12952 54432
rect 13128 54398 13144 54432
rect 13434 54398 13450 54432
rect 13626 54398 13642 54432
rect 12868 54338 12902 54354
rect 13685 54388 13719 54404
rect 12936 54310 12952 54344
rect 13128 54310 13144 54344
rect 13434 54310 13450 54344
rect 13626 54310 13642 54344
rect 13685 54338 13719 54354
rect 12780 54240 12810 54292
rect 12720 54180 12810 54240
rect 12720 53940 12740 54180
rect 12780 54140 12810 54180
rect 12800 53982 12810 54140
rect 13780 54292 13788 54450
rect 13780 54260 13810 54292
rect 13850 54260 13870 54500
rect 13780 54180 13870 54260
rect 13780 54140 13810 54180
rect 12868 54078 12902 54094
rect 12936 54088 12952 54122
rect 13128 54088 13144 54122
rect 13434 54088 13450 54122
rect 13626 54088 13642 54122
rect 12868 54028 12902 54044
rect 13685 54078 13719 54094
rect 12936 54000 12952 54034
rect 13128 54000 13144 54034
rect 13434 54000 13450 54034
rect 13626 54000 13642 54034
rect 13685 54028 13719 54044
rect 12780 53940 12810 53982
rect 12720 53810 12810 53940
rect 13780 53982 13788 54140
rect 13780 53940 13810 53982
rect 13850 53940 13870 54180
rect 13780 53810 13870 53940
rect 17710 54500 17800 54620
rect 17710 54240 17730 54500
rect 17770 54450 17800 54500
rect 17790 54292 17800 54450
rect 18770 54500 18860 54620
rect 18770 54450 18800 54500
rect 17858 54388 17892 54404
rect 17926 54398 17942 54432
rect 18118 54398 18134 54432
rect 18424 54398 18440 54432
rect 18616 54398 18632 54432
rect 17858 54338 17892 54354
rect 18675 54388 18709 54404
rect 17926 54310 17942 54344
rect 18118 54310 18134 54344
rect 18424 54310 18440 54344
rect 18616 54310 18632 54344
rect 18675 54338 18709 54354
rect 17770 54240 17800 54292
rect 17710 54180 17800 54240
rect 17710 53940 17730 54180
rect 17770 54140 17800 54180
rect 17790 53982 17800 54140
rect 18770 54292 18778 54450
rect 18770 54260 18800 54292
rect 18840 54260 18860 54500
rect 18770 54180 18860 54260
rect 18770 54140 18800 54180
rect 17858 54078 17892 54094
rect 17926 54088 17942 54122
rect 18118 54088 18134 54122
rect 18424 54088 18440 54122
rect 18616 54088 18632 54122
rect 17858 54028 17892 54044
rect 18675 54078 18709 54094
rect 17926 54000 17942 54034
rect 18118 54000 18134 54034
rect 18424 54000 18440 54034
rect 18616 54000 18632 54034
rect 18675 54028 18709 54044
rect 17770 53940 17800 53982
rect 17710 53810 17800 53940
rect 18770 53982 18778 54140
rect 18770 53940 18800 53982
rect 18840 53940 18860 54180
rect 18770 53810 18860 53940
rect 22700 54500 22790 54620
rect 22700 54240 22720 54500
rect 22760 54450 22790 54500
rect 22780 54292 22790 54450
rect 23760 54500 23850 54620
rect 23760 54450 23790 54500
rect 22848 54388 22882 54404
rect 22916 54398 22932 54432
rect 23108 54398 23124 54432
rect 23414 54398 23430 54432
rect 23606 54398 23622 54432
rect 22848 54338 22882 54354
rect 23665 54388 23699 54404
rect 22916 54310 22932 54344
rect 23108 54310 23124 54344
rect 23414 54310 23430 54344
rect 23606 54310 23622 54344
rect 23665 54338 23699 54354
rect 22760 54240 22790 54292
rect 22700 54180 22790 54240
rect 22700 53940 22720 54180
rect 22760 54140 22790 54180
rect 22780 53982 22790 54140
rect 23760 54292 23768 54450
rect 23760 54260 23790 54292
rect 23830 54260 23850 54500
rect 23760 54180 23850 54260
rect 23760 54140 23790 54180
rect 22848 54078 22882 54094
rect 22916 54088 22932 54122
rect 23108 54088 23124 54122
rect 23414 54088 23430 54122
rect 23606 54088 23622 54122
rect 22848 54028 22882 54044
rect 23665 54078 23699 54094
rect 22916 54000 22932 54034
rect 23108 54000 23124 54034
rect 23414 54000 23430 54034
rect 23606 54000 23622 54034
rect 23665 54028 23699 54044
rect 22760 53940 22790 53982
rect 22700 53810 22790 53940
rect 23760 53982 23768 54140
rect 23760 53940 23790 53982
rect 23830 53940 23850 54180
rect 23760 53810 23850 53940
rect 27690 54500 27780 54620
rect 27690 54240 27710 54500
rect 27750 54450 27780 54500
rect 27770 54292 27780 54450
rect 28750 54500 28840 54620
rect 28750 54450 28780 54500
rect 27838 54388 27872 54404
rect 27906 54398 27922 54432
rect 28098 54398 28114 54432
rect 28404 54398 28420 54432
rect 28596 54398 28612 54432
rect 27838 54338 27872 54354
rect 28655 54388 28689 54404
rect 27906 54310 27922 54344
rect 28098 54310 28114 54344
rect 28404 54310 28420 54344
rect 28596 54310 28612 54344
rect 28655 54338 28689 54354
rect 27750 54240 27780 54292
rect 27690 54180 27780 54240
rect 27690 53940 27710 54180
rect 27750 54140 27780 54180
rect 27770 53982 27780 54140
rect 28750 54292 28758 54450
rect 28750 54260 28780 54292
rect 28820 54260 28840 54500
rect 28750 54180 28840 54260
rect 28750 54140 28780 54180
rect 27838 54078 27872 54094
rect 27906 54088 27922 54122
rect 28098 54088 28114 54122
rect 28404 54088 28420 54122
rect 28596 54088 28612 54122
rect 27838 54028 27872 54044
rect 28655 54078 28689 54094
rect 27906 54000 27922 54034
rect 28098 54000 28114 54034
rect 28404 54000 28420 54034
rect 28596 54000 28612 54034
rect 28655 54028 28689 54044
rect 27750 53940 27780 53982
rect 27690 53810 27780 53940
rect 28750 53982 28758 54140
rect 28750 53940 28780 53982
rect 28820 53940 28840 54180
rect 28750 53810 28840 53940
rect 32680 54500 32770 54620
rect 32680 54240 32700 54500
rect 32740 54450 32770 54500
rect 32760 54292 32770 54450
rect 33740 54500 33830 54620
rect 33740 54450 33770 54500
rect 32828 54388 32862 54404
rect 32896 54398 32912 54432
rect 33088 54398 33104 54432
rect 33394 54398 33410 54432
rect 33586 54398 33602 54432
rect 32828 54338 32862 54354
rect 33645 54388 33679 54404
rect 32896 54310 32912 54344
rect 33088 54310 33104 54344
rect 33394 54310 33410 54344
rect 33586 54310 33602 54344
rect 33645 54338 33679 54354
rect 32740 54240 32770 54292
rect 32680 54180 32770 54240
rect 32680 53940 32700 54180
rect 32740 54140 32770 54180
rect 32760 53982 32770 54140
rect 33740 54292 33748 54450
rect 33740 54260 33770 54292
rect 33810 54260 33830 54500
rect 33740 54180 33830 54260
rect 33740 54140 33770 54180
rect 32828 54078 32862 54094
rect 32896 54088 32912 54122
rect 33088 54088 33104 54122
rect 33394 54088 33410 54122
rect 33586 54088 33602 54122
rect 32828 54028 32862 54044
rect 33645 54078 33679 54094
rect 32896 54000 32912 54034
rect 33088 54000 33104 54034
rect 33394 54000 33410 54034
rect 33586 54000 33602 54034
rect 33645 54028 33679 54044
rect 32740 53940 32770 53982
rect 32680 53810 32770 53940
rect 33740 53982 33748 54140
rect 33740 53940 33770 53982
rect 33810 53940 33830 54180
rect 33740 53810 33830 53940
rect 37670 54500 37760 54620
rect 37670 54240 37690 54500
rect 37730 54450 37760 54500
rect 37750 54292 37760 54450
rect 38730 54500 38820 54620
rect 38730 54450 38760 54500
rect 37818 54388 37852 54404
rect 37886 54398 37902 54432
rect 38078 54398 38094 54432
rect 38384 54398 38400 54432
rect 38576 54398 38592 54432
rect 37818 54338 37852 54354
rect 38635 54388 38669 54404
rect 37886 54310 37902 54344
rect 38078 54310 38094 54344
rect 38384 54310 38400 54344
rect 38576 54310 38592 54344
rect 38635 54338 38669 54354
rect 37730 54240 37760 54292
rect 37670 54180 37760 54240
rect 37670 53940 37690 54180
rect 37730 54140 37760 54180
rect 37750 53982 37760 54140
rect 38730 54292 38738 54450
rect 38730 54260 38760 54292
rect 38800 54260 38820 54500
rect 38730 54180 38820 54260
rect 38730 54140 38760 54180
rect 37818 54078 37852 54094
rect 37886 54088 37902 54122
rect 38078 54088 38094 54122
rect 38384 54088 38400 54122
rect 38576 54088 38592 54122
rect 37818 54028 37852 54044
rect 38635 54078 38669 54094
rect 37886 54000 37902 54034
rect 38078 54000 38094 54034
rect 38384 54000 38400 54034
rect 38576 54000 38592 54034
rect 38635 54028 38669 54044
rect 37730 53940 37760 53982
rect 37670 53810 37760 53940
rect 38730 53982 38738 54140
rect 38730 53940 38760 53982
rect 38800 53940 38820 54180
rect 38730 53810 38820 53940
rect 42660 54500 42750 54620
rect 42660 54240 42680 54500
rect 42720 54450 42750 54500
rect 42740 54292 42750 54450
rect 43720 54500 43810 54620
rect 43720 54450 43750 54500
rect 42808 54388 42842 54404
rect 42876 54398 42892 54432
rect 43068 54398 43084 54432
rect 43374 54398 43390 54432
rect 43566 54398 43582 54432
rect 42808 54338 42842 54354
rect 43625 54388 43659 54404
rect 42876 54310 42892 54344
rect 43068 54310 43084 54344
rect 43374 54310 43390 54344
rect 43566 54310 43582 54344
rect 43625 54338 43659 54354
rect 42720 54240 42750 54292
rect 42660 54180 42750 54240
rect 42660 53940 42680 54180
rect 42720 54140 42750 54180
rect 42740 53982 42750 54140
rect 43720 54292 43728 54450
rect 43720 54260 43750 54292
rect 43790 54260 43810 54500
rect 43720 54180 43810 54260
rect 43720 54140 43750 54180
rect 42808 54078 42842 54094
rect 42876 54088 42892 54122
rect 43068 54088 43084 54122
rect 43374 54088 43390 54122
rect 43566 54088 43582 54122
rect 42808 54028 42842 54044
rect 43625 54078 43659 54094
rect 42876 54000 42892 54034
rect 43068 54000 43084 54034
rect 43374 54000 43390 54034
rect 43566 54000 43582 54034
rect 43625 54028 43659 54044
rect 42720 53940 42750 53982
rect 42660 53810 42750 53940
rect 43720 53982 43728 54140
rect 43720 53940 43750 53982
rect 43790 53940 43810 54180
rect 43720 53810 43810 53940
rect 47650 54500 47740 54620
rect 47650 54240 47670 54500
rect 47710 54450 47740 54500
rect 47730 54292 47740 54450
rect 48710 54500 48800 54620
rect 48710 54450 48740 54500
rect 47798 54388 47832 54404
rect 47866 54398 47882 54432
rect 48058 54398 48074 54432
rect 48364 54398 48380 54432
rect 48556 54398 48572 54432
rect 47798 54338 47832 54354
rect 48615 54388 48649 54404
rect 47866 54310 47882 54344
rect 48058 54310 48074 54344
rect 48364 54310 48380 54344
rect 48556 54310 48572 54344
rect 48615 54338 48649 54354
rect 47710 54240 47740 54292
rect 47650 54180 47740 54240
rect 47650 53940 47670 54180
rect 47710 54140 47740 54180
rect 47730 53982 47740 54140
rect 48710 54292 48718 54450
rect 48710 54260 48740 54292
rect 48780 54260 48800 54500
rect 48710 54180 48800 54260
rect 48710 54140 48740 54180
rect 47798 54078 47832 54094
rect 47866 54088 47882 54122
rect 48058 54088 48074 54122
rect 48364 54088 48380 54122
rect 48556 54088 48572 54122
rect 47798 54028 47832 54044
rect 48615 54078 48649 54094
rect 47866 54000 47882 54034
rect 48058 54000 48074 54034
rect 48364 54000 48380 54034
rect 48556 54000 48572 54034
rect 48615 54028 48649 54044
rect 47710 53940 47740 53982
rect 47650 53810 47740 53940
rect 48710 53982 48718 54140
rect 48710 53940 48740 53982
rect 48780 53940 48800 54180
rect 48710 53810 48800 53940
rect 52640 54500 52730 54620
rect 52640 54240 52660 54500
rect 52700 54450 52730 54500
rect 52720 54292 52730 54450
rect 53700 54500 53790 54620
rect 53700 54450 53730 54500
rect 52788 54388 52822 54404
rect 52856 54398 52872 54432
rect 53048 54398 53064 54432
rect 53354 54398 53370 54432
rect 53546 54398 53562 54432
rect 52788 54338 52822 54354
rect 53605 54388 53639 54404
rect 52856 54310 52872 54344
rect 53048 54310 53064 54344
rect 53354 54310 53370 54344
rect 53546 54310 53562 54344
rect 53605 54338 53639 54354
rect 52700 54240 52730 54292
rect 52640 54180 52730 54240
rect 52640 53940 52660 54180
rect 52700 54140 52730 54180
rect 52720 53982 52730 54140
rect 53700 54292 53708 54450
rect 53700 54260 53730 54292
rect 53770 54260 53790 54500
rect 53700 54180 53790 54260
rect 53700 54140 53730 54180
rect 52788 54078 52822 54094
rect 52856 54088 52872 54122
rect 53048 54088 53064 54122
rect 53354 54088 53370 54122
rect 53546 54088 53562 54122
rect 52788 54028 52822 54044
rect 53605 54078 53639 54094
rect 52856 54000 52872 54034
rect 53048 54000 53064 54034
rect 53354 54000 53370 54034
rect 53546 54000 53562 54034
rect 53605 54028 53639 54044
rect 52700 53940 52730 53982
rect 52640 53810 52730 53940
rect 53700 53982 53708 54140
rect 53700 53940 53730 53982
rect 53770 53940 53790 54180
rect 53700 53810 53790 53940
rect 57630 54500 57720 54620
rect 57630 54240 57650 54500
rect 57690 54450 57720 54500
rect 57710 54292 57720 54450
rect 58690 54500 58780 54620
rect 58690 54450 58720 54500
rect 57778 54388 57812 54404
rect 57846 54398 57862 54432
rect 58038 54398 58054 54432
rect 58344 54398 58360 54432
rect 58536 54398 58552 54432
rect 57778 54338 57812 54354
rect 58595 54388 58629 54404
rect 57846 54310 57862 54344
rect 58038 54310 58054 54344
rect 58344 54310 58360 54344
rect 58536 54310 58552 54344
rect 58595 54338 58629 54354
rect 57690 54240 57720 54292
rect 57630 54180 57720 54240
rect 57630 53940 57650 54180
rect 57690 54140 57720 54180
rect 57710 53982 57720 54140
rect 58690 54292 58698 54450
rect 58690 54260 58720 54292
rect 58760 54260 58780 54500
rect 58690 54180 58780 54260
rect 58690 54140 58720 54180
rect 57778 54078 57812 54094
rect 57846 54088 57862 54122
rect 58038 54088 58054 54122
rect 58344 54088 58360 54122
rect 58536 54088 58552 54122
rect 57778 54028 57812 54044
rect 58595 54078 58629 54094
rect 57846 54000 57862 54034
rect 58038 54000 58054 54034
rect 58344 54000 58360 54034
rect 58536 54000 58552 54034
rect 58595 54028 58629 54044
rect 57690 53940 57720 53982
rect 57630 53810 57720 53940
rect 58690 53982 58698 54140
rect 58690 53940 58720 53982
rect 58760 53940 58780 54180
rect 58690 53810 58780 53940
rect 62620 54500 62710 54620
rect 62620 54240 62640 54500
rect 62680 54450 62710 54500
rect 62700 54292 62710 54450
rect 63680 54500 63770 54620
rect 63680 54450 63710 54500
rect 62768 54388 62802 54404
rect 62836 54398 62852 54432
rect 63028 54398 63044 54432
rect 63334 54398 63350 54432
rect 63526 54398 63542 54432
rect 62768 54338 62802 54354
rect 63585 54388 63619 54404
rect 62836 54310 62852 54344
rect 63028 54310 63044 54344
rect 63334 54310 63350 54344
rect 63526 54310 63542 54344
rect 63585 54338 63619 54354
rect 62680 54240 62710 54292
rect 62620 54180 62710 54240
rect 62620 53940 62640 54180
rect 62680 54140 62710 54180
rect 62700 53982 62710 54140
rect 63680 54292 63688 54450
rect 63680 54260 63710 54292
rect 63750 54260 63770 54500
rect 63680 54180 63770 54260
rect 63680 54140 63710 54180
rect 62768 54078 62802 54094
rect 62836 54088 62852 54122
rect 63028 54088 63044 54122
rect 63334 54088 63350 54122
rect 63526 54088 63542 54122
rect 62768 54028 62802 54044
rect 63585 54078 63619 54094
rect 62836 54000 62852 54034
rect 63028 54000 63044 54034
rect 63334 54000 63350 54034
rect 63526 54000 63542 54034
rect 63585 54028 63619 54044
rect 62680 53940 62710 53982
rect 62620 53810 62710 53940
rect 63680 53982 63688 54140
rect 63680 53940 63710 53982
rect 63750 53940 63770 54180
rect 63680 53810 63770 53940
rect 67610 54500 67700 54620
rect 67610 54240 67630 54500
rect 67670 54450 67700 54500
rect 67690 54292 67700 54450
rect 68670 54500 68760 54620
rect 68670 54450 68700 54500
rect 67758 54388 67792 54404
rect 67826 54398 67842 54432
rect 68018 54398 68034 54432
rect 68324 54398 68340 54432
rect 68516 54398 68532 54432
rect 67758 54338 67792 54354
rect 68575 54388 68609 54404
rect 67826 54310 67842 54344
rect 68018 54310 68034 54344
rect 68324 54310 68340 54344
rect 68516 54310 68532 54344
rect 68575 54338 68609 54354
rect 67670 54240 67700 54292
rect 67610 54180 67700 54240
rect 67610 53940 67630 54180
rect 67670 54140 67700 54180
rect 67690 53982 67700 54140
rect 68670 54292 68678 54450
rect 68670 54260 68700 54292
rect 68740 54260 68760 54500
rect 68670 54180 68760 54260
rect 68670 54140 68700 54180
rect 67758 54078 67792 54094
rect 67826 54088 67842 54122
rect 68018 54088 68034 54122
rect 68324 54088 68340 54122
rect 68516 54088 68532 54122
rect 67758 54028 67792 54044
rect 68575 54078 68609 54094
rect 67826 54000 67842 54034
rect 68018 54000 68034 54034
rect 68324 54000 68340 54034
rect 68516 54000 68532 54034
rect 68575 54028 68609 54044
rect 67670 53940 67700 53982
rect 67610 53810 67700 53940
rect 68670 53982 68678 54140
rect 68670 53940 68700 53982
rect 68740 53940 68760 54180
rect 68670 53810 68760 53940
rect 72600 54500 72690 54620
rect 72600 54240 72620 54500
rect 72660 54450 72690 54500
rect 72680 54292 72690 54450
rect 73660 54500 73750 54620
rect 73660 54450 73690 54500
rect 72748 54388 72782 54404
rect 72816 54398 72832 54432
rect 73008 54398 73024 54432
rect 73314 54398 73330 54432
rect 73506 54398 73522 54432
rect 72748 54338 72782 54354
rect 73565 54388 73599 54404
rect 72816 54310 72832 54344
rect 73008 54310 73024 54344
rect 73314 54310 73330 54344
rect 73506 54310 73522 54344
rect 73565 54338 73599 54354
rect 72660 54240 72690 54292
rect 72600 54180 72690 54240
rect 72600 53940 72620 54180
rect 72660 54140 72690 54180
rect 72680 53982 72690 54140
rect 73660 54292 73668 54450
rect 73660 54260 73690 54292
rect 73730 54260 73750 54500
rect 73660 54180 73750 54260
rect 73660 54140 73690 54180
rect 72748 54078 72782 54094
rect 72816 54088 72832 54122
rect 73008 54088 73024 54122
rect 73314 54088 73330 54122
rect 73506 54088 73522 54122
rect 72748 54028 72782 54044
rect 73565 54078 73599 54094
rect 72816 54000 72832 54034
rect 73008 54000 73024 54034
rect 73314 54000 73330 54034
rect 73506 54000 73522 54034
rect 73565 54028 73599 54044
rect 72660 53940 72690 53982
rect 72600 53810 72690 53940
rect 73660 53982 73668 54140
rect 73660 53940 73690 53982
rect 73730 53940 73750 54180
rect 73660 53810 73750 53940
rect 77590 54500 77680 54620
rect 77590 54240 77610 54500
rect 77650 54450 77680 54500
rect 77670 54292 77680 54450
rect 78650 54500 78740 54620
rect 78650 54450 78680 54500
rect 77738 54388 77772 54404
rect 77806 54398 77822 54432
rect 77998 54398 78014 54432
rect 78304 54398 78320 54432
rect 78496 54398 78512 54432
rect 77738 54338 77772 54354
rect 78555 54388 78589 54404
rect 77806 54310 77822 54344
rect 77998 54310 78014 54344
rect 78304 54310 78320 54344
rect 78496 54310 78512 54344
rect 78555 54338 78589 54354
rect 77650 54240 77680 54292
rect 77590 54180 77680 54240
rect 77590 53940 77610 54180
rect 77650 54140 77680 54180
rect 77670 53982 77680 54140
rect 78650 54292 78658 54450
rect 78650 54260 78680 54292
rect 78720 54260 78740 54500
rect 78650 54180 78740 54260
rect 78650 54140 78680 54180
rect 77738 54078 77772 54094
rect 77806 54088 77822 54122
rect 77998 54088 78014 54122
rect 78304 54088 78320 54122
rect 78496 54088 78512 54122
rect 77738 54028 77772 54044
rect 78555 54078 78589 54094
rect 77806 54000 77822 54034
rect 77998 54000 78014 54034
rect 78304 54000 78320 54034
rect 78496 54000 78512 54034
rect 78555 54028 78589 54044
rect 77650 53940 77680 53982
rect 77590 53810 77680 53940
rect 78650 53982 78658 54140
rect 78650 53940 78680 53982
rect 78720 53940 78740 54180
rect 78650 53810 78740 53940
rect 2740 52790 2830 52910
rect 2740 52530 2760 52790
rect 2800 52740 2830 52790
rect 2820 52582 2830 52740
rect 3800 52790 3890 52910
rect 3800 52740 3830 52790
rect 2888 52678 2922 52694
rect 2956 52688 2972 52722
rect 3148 52688 3164 52722
rect 3454 52688 3470 52722
rect 3646 52688 3662 52722
rect 2888 52628 2922 52644
rect 3705 52678 3739 52694
rect 2956 52600 2972 52634
rect 3148 52600 3164 52634
rect 3454 52600 3470 52634
rect 3646 52600 3662 52634
rect 3705 52628 3739 52644
rect 2800 52530 2830 52582
rect 2740 52470 2830 52530
rect 2740 52230 2760 52470
rect 2800 52430 2830 52470
rect 2820 52272 2830 52430
rect 3800 52582 3808 52740
rect 3800 52550 3830 52582
rect 3870 52550 3890 52790
rect 3800 52470 3890 52550
rect 3800 52430 3830 52470
rect 2888 52368 2922 52384
rect 2956 52378 2972 52412
rect 3148 52378 3164 52412
rect 3454 52378 3470 52412
rect 3646 52378 3662 52412
rect 2888 52318 2922 52334
rect 3705 52368 3739 52384
rect 2956 52290 2972 52324
rect 3148 52290 3164 52324
rect 3454 52290 3470 52324
rect 3646 52290 3662 52324
rect 3705 52318 3739 52334
rect 2800 52230 2830 52272
rect 2740 52100 2830 52230
rect 3800 52272 3808 52430
rect 3800 52230 3830 52272
rect 3870 52230 3890 52470
rect 3800 52100 3890 52230
rect 7730 52790 7820 52910
rect 7730 52530 7750 52790
rect 7790 52740 7820 52790
rect 7810 52582 7820 52740
rect 8790 52790 8880 52910
rect 8790 52740 8820 52790
rect 7878 52678 7912 52694
rect 7946 52688 7962 52722
rect 8138 52688 8154 52722
rect 8444 52688 8460 52722
rect 8636 52688 8652 52722
rect 7878 52628 7912 52644
rect 8695 52678 8729 52694
rect 7946 52600 7962 52634
rect 8138 52600 8154 52634
rect 8444 52600 8460 52634
rect 8636 52600 8652 52634
rect 8695 52628 8729 52644
rect 7790 52530 7820 52582
rect 7730 52470 7820 52530
rect 7730 52230 7750 52470
rect 7790 52430 7820 52470
rect 7810 52272 7820 52430
rect 8790 52582 8798 52740
rect 8790 52550 8820 52582
rect 8860 52550 8880 52790
rect 8790 52470 8880 52550
rect 8790 52430 8820 52470
rect 7878 52368 7912 52384
rect 7946 52378 7962 52412
rect 8138 52378 8154 52412
rect 8444 52378 8460 52412
rect 8636 52378 8652 52412
rect 7878 52318 7912 52334
rect 8695 52368 8729 52384
rect 7946 52290 7962 52324
rect 8138 52290 8154 52324
rect 8444 52290 8460 52324
rect 8636 52290 8652 52324
rect 8695 52318 8729 52334
rect 7790 52230 7820 52272
rect 7730 52100 7820 52230
rect 8790 52272 8798 52430
rect 8790 52230 8820 52272
rect 8860 52230 8880 52470
rect 8790 52100 8880 52230
rect 12720 52790 12810 52910
rect 12720 52530 12740 52790
rect 12780 52740 12810 52790
rect 12800 52582 12810 52740
rect 13780 52790 13870 52910
rect 13780 52740 13810 52790
rect 12868 52678 12902 52694
rect 12936 52688 12952 52722
rect 13128 52688 13144 52722
rect 13434 52688 13450 52722
rect 13626 52688 13642 52722
rect 12868 52628 12902 52644
rect 13685 52678 13719 52694
rect 12936 52600 12952 52634
rect 13128 52600 13144 52634
rect 13434 52600 13450 52634
rect 13626 52600 13642 52634
rect 13685 52628 13719 52644
rect 12780 52530 12810 52582
rect 12720 52470 12810 52530
rect 12720 52230 12740 52470
rect 12780 52430 12810 52470
rect 12800 52272 12810 52430
rect 13780 52582 13788 52740
rect 13780 52550 13810 52582
rect 13850 52550 13870 52790
rect 13780 52470 13870 52550
rect 13780 52430 13810 52470
rect 12868 52368 12902 52384
rect 12936 52378 12952 52412
rect 13128 52378 13144 52412
rect 13434 52378 13450 52412
rect 13626 52378 13642 52412
rect 12868 52318 12902 52334
rect 13685 52368 13719 52384
rect 12936 52290 12952 52324
rect 13128 52290 13144 52324
rect 13434 52290 13450 52324
rect 13626 52290 13642 52324
rect 13685 52318 13719 52334
rect 12780 52230 12810 52272
rect 12720 52100 12810 52230
rect 13780 52272 13788 52430
rect 13780 52230 13810 52272
rect 13850 52230 13870 52470
rect 13780 52100 13870 52230
rect 17710 52790 17800 52910
rect 17710 52530 17730 52790
rect 17770 52740 17800 52790
rect 17790 52582 17800 52740
rect 18770 52790 18860 52910
rect 18770 52740 18800 52790
rect 17858 52678 17892 52694
rect 17926 52688 17942 52722
rect 18118 52688 18134 52722
rect 18424 52688 18440 52722
rect 18616 52688 18632 52722
rect 17858 52628 17892 52644
rect 18675 52678 18709 52694
rect 17926 52600 17942 52634
rect 18118 52600 18134 52634
rect 18424 52600 18440 52634
rect 18616 52600 18632 52634
rect 18675 52628 18709 52644
rect 17770 52530 17800 52582
rect 17710 52470 17800 52530
rect 17710 52230 17730 52470
rect 17770 52430 17800 52470
rect 17790 52272 17800 52430
rect 18770 52582 18778 52740
rect 18770 52550 18800 52582
rect 18840 52550 18860 52790
rect 18770 52470 18860 52550
rect 18770 52430 18800 52470
rect 17858 52368 17892 52384
rect 17926 52378 17942 52412
rect 18118 52378 18134 52412
rect 18424 52378 18440 52412
rect 18616 52378 18632 52412
rect 17858 52318 17892 52334
rect 18675 52368 18709 52384
rect 17926 52290 17942 52324
rect 18118 52290 18134 52324
rect 18424 52290 18440 52324
rect 18616 52290 18632 52324
rect 18675 52318 18709 52334
rect 17770 52230 17800 52272
rect 17710 52100 17800 52230
rect 18770 52272 18778 52430
rect 18770 52230 18800 52272
rect 18840 52230 18860 52470
rect 18770 52100 18860 52230
rect 22700 52790 22790 52910
rect 22700 52530 22720 52790
rect 22760 52740 22790 52790
rect 22780 52582 22790 52740
rect 23760 52790 23850 52910
rect 23760 52740 23790 52790
rect 22848 52678 22882 52694
rect 22916 52688 22932 52722
rect 23108 52688 23124 52722
rect 23414 52688 23430 52722
rect 23606 52688 23622 52722
rect 22848 52628 22882 52644
rect 23665 52678 23699 52694
rect 22916 52600 22932 52634
rect 23108 52600 23124 52634
rect 23414 52600 23430 52634
rect 23606 52600 23622 52634
rect 23665 52628 23699 52644
rect 22760 52530 22790 52582
rect 22700 52470 22790 52530
rect 22700 52230 22720 52470
rect 22760 52430 22790 52470
rect 22780 52272 22790 52430
rect 23760 52582 23768 52740
rect 23760 52550 23790 52582
rect 23830 52550 23850 52790
rect 23760 52470 23850 52550
rect 23760 52430 23790 52470
rect 22848 52368 22882 52384
rect 22916 52378 22932 52412
rect 23108 52378 23124 52412
rect 23414 52378 23430 52412
rect 23606 52378 23622 52412
rect 22848 52318 22882 52334
rect 23665 52368 23699 52384
rect 22916 52290 22932 52324
rect 23108 52290 23124 52324
rect 23414 52290 23430 52324
rect 23606 52290 23622 52324
rect 23665 52318 23699 52334
rect 22760 52230 22790 52272
rect 22700 52100 22790 52230
rect 23760 52272 23768 52430
rect 23760 52230 23790 52272
rect 23830 52230 23850 52470
rect 23760 52100 23850 52230
rect 27690 52790 27780 52910
rect 27690 52530 27710 52790
rect 27750 52740 27780 52790
rect 27770 52582 27780 52740
rect 28750 52790 28840 52910
rect 28750 52740 28780 52790
rect 27838 52678 27872 52694
rect 27906 52688 27922 52722
rect 28098 52688 28114 52722
rect 28404 52688 28420 52722
rect 28596 52688 28612 52722
rect 27838 52628 27872 52644
rect 28655 52678 28689 52694
rect 27906 52600 27922 52634
rect 28098 52600 28114 52634
rect 28404 52600 28420 52634
rect 28596 52600 28612 52634
rect 28655 52628 28689 52644
rect 27750 52530 27780 52582
rect 27690 52470 27780 52530
rect 27690 52230 27710 52470
rect 27750 52430 27780 52470
rect 27770 52272 27780 52430
rect 28750 52582 28758 52740
rect 28750 52550 28780 52582
rect 28820 52550 28840 52790
rect 28750 52470 28840 52550
rect 28750 52430 28780 52470
rect 27838 52368 27872 52384
rect 27906 52378 27922 52412
rect 28098 52378 28114 52412
rect 28404 52378 28420 52412
rect 28596 52378 28612 52412
rect 27838 52318 27872 52334
rect 28655 52368 28689 52384
rect 27906 52290 27922 52324
rect 28098 52290 28114 52324
rect 28404 52290 28420 52324
rect 28596 52290 28612 52324
rect 28655 52318 28689 52334
rect 27750 52230 27780 52272
rect 27690 52100 27780 52230
rect 28750 52272 28758 52430
rect 28750 52230 28780 52272
rect 28820 52230 28840 52470
rect 28750 52100 28840 52230
rect 32680 52790 32770 52910
rect 32680 52530 32700 52790
rect 32740 52740 32770 52790
rect 32760 52582 32770 52740
rect 33740 52790 33830 52910
rect 33740 52740 33770 52790
rect 32828 52678 32862 52694
rect 32896 52688 32912 52722
rect 33088 52688 33104 52722
rect 33394 52688 33410 52722
rect 33586 52688 33602 52722
rect 32828 52628 32862 52644
rect 33645 52678 33679 52694
rect 32896 52600 32912 52634
rect 33088 52600 33104 52634
rect 33394 52600 33410 52634
rect 33586 52600 33602 52634
rect 33645 52628 33679 52644
rect 32740 52530 32770 52582
rect 32680 52470 32770 52530
rect 32680 52230 32700 52470
rect 32740 52430 32770 52470
rect 32760 52272 32770 52430
rect 33740 52582 33748 52740
rect 33740 52550 33770 52582
rect 33810 52550 33830 52790
rect 33740 52470 33830 52550
rect 33740 52430 33770 52470
rect 32828 52368 32862 52384
rect 32896 52378 32912 52412
rect 33088 52378 33104 52412
rect 33394 52378 33410 52412
rect 33586 52378 33602 52412
rect 32828 52318 32862 52334
rect 33645 52368 33679 52384
rect 32896 52290 32912 52324
rect 33088 52290 33104 52324
rect 33394 52290 33410 52324
rect 33586 52290 33602 52324
rect 33645 52318 33679 52334
rect 32740 52230 32770 52272
rect 32680 52100 32770 52230
rect 33740 52272 33748 52430
rect 33740 52230 33770 52272
rect 33810 52230 33830 52470
rect 33740 52100 33830 52230
rect 37670 52790 37760 52910
rect 37670 52530 37690 52790
rect 37730 52740 37760 52790
rect 37750 52582 37760 52740
rect 38730 52790 38820 52910
rect 38730 52740 38760 52790
rect 37818 52678 37852 52694
rect 37886 52688 37902 52722
rect 38078 52688 38094 52722
rect 38384 52688 38400 52722
rect 38576 52688 38592 52722
rect 37818 52628 37852 52644
rect 38635 52678 38669 52694
rect 37886 52600 37902 52634
rect 38078 52600 38094 52634
rect 38384 52600 38400 52634
rect 38576 52600 38592 52634
rect 38635 52628 38669 52644
rect 37730 52530 37760 52582
rect 37670 52470 37760 52530
rect 37670 52230 37690 52470
rect 37730 52430 37760 52470
rect 37750 52272 37760 52430
rect 38730 52582 38738 52740
rect 38730 52550 38760 52582
rect 38800 52550 38820 52790
rect 38730 52470 38820 52550
rect 38730 52430 38760 52470
rect 37818 52368 37852 52384
rect 37886 52378 37902 52412
rect 38078 52378 38094 52412
rect 38384 52378 38400 52412
rect 38576 52378 38592 52412
rect 37818 52318 37852 52334
rect 38635 52368 38669 52384
rect 37886 52290 37902 52324
rect 38078 52290 38094 52324
rect 38384 52290 38400 52324
rect 38576 52290 38592 52324
rect 38635 52318 38669 52334
rect 37730 52230 37760 52272
rect 37670 52100 37760 52230
rect 38730 52272 38738 52430
rect 38730 52230 38760 52272
rect 38800 52230 38820 52470
rect 38730 52100 38820 52230
rect 42660 52790 42750 52910
rect 42660 52530 42680 52790
rect 42720 52740 42750 52790
rect 42740 52582 42750 52740
rect 43720 52790 43810 52910
rect 43720 52740 43750 52790
rect 42808 52678 42842 52694
rect 42876 52688 42892 52722
rect 43068 52688 43084 52722
rect 43374 52688 43390 52722
rect 43566 52688 43582 52722
rect 42808 52628 42842 52644
rect 43625 52678 43659 52694
rect 42876 52600 42892 52634
rect 43068 52600 43084 52634
rect 43374 52600 43390 52634
rect 43566 52600 43582 52634
rect 43625 52628 43659 52644
rect 42720 52530 42750 52582
rect 42660 52470 42750 52530
rect 42660 52230 42680 52470
rect 42720 52430 42750 52470
rect 42740 52272 42750 52430
rect 43720 52582 43728 52740
rect 43720 52550 43750 52582
rect 43790 52550 43810 52790
rect 43720 52470 43810 52550
rect 43720 52430 43750 52470
rect 42808 52368 42842 52384
rect 42876 52378 42892 52412
rect 43068 52378 43084 52412
rect 43374 52378 43390 52412
rect 43566 52378 43582 52412
rect 42808 52318 42842 52334
rect 43625 52368 43659 52384
rect 42876 52290 42892 52324
rect 43068 52290 43084 52324
rect 43374 52290 43390 52324
rect 43566 52290 43582 52324
rect 43625 52318 43659 52334
rect 42720 52230 42750 52272
rect 42660 52100 42750 52230
rect 43720 52272 43728 52430
rect 43720 52230 43750 52272
rect 43790 52230 43810 52470
rect 43720 52100 43810 52230
rect 47650 52790 47740 52910
rect 47650 52530 47670 52790
rect 47710 52740 47740 52790
rect 47730 52582 47740 52740
rect 48710 52790 48800 52910
rect 48710 52740 48740 52790
rect 47798 52678 47832 52694
rect 47866 52688 47882 52722
rect 48058 52688 48074 52722
rect 48364 52688 48380 52722
rect 48556 52688 48572 52722
rect 47798 52628 47832 52644
rect 48615 52678 48649 52694
rect 47866 52600 47882 52634
rect 48058 52600 48074 52634
rect 48364 52600 48380 52634
rect 48556 52600 48572 52634
rect 48615 52628 48649 52644
rect 47710 52530 47740 52582
rect 47650 52470 47740 52530
rect 47650 52230 47670 52470
rect 47710 52430 47740 52470
rect 47730 52272 47740 52430
rect 48710 52582 48718 52740
rect 48710 52550 48740 52582
rect 48780 52550 48800 52790
rect 48710 52470 48800 52550
rect 48710 52430 48740 52470
rect 47798 52368 47832 52384
rect 47866 52378 47882 52412
rect 48058 52378 48074 52412
rect 48364 52378 48380 52412
rect 48556 52378 48572 52412
rect 47798 52318 47832 52334
rect 48615 52368 48649 52384
rect 47866 52290 47882 52324
rect 48058 52290 48074 52324
rect 48364 52290 48380 52324
rect 48556 52290 48572 52324
rect 48615 52318 48649 52334
rect 47710 52230 47740 52272
rect 47650 52100 47740 52230
rect 48710 52272 48718 52430
rect 48710 52230 48740 52272
rect 48780 52230 48800 52470
rect 48710 52100 48800 52230
rect 52640 52790 52730 52910
rect 52640 52530 52660 52790
rect 52700 52740 52730 52790
rect 52720 52582 52730 52740
rect 53700 52790 53790 52910
rect 53700 52740 53730 52790
rect 52788 52678 52822 52694
rect 52856 52688 52872 52722
rect 53048 52688 53064 52722
rect 53354 52688 53370 52722
rect 53546 52688 53562 52722
rect 52788 52628 52822 52644
rect 53605 52678 53639 52694
rect 52856 52600 52872 52634
rect 53048 52600 53064 52634
rect 53354 52600 53370 52634
rect 53546 52600 53562 52634
rect 53605 52628 53639 52644
rect 52700 52530 52730 52582
rect 52640 52470 52730 52530
rect 52640 52230 52660 52470
rect 52700 52430 52730 52470
rect 52720 52272 52730 52430
rect 53700 52582 53708 52740
rect 53700 52550 53730 52582
rect 53770 52550 53790 52790
rect 53700 52470 53790 52550
rect 53700 52430 53730 52470
rect 52788 52368 52822 52384
rect 52856 52378 52872 52412
rect 53048 52378 53064 52412
rect 53354 52378 53370 52412
rect 53546 52378 53562 52412
rect 52788 52318 52822 52334
rect 53605 52368 53639 52384
rect 52856 52290 52872 52324
rect 53048 52290 53064 52324
rect 53354 52290 53370 52324
rect 53546 52290 53562 52324
rect 53605 52318 53639 52334
rect 52700 52230 52730 52272
rect 52640 52100 52730 52230
rect 53700 52272 53708 52430
rect 53700 52230 53730 52272
rect 53770 52230 53790 52470
rect 53700 52100 53790 52230
rect 57630 52790 57720 52910
rect 57630 52530 57650 52790
rect 57690 52740 57720 52790
rect 57710 52582 57720 52740
rect 58690 52790 58780 52910
rect 58690 52740 58720 52790
rect 57778 52678 57812 52694
rect 57846 52688 57862 52722
rect 58038 52688 58054 52722
rect 58344 52688 58360 52722
rect 58536 52688 58552 52722
rect 57778 52628 57812 52644
rect 58595 52678 58629 52694
rect 57846 52600 57862 52634
rect 58038 52600 58054 52634
rect 58344 52600 58360 52634
rect 58536 52600 58552 52634
rect 58595 52628 58629 52644
rect 57690 52530 57720 52582
rect 57630 52470 57720 52530
rect 57630 52230 57650 52470
rect 57690 52430 57720 52470
rect 57710 52272 57720 52430
rect 58690 52582 58698 52740
rect 58690 52550 58720 52582
rect 58760 52550 58780 52790
rect 58690 52470 58780 52550
rect 58690 52430 58720 52470
rect 57778 52368 57812 52384
rect 57846 52378 57862 52412
rect 58038 52378 58054 52412
rect 58344 52378 58360 52412
rect 58536 52378 58552 52412
rect 57778 52318 57812 52334
rect 58595 52368 58629 52384
rect 57846 52290 57862 52324
rect 58038 52290 58054 52324
rect 58344 52290 58360 52324
rect 58536 52290 58552 52324
rect 58595 52318 58629 52334
rect 57690 52230 57720 52272
rect 57630 52100 57720 52230
rect 58690 52272 58698 52430
rect 58690 52230 58720 52272
rect 58760 52230 58780 52470
rect 58690 52100 58780 52230
rect 62620 52790 62710 52910
rect 62620 52530 62640 52790
rect 62680 52740 62710 52790
rect 62700 52582 62710 52740
rect 63680 52790 63770 52910
rect 63680 52740 63710 52790
rect 62768 52678 62802 52694
rect 62836 52688 62852 52722
rect 63028 52688 63044 52722
rect 63334 52688 63350 52722
rect 63526 52688 63542 52722
rect 62768 52628 62802 52644
rect 63585 52678 63619 52694
rect 62836 52600 62852 52634
rect 63028 52600 63044 52634
rect 63334 52600 63350 52634
rect 63526 52600 63542 52634
rect 63585 52628 63619 52644
rect 62680 52530 62710 52582
rect 62620 52470 62710 52530
rect 62620 52230 62640 52470
rect 62680 52430 62710 52470
rect 62700 52272 62710 52430
rect 63680 52582 63688 52740
rect 63680 52550 63710 52582
rect 63750 52550 63770 52790
rect 63680 52470 63770 52550
rect 63680 52430 63710 52470
rect 62768 52368 62802 52384
rect 62836 52378 62852 52412
rect 63028 52378 63044 52412
rect 63334 52378 63350 52412
rect 63526 52378 63542 52412
rect 62768 52318 62802 52334
rect 63585 52368 63619 52384
rect 62836 52290 62852 52324
rect 63028 52290 63044 52324
rect 63334 52290 63350 52324
rect 63526 52290 63542 52324
rect 63585 52318 63619 52334
rect 62680 52230 62710 52272
rect 62620 52100 62710 52230
rect 63680 52272 63688 52430
rect 63680 52230 63710 52272
rect 63750 52230 63770 52470
rect 63680 52100 63770 52230
rect 67610 52790 67700 52910
rect 67610 52530 67630 52790
rect 67670 52740 67700 52790
rect 67690 52582 67700 52740
rect 68670 52790 68760 52910
rect 68670 52740 68700 52790
rect 67758 52678 67792 52694
rect 67826 52688 67842 52722
rect 68018 52688 68034 52722
rect 68324 52688 68340 52722
rect 68516 52688 68532 52722
rect 67758 52628 67792 52644
rect 68575 52678 68609 52694
rect 67826 52600 67842 52634
rect 68018 52600 68034 52634
rect 68324 52600 68340 52634
rect 68516 52600 68532 52634
rect 68575 52628 68609 52644
rect 67670 52530 67700 52582
rect 67610 52470 67700 52530
rect 67610 52230 67630 52470
rect 67670 52430 67700 52470
rect 67690 52272 67700 52430
rect 68670 52582 68678 52740
rect 68670 52550 68700 52582
rect 68740 52550 68760 52790
rect 68670 52470 68760 52550
rect 68670 52430 68700 52470
rect 67758 52368 67792 52384
rect 67826 52378 67842 52412
rect 68018 52378 68034 52412
rect 68324 52378 68340 52412
rect 68516 52378 68532 52412
rect 67758 52318 67792 52334
rect 68575 52368 68609 52384
rect 67826 52290 67842 52324
rect 68018 52290 68034 52324
rect 68324 52290 68340 52324
rect 68516 52290 68532 52324
rect 68575 52318 68609 52334
rect 67670 52230 67700 52272
rect 67610 52100 67700 52230
rect 68670 52272 68678 52430
rect 68670 52230 68700 52272
rect 68740 52230 68760 52470
rect 68670 52100 68760 52230
rect 72600 52790 72690 52910
rect 72600 52530 72620 52790
rect 72660 52740 72690 52790
rect 72680 52582 72690 52740
rect 73660 52790 73750 52910
rect 73660 52740 73690 52790
rect 72748 52678 72782 52694
rect 72816 52688 72832 52722
rect 73008 52688 73024 52722
rect 73314 52688 73330 52722
rect 73506 52688 73522 52722
rect 72748 52628 72782 52644
rect 73565 52678 73599 52694
rect 72816 52600 72832 52634
rect 73008 52600 73024 52634
rect 73314 52600 73330 52634
rect 73506 52600 73522 52634
rect 73565 52628 73599 52644
rect 72660 52530 72690 52582
rect 72600 52470 72690 52530
rect 72600 52230 72620 52470
rect 72660 52430 72690 52470
rect 72680 52272 72690 52430
rect 73660 52582 73668 52740
rect 73660 52550 73690 52582
rect 73730 52550 73750 52790
rect 73660 52470 73750 52550
rect 73660 52430 73690 52470
rect 72748 52368 72782 52384
rect 72816 52378 72832 52412
rect 73008 52378 73024 52412
rect 73314 52378 73330 52412
rect 73506 52378 73522 52412
rect 72748 52318 72782 52334
rect 73565 52368 73599 52384
rect 72816 52290 72832 52324
rect 73008 52290 73024 52324
rect 73314 52290 73330 52324
rect 73506 52290 73522 52324
rect 73565 52318 73599 52334
rect 72660 52230 72690 52272
rect 72600 52100 72690 52230
rect 73660 52272 73668 52430
rect 73660 52230 73690 52272
rect 73730 52230 73750 52470
rect 73660 52100 73750 52230
rect 77590 52790 77680 52910
rect 77590 52530 77610 52790
rect 77650 52740 77680 52790
rect 77670 52582 77680 52740
rect 78650 52790 78740 52910
rect 78650 52740 78680 52790
rect 77738 52678 77772 52694
rect 77806 52688 77822 52722
rect 77998 52688 78014 52722
rect 78304 52688 78320 52722
rect 78496 52688 78512 52722
rect 77738 52628 77772 52644
rect 78555 52678 78589 52694
rect 77806 52600 77822 52634
rect 77998 52600 78014 52634
rect 78304 52600 78320 52634
rect 78496 52600 78512 52634
rect 78555 52628 78589 52644
rect 77650 52530 77680 52582
rect 77590 52470 77680 52530
rect 77590 52230 77610 52470
rect 77650 52430 77680 52470
rect 77670 52272 77680 52430
rect 78650 52582 78658 52740
rect 78650 52550 78680 52582
rect 78720 52550 78740 52790
rect 78650 52470 78740 52550
rect 78650 52430 78680 52470
rect 77738 52368 77772 52384
rect 77806 52378 77822 52412
rect 77998 52378 78014 52412
rect 78304 52378 78320 52412
rect 78496 52378 78512 52412
rect 77738 52318 77772 52334
rect 78555 52368 78589 52384
rect 77806 52290 77822 52324
rect 77998 52290 78014 52324
rect 78304 52290 78320 52324
rect 78496 52290 78512 52324
rect 78555 52318 78589 52334
rect 77650 52230 77680 52272
rect 77590 52100 77680 52230
rect 78650 52272 78658 52430
rect 78650 52230 78680 52272
rect 78720 52230 78740 52470
rect 78650 52100 78740 52230
rect 2740 51080 2830 51200
rect 2740 50820 2760 51080
rect 2800 51030 2830 51080
rect 2820 50872 2830 51030
rect 3800 51080 3890 51200
rect 3800 51030 3830 51080
rect 2888 50968 2922 50984
rect 2956 50978 2972 51012
rect 3148 50978 3164 51012
rect 3454 50978 3470 51012
rect 3646 50978 3662 51012
rect 2888 50918 2922 50934
rect 3705 50968 3739 50984
rect 2956 50890 2972 50924
rect 3148 50890 3164 50924
rect 3454 50890 3470 50924
rect 3646 50890 3662 50924
rect 3705 50918 3739 50934
rect 2800 50820 2830 50872
rect 2740 50760 2830 50820
rect 2740 50520 2760 50760
rect 2800 50720 2830 50760
rect 2820 50562 2830 50720
rect 3800 50872 3808 51030
rect 3800 50840 3830 50872
rect 3870 50840 3890 51080
rect 3800 50760 3890 50840
rect 3800 50720 3830 50760
rect 2888 50658 2922 50674
rect 2956 50668 2972 50702
rect 3148 50668 3164 50702
rect 3454 50668 3470 50702
rect 3646 50668 3662 50702
rect 2888 50608 2922 50624
rect 3705 50658 3739 50674
rect 2956 50580 2972 50614
rect 3148 50580 3164 50614
rect 3454 50580 3470 50614
rect 3646 50580 3662 50614
rect 3705 50608 3739 50624
rect 2800 50520 2830 50562
rect 2740 50390 2830 50520
rect 3800 50562 3808 50720
rect 3800 50520 3830 50562
rect 3870 50520 3890 50760
rect 3800 50390 3890 50520
rect 7730 51080 7820 51200
rect 7730 50820 7750 51080
rect 7790 51030 7820 51080
rect 7810 50872 7820 51030
rect 8790 51080 8880 51200
rect 8790 51030 8820 51080
rect 7878 50968 7912 50984
rect 7946 50978 7962 51012
rect 8138 50978 8154 51012
rect 8444 50978 8460 51012
rect 8636 50978 8652 51012
rect 7878 50918 7912 50934
rect 8695 50968 8729 50984
rect 7946 50890 7962 50924
rect 8138 50890 8154 50924
rect 8444 50890 8460 50924
rect 8636 50890 8652 50924
rect 8695 50918 8729 50934
rect 7790 50820 7820 50872
rect 7730 50760 7820 50820
rect 7730 50520 7750 50760
rect 7790 50720 7820 50760
rect 7810 50562 7820 50720
rect 8790 50872 8798 51030
rect 8790 50840 8820 50872
rect 8860 50840 8880 51080
rect 8790 50760 8880 50840
rect 8790 50720 8820 50760
rect 7878 50658 7912 50674
rect 7946 50668 7962 50702
rect 8138 50668 8154 50702
rect 8444 50668 8460 50702
rect 8636 50668 8652 50702
rect 7878 50608 7912 50624
rect 8695 50658 8729 50674
rect 7946 50580 7962 50614
rect 8138 50580 8154 50614
rect 8444 50580 8460 50614
rect 8636 50580 8652 50614
rect 8695 50608 8729 50624
rect 7790 50520 7820 50562
rect 7730 50390 7820 50520
rect 8790 50562 8798 50720
rect 8790 50520 8820 50562
rect 8860 50520 8880 50760
rect 8790 50390 8880 50520
rect 12720 51080 12810 51200
rect 12720 50820 12740 51080
rect 12780 51030 12810 51080
rect 12800 50872 12810 51030
rect 13780 51080 13870 51200
rect 13780 51030 13810 51080
rect 12868 50968 12902 50984
rect 12936 50978 12952 51012
rect 13128 50978 13144 51012
rect 13434 50978 13450 51012
rect 13626 50978 13642 51012
rect 12868 50918 12902 50934
rect 13685 50968 13719 50984
rect 12936 50890 12952 50924
rect 13128 50890 13144 50924
rect 13434 50890 13450 50924
rect 13626 50890 13642 50924
rect 13685 50918 13719 50934
rect 12780 50820 12810 50872
rect 12720 50760 12810 50820
rect 12720 50520 12740 50760
rect 12780 50720 12810 50760
rect 12800 50562 12810 50720
rect 13780 50872 13788 51030
rect 13780 50840 13810 50872
rect 13850 50840 13870 51080
rect 13780 50760 13870 50840
rect 13780 50720 13810 50760
rect 12868 50658 12902 50674
rect 12936 50668 12952 50702
rect 13128 50668 13144 50702
rect 13434 50668 13450 50702
rect 13626 50668 13642 50702
rect 12868 50608 12902 50624
rect 13685 50658 13719 50674
rect 12936 50580 12952 50614
rect 13128 50580 13144 50614
rect 13434 50580 13450 50614
rect 13626 50580 13642 50614
rect 13685 50608 13719 50624
rect 12780 50520 12810 50562
rect 12720 50390 12810 50520
rect 13780 50562 13788 50720
rect 13780 50520 13810 50562
rect 13850 50520 13870 50760
rect 13780 50390 13870 50520
rect 17710 51080 17800 51200
rect 17710 50820 17730 51080
rect 17770 51030 17800 51080
rect 17790 50872 17800 51030
rect 18770 51080 18860 51200
rect 18770 51030 18800 51080
rect 17858 50968 17892 50984
rect 17926 50978 17942 51012
rect 18118 50978 18134 51012
rect 18424 50978 18440 51012
rect 18616 50978 18632 51012
rect 17858 50918 17892 50934
rect 18675 50968 18709 50984
rect 17926 50890 17942 50924
rect 18118 50890 18134 50924
rect 18424 50890 18440 50924
rect 18616 50890 18632 50924
rect 18675 50918 18709 50934
rect 17770 50820 17800 50872
rect 17710 50760 17800 50820
rect 17710 50520 17730 50760
rect 17770 50720 17800 50760
rect 17790 50562 17800 50720
rect 18770 50872 18778 51030
rect 18770 50840 18800 50872
rect 18840 50840 18860 51080
rect 18770 50760 18860 50840
rect 18770 50720 18800 50760
rect 17858 50658 17892 50674
rect 17926 50668 17942 50702
rect 18118 50668 18134 50702
rect 18424 50668 18440 50702
rect 18616 50668 18632 50702
rect 17858 50608 17892 50624
rect 18675 50658 18709 50674
rect 17926 50580 17942 50614
rect 18118 50580 18134 50614
rect 18424 50580 18440 50614
rect 18616 50580 18632 50614
rect 18675 50608 18709 50624
rect 17770 50520 17800 50562
rect 17710 50390 17800 50520
rect 18770 50562 18778 50720
rect 18770 50520 18800 50562
rect 18840 50520 18860 50760
rect 18770 50390 18860 50520
rect 22700 51080 22790 51200
rect 22700 50820 22720 51080
rect 22760 51030 22790 51080
rect 22780 50872 22790 51030
rect 23760 51080 23850 51200
rect 23760 51030 23790 51080
rect 22848 50968 22882 50984
rect 22916 50978 22932 51012
rect 23108 50978 23124 51012
rect 23414 50978 23430 51012
rect 23606 50978 23622 51012
rect 22848 50918 22882 50934
rect 23665 50968 23699 50984
rect 22916 50890 22932 50924
rect 23108 50890 23124 50924
rect 23414 50890 23430 50924
rect 23606 50890 23622 50924
rect 23665 50918 23699 50934
rect 22760 50820 22790 50872
rect 22700 50760 22790 50820
rect 22700 50520 22720 50760
rect 22760 50720 22790 50760
rect 22780 50562 22790 50720
rect 23760 50872 23768 51030
rect 23760 50840 23790 50872
rect 23830 50840 23850 51080
rect 23760 50760 23850 50840
rect 23760 50720 23790 50760
rect 22848 50658 22882 50674
rect 22916 50668 22932 50702
rect 23108 50668 23124 50702
rect 23414 50668 23430 50702
rect 23606 50668 23622 50702
rect 22848 50608 22882 50624
rect 23665 50658 23699 50674
rect 22916 50580 22932 50614
rect 23108 50580 23124 50614
rect 23414 50580 23430 50614
rect 23606 50580 23622 50614
rect 23665 50608 23699 50624
rect 22760 50520 22790 50562
rect 22700 50390 22790 50520
rect 23760 50562 23768 50720
rect 23760 50520 23790 50562
rect 23830 50520 23850 50760
rect 23760 50390 23850 50520
rect 27690 51080 27780 51200
rect 27690 50820 27710 51080
rect 27750 51030 27780 51080
rect 27770 50872 27780 51030
rect 28750 51080 28840 51200
rect 28750 51030 28780 51080
rect 27838 50968 27872 50984
rect 27906 50978 27922 51012
rect 28098 50978 28114 51012
rect 28404 50978 28420 51012
rect 28596 50978 28612 51012
rect 27838 50918 27872 50934
rect 28655 50968 28689 50984
rect 27906 50890 27922 50924
rect 28098 50890 28114 50924
rect 28404 50890 28420 50924
rect 28596 50890 28612 50924
rect 28655 50918 28689 50934
rect 27750 50820 27780 50872
rect 27690 50760 27780 50820
rect 27690 50520 27710 50760
rect 27750 50720 27780 50760
rect 27770 50562 27780 50720
rect 28750 50872 28758 51030
rect 28750 50840 28780 50872
rect 28820 50840 28840 51080
rect 28750 50760 28840 50840
rect 28750 50720 28780 50760
rect 27838 50658 27872 50674
rect 27906 50668 27922 50702
rect 28098 50668 28114 50702
rect 28404 50668 28420 50702
rect 28596 50668 28612 50702
rect 27838 50608 27872 50624
rect 28655 50658 28689 50674
rect 27906 50580 27922 50614
rect 28098 50580 28114 50614
rect 28404 50580 28420 50614
rect 28596 50580 28612 50614
rect 28655 50608 28689 50624
rect 27750 50520 27780 50562
rect 27690 50390 27780 50520
rect 28750 50562 28758 50720
rect 28750 50520 28780 50562
rect 28820 50520 28840 50760
rect 28750 50390 28840 50520
rect 32680 51080 32770 51200
rect 32680 50820 32700 51080
rect 32740 51030 32770 51080
rect 32760 50872 32770 51030
rect 33740 51080 33830 51200
rect 33740 51030 33770 51080
rect 32828 50968 32862 50984
rect 32896 50978 32912 51012
rect 33088 50978 33104 51012
rect 33394 50978 33410 51012
rect 33586 50978 33602 51012
rect 32828 50918 32862 50934
rect 33645 50968 33679 50984
rect 32896 50890 32912 50924
rect 33088 50890 33104 50924
rect 33394 50890 33410 50924
rect 33586 50890 33602 50924
rect 33645 50918 33679 50934
rect 32740 50820 32770 50872
rect 32680 50760 32770 50820
rect 32680 50520 32700 50760
rect 32740 50720 32770 50760
rect 32760 50562 32770 50720
rect 33740 50872 33748 51030
rect 33740 50840 33770 50872
rect 33810 50840 33830 51080
rect 33740 50760 33830 50840
rect 33740 50720 33770 50760
rect 32828 50658 32862 50674
rect 32896 50668 32912 50702
rect 33088 50668 33104 50702
rect 33394 50668 33410 50702
rect 33586 50668 33602 50702
rect 32828 50608 32862 50624
rect 33645 50658 33679 50674
rect 32896 50580 32912 50614
rect 33088 50580 33104 50614
rect 33394 50580 33410 50614
rect 33586 50580 33602 50614
rect 33645 50608 33679 50624
rect 32740 50520 32770 50562
rect 32680 50390 32770 50520
rect 33740 50562 33748 50720
rect 33740 50520 33770 50562
rect 33810 50520 33830 50760
rect 33740 50390 33830 50520
rect 37670 51080 37760 51200
rect 37670 50820 37690 51080
rect 37730 51030 37760 51080
rect 37750 50872 37760 51030
rect 38730 51080 38820 51200
rect 38730 51030 38760 51080
rect 37818 50968 37852 50984
rect 37886 50978 37902 51012
rect 38078 50978 38094 51012
rect 38384 50978 38400 51012
rect 38576 50978 38592 51012
rect 37818 50918 37852 50934
rect 38635 50968 38669 50984
rect 37886 50890 37902 50924
rect 38078 50890 38094 50924
rect 38384 50890 38400 50924
rect 38576 50890 38592 50924
rect 38635 50918 38669 50934
rect 37730 50820 37760 50872
rect 37670 50760 37760 50820
rect 37670 50520 37690 50760
rect 37730 50720 37760 50760
rect 37750 50562 37760 50720
rect 38730 50872 38738 51030
rect 38730 50840 38760 50872
rect 38800 50840 38820 51080
rect 38730 50760 38820 50840
rect 38730 50720 38760 50760
rect 37818 50658 37852 50674
rect 37886 50668 37902 50702
rect 38078 50668 38094 50702
rect 38384 50668 38400 50702
rect 38576 50668 38592 50702
rect 37818 50608 37852 50624
rect 38635 50658 38669 50674
rect 37886 50580 37902 50614
rect 38078 50580 38094 50614
rect 38384 50580 38400 50614
rect 38576 50580 38592 50614
rect 38635 50608 38669 50624
rect 37730 50520 37760 50562
rect 37670 50390 37760 50520
rect 38730 50562 38738 50720
rect 38730 50520 38760 50562
rect 38800 50520 38820 50760
rect 38730 50390 38820 50520
rect 42660 51080 42750 51200
rect 42660 50820 42680 51080
rect 42720 51030 42750 51080
rect 42740 50872 42750 51030
rect 43720 51080 43810 51200
rect 43720 51030 43750 51080
rect 42808 50968 42842 50984
rect 42876 50978 42892 51012
rect 43068 50978 43084 51012
rect 43374 50978 43390 51012
rect 43566 50978 43582 51012
rect 42808 50918 42842 50934
rect 43625 50968 43659 50984
rect 42876 50890 42892 50924
rect 43068 50890 43084 50924
rect 43374 50890 43390 50924
rect 43566 50890 43582 50924
rect 43625 50918 43659 50934
rect 42720 50820 42750 50872
rect 42660 50760 42750 50820
rect 42660 50520 42680 50760
rect 42720 50720 42750 50760
rect 42740 50562 42750 50720
rect 43720 50872 43728 51030
rect 43720 50840 43750 50872
rect 43790 50840 43810 51080
rect 43720 50760 43810 50840
rect 43720 50720 43750 50760
rect 42808 50658 42842 50674
rect 42876 50668 42892 50702
rect 43068 50668 43084 50702
rect 43374 50668 43390 50702
rect 43566 50668 43582 50702
rect 42808 50608 42842 50624
rect 43625 50658 43659 50674
rect 42876 50580 42892 50614
rect 43068 50580 43084 50614
rect 43374 50580 43390 50614
rect 43566 50580 43582 50614
rect 43625 50608 43659 50624
rect 42720 50520 42750 50562
rect 42660 50390 42750 50520
rect 43720 50562 43728 50720
rect 43720 50520 43750 50562
rect 43790 50520 43810 50760
rect 43720 50390 43810 50520
rect 47650 51080 47740 51200
rect 47650 50820 47670 51080
rect 47710 51030 47740 51080
rect 47730 50872 47740 51030
rect 48710 51080 48800 51200
rect 48710 51030 48740 51080
rect 47798 50968 47832 50984
rect 47866 50978 47882 51012
rect 48058 50978 48074 51012
rect 48364 50978 48380 51012
rect 48556 50978 48572 51012
rect 47798 50918 47832 50934
rect 48615 50968 48649 50984
rect 47866 50890 47882 50924
rect 48058 50890 48074 50924
rect 48364 50890 48380 50924
rect 48556 50890 48572 50924
rect 48615 50918 48649 50934
rect 47710 50820 47740 50872
rect 47650 50760 47740 50820
rect 47650 50520 47670 50760
rect 47710 50720 47740 50760
rect 47730 50562 47740 50720
rect 48710 50872 48718 51030
rect 48710 50840 48740 50872
rect 48780 50840 48800 51080
rect 48710 50760 48800 50840
rect 48710 50720 48740 50760
rect 47798 50658 47832 50674
rect 47866 50668 47882 50702
rect 48058 50668 48074 50702
rect 48364 50668 48380 50702
rect 48556 50668 48572 50702
rect 47798 50608 47832 50624
rect 48615 50658 48649 50674
rect 47866 50580 47882 50614
rect 48058 50580 48074 50614
rect 48364 50580 48380 50614
rect 48556 50580 48572 50614
rect 48615 50608 48649 50624
rect 47710 50520 47740 50562
rect 47650 50390 47740 50520
rect 48710 50562 48718 50720
rect 48710 50520 48740 50562
rect 48780 50520 48800 50760
rect 48710 50390 48800 50520
rect 52640 51080 52730 51200
rect 52640 50820 52660 51080
rect 52700 51030 52730 51080
rect 52720 50872 52730 51030
rect 53700 51080 53790 51200
rect 53700 51030 53730 51080
rect 52788 50968 52822 50984
rect 52856 50978 52872 51012
rect 53048 50978 53064 51012
rect 53354 50978 53370 51012
rect 53546 50978 53562 51012
rect 52788 50918 52822 50934
rect 53605 50968 53639 50984
rect 52856 50890 52872 50924
rect 53048 50890 53064 50924
rect 53354 50890 53370 50924
rect 53546 50890 53562 50924
rect 53605 50918 53639 50934
rect 52700 50820 52730 50872
rect 52640 50760 52730 50820
rect 52640 50520 52660 50760
rect 52700 50720 52730 50760
rect 52720 50562 52730 50720
rect 53700 50872 53708 51030
rect 53700 50840 53730 50872
rect 53770 50840 53790 51080
rect 53700 50760 53790 50840
rect 53700 50720 53730 50760
rect 52788 50658 52822 50674
rect 52856 50668 52872 50702
rect 53048 50668 53064 50702
rect 53354 50668 53370 50702
rect 53546 50668 53562 50702
rect 52788 50608 52822 50624
rect 53605 50658 53639 50674
rect 52856 50580 52872 50614
rect 53048 50580 53064 50614
rect 53354 50580 53370 50614
rect 53546 50580 53562 50614
rect 53605 50608 53639 50624
rect 52700 50520 52730 50562
rect 52640 50390 52730 50520
rect 53700 50562 53708 50720
rect 53700 50520 53730 50562
rect 53770 50520 53790 50760
rect 53700 50390 53790 50520
rect 57630 51080 57720 51200
rect 57630 50820 57650 51080
rect 57690 51030 57720 51080
rect 57710 50872 57720 51030
rect 58690 51080 58780 51200
rect 58690 51030 58720 51080
rect 57778 50968 57812 50984
rect 57846 50978 57862 51012
rect 58038 50978 58054 51012
rect 58344 50978 58360 51012
rect 58536 50978 58552 51012
rect 57778 50918 57812 50934
rect 58595 50968 58629 50984
rect 57846 50890 57862 50924
rect 58038 50890 58054 50924
rect 58344 50890 58360 50924
rect 58536 50890 58552 50924
rect 58595 50918 58629 50934
rect 57690 50820 57720 50872
rect 57630 50760 57720 50820
rect 57630 50520 57650 50760
rect 57690 50720 57720 50760
rect 57710 50562 57720 50720
rect 58690 50872 58698 51030
rect 58690 50840 58720 50872
rect 58760 50840 58780 51080
rect 58690 50760 58780 50840
rect 58690 50720 58720 50760
rect 57778 50658 57812 50674
rect 57846 50668 57862 50702
rect 58038 50668 58054 50702
rect 58344 50668 58360 50702
rect 58536 50668 58552 50702
rect 57778 50608 57812 50624
rect 58595 50658 58629 50674
rect 57846 50580 57862 50614
rect 58038 50580 58054 50614
rect 58344 50580 58360 50614
rect 58536 50580 58552 50614
rect 58595 50608 58629 50624
rect 57690 50520 57720 50562
rect 57630 50390 57720 50520
rect 58690 50562 58698 50720
rect 58690 50520 58720 50562
rect 58760 50520 58780 50760
rect 58690 50390 58780 50520
rect 62620 51080 62710 51200
rect 62620 50820 62640 51080
rect 62680 51030 62710 51080
rect 62700 50872 62710 51030
rect 63680 51080 63770 51200
rect 63680 51030 63710 51080
rect 62768 50968 62802 50984
rect 62836 50978 62852 51012
rect 63028 50978 63044 51012
rect 63334 50978 63350 51012
rect 63526 50978 63542 51012
rect 62768 50918 62802 50934
rect 63585 50968 63619 50984
rect 62836 50890 62852 50924
rect 63028 50890 63044 50924
rect 63334 50890 63350 50924
rect 63526 50890 63542 50924
rect 63585 50918 63619 50934
rect 62680 50820 62710 50872
rect 62620 50760 62710 50820
rect 62620 50520 62640 50760
rect 62680 50720 62710 50760
rect 62700 50562 62710 50720
rect 63680 50872 63688 51030
rect 63680 50840 63710 50872
rect 63750 50840 63770 51080
rect 63680 50760 63770 50840
rect 63680 50720 63710 50760
rect 62768 50658 62802 50674
rect 62836 50668 62852 50702
rect 63028 50668 63044 50702
rect 63334 50668 63350 50702
rect 63526 50668 63542 50702
rect 62768 50608 62802 50624
rect 63585 50658 63619 50674
rect 62836 50580 62852 50614
rect 63028 50580 63044 50614
rect 63334 50580 63350 50614
rect 63526 50580 63542 50614
rect 63585 50608 63619 50624
rect 62680 50520 62710 50562
rect 62620 50390 62710 50520
rect 63680 50562 63688 50720
rect 63680 50520 63710 50562
rect 63750 50520 63770 50760
rect 63680 50390 63770 50520
rect 67610 51080 67700 51200
rect 67610 50820 67630 51080
rect 67670 51030 67700 51080
rect 67690 50872 67700 51030
rect 68670 51080 68760 51200
rect 68670 51030 68700 51080
rect 67758 50968 67792 50984
rect 67826 50978 67842 51012
rect 68018 50978 68034 51012
rect 68324 50978 68340 51012
rect 68516 50978 68532 51012
rect 67758 50918 67792 50934
rect 68575 50968 68609 50984
rect 67826 50890 67842 50924
rect 68018 50890 68034 50924
rect 68324 50890 68340 50924
rect 68516 50890 68532 50924
rect 68575 50918 68609 50934
rect 67670 50820 67700 50872
rect 67610 50760 67700 50820
rect 67610 50520 67630 50760
rect 67670 50720 67700 50760
rect 67690 50562 67700 50720
rect 68670 50872 68678 51030
rect 68670 50840 68700 50872
rect 68740 50840 68760 51080
rect 68670 50760 68760 50840
rect 68670 50720 68700 50760
rect 67758 50658 67792 50674
rect 67826 50668 67842 50702
rect 68018 50668 68034 50702
rect 68324 50668 68340 50702
rect 68516 50668 68532 50702
rect 67758 50608 67792 50624
rect 68575 50658 68609 50674
rect 67826 50580 67842 50614
rect 68018 50580 68034 50614
rect 68324 50580 68340 50614
rect 68516 50580 68532 50614
rect 68575 50608 68609 50624
rect 67670 50520 67700 50562
rect 67610 50390 67700 50520
rect 68670 50562 68678 50720
rect 68670 50520 68700 50562
rect 68740 50520 68760 50760
rect 68670 50390 68760 50520
rect 72600 51080 72690 51200
rect 72600 50820 72620 51080
rect 72660 51030 72690 51080
rect 72680 50872 72690 51030
rect 73660 51080 73750 51200
rect 73660 51030 73690 51080
rect 72748 50968 72782 50984
rect 72816 50978 72832 51012
rect 73008 50978 73024 51012
rect 73314 50978 73330 51012
rect 73506 50978 73522 51012
rect 72748 50918 72782 50934
rect 73565 50968 73599 50984
rect 72816 50890 72832 50924
rect 73008 50890 73024 50924
rect 73314 50890 73330 50924
rect 73506 50890 73522 50924
rect 73565 50918 73599 50934
rect 72660 50820 72690 50872
rect 72600 50760 72690 50820
rect 72600 50520 72620 50760
rect 72660 50720 72690 50760
rect 72680 50562 72690 50720
rect 73660 50872 73668 51030
rect 73660 50840 73690 50872
rect 73730 50840 73750 51080
rect 73660 50760 73750 50840
rect 73660 50720 73690 50760
rect 72748 50658 72782 50674
rect 72816 50668 72832 50702
rect 73008 50668 73024 50702
rect 73314 50668 73330 50702
rect 73506 50668 73522 50702
rect 72748 50608 72782 50624
rect 73565 50658 73599 50674
rect 72816 50580 72832 50614
rect 73008 50580 73024 50614
rect 73314 50580 73330 50614
rect 73506 50580 73522 50614
rect 73565 50608 73599 50624
rect 72660 50520 72690 50562
rect 72600 50390 72690 50520
rect 73660 50562 73668 50720
rect 73660 50520 73690 50562
rect 73730 50520 73750 50760
rect 73660 50390 73750 50520
rect 77590 51080 77680 51200
rect 77590 50820 77610 51080
rect 77650 51030 77680 51080
rect 77670 50872 77680 51030
rect 78650 51080 78740 51200
rect 78650 51030 78680 51080
rect 77738 50968 77772 50984
rect 77806 50978 77822 51012
rect 77998 50978 78014 51012
rect 78304 50978 78320 51012
rect 78496 50978 78512 51012
rect 77738 50918 77772 50934
rect 78555 50968 78589 50984
rect 77806 50890 77822 50924
rect 77998 50890 78014 50924
rect 78304 50890 78320 50924
rect 78496 50890 78512 50924
rect 78555 50918 78589 50934
rect 77650 50820 77680 50872
rect 77590 50760 77680 50820
rect 77590 50520 77610 50760
rect 77650 50720 77680 50760
rect 77670 50562 77680 50720
rect 78650 50872 78658 51030
rect 78650 50840 78680 50872
rect 78720 50840 78740 51080
rect 78650 50760 78740 50840
rect 78650 50720 78680 50760
rect 77738 50658 77772 50674
rect 77806 50668 77822 50702
rect 77998 50668 78014 50702
rect 78304 50668 78320 50702
rect 78496 50668 78512 50702
rect 77738 50608 77772 50624
rect 78555 50658 78589 50674
rect 77806 50580 77822 50614
rect 77998 50580 78014 50614
rect 78304 50580 78320 50614
rect 78496 50580 78512 50614
rect 78555 50608 78589 50624
rect 77650 50520 77680 50562
rect 77590 50390 77680 50520
rect 78650 50562 78658 50720
rect 78650 50520 78680 50562
rect 78720 50520 78740 50760
rect 78650 50390 78740 50520
rect 2740 49370 2830 49490
rect 2740 49110 2760 49370
rect 2800 49320 2830 49370
rect 2820 49162 2830 49320
rect 3800 49370 3890 49490
rect 3800 49320 3830 49370
rect 2888 49258 2922 49274
rect 2956 49268 2972 49302
rect 3148 49268 3164 49302
rect 3454 49268 3470 49302
rect 3646 49268 3662 49302
rect 2888 49208 2922 49224
rect 3705 49258 3739 49274
rect 2956 49180 2972 49214
rect 3148 49180 3164 49214
rect 3454 49180 3470 49214
rect 3646 49180 3662 49214
rect 3705 49208 3739 49224
rect 2800 49110 2830 49162
rect 2740 49050 2830 49110
rect 2740 48810 2760 49050
rect 2800 49010 2830 49050
rect 2820 48852 2830 49010
rect 3800 49162 3808 49320
rect 3800 49130 3830 49162
rect 3870 49130 3890 49370
rect 3800 49050 3890 49130
rect 3800 49010 3830 49050
rect 2888 48948 2922 48964
rect 2956 48958 2972 48992
rect 3148 48958 3164 48992
rect 3454 48958 3470 48992
rect 3646 48958 3662 48992
rect 2888 48898 2922 48914
rect 3705 48948 3739 48964
rect 2956 48870 2972 48904
rect 3148 48870 3164 48904
rect 3454 48870 3470 48904
rect 3646 48870 3662 48904
rect 3705 48898 3739 48914
rect 2800 48810 2830 48852
rect 2740 48680 2830 48810
rect 3800 48852 3808 49010
rect 3800 48810 3830 48852
rect 3870 48810 3890 49050
rect 3800 48680 3890 48810
rect 7730 49370 7820 49490
rect 7730 49110 7750 49370
rect 7790 49320 7820 49370
rect 7810 49162 7820 49320
rect 8790 49370 8880 49490
rect 8790 49320 8820 49370
rect 7878 49258 7912 49274
rect 7946 49268 7962 49302
rect 8138 49268 8154 49302
rect 8444 49268 8460 49302
rect 8636 49268 8652 49302
rect 7878 49208 7912 49224
rect 8695 49258 8729 49274
rect 7946 49180 7962 49214
rect 8138 49180 8154 49214
rect 8444 49180 8460 49214
rect 8636 49180 8652 49214
rect 8695 49208 8729 49224
rect 7790 49110 7820 49162
rect 7730 49050 7820 49110
rect 7730 48810 7750 49050
rect 7790 49010 7820 49050
rect 7810 48852 7820 49010
rect 8790 49162 8798 49320
rect 8790 49130 8820 49162
rect 8860 49130 8880 49370
rect 8790 49050 8880 49130
rect 8790 49010 8820 49050
rect 7878 48948 7912 48964
rect 7946 48958 7962 48992
rect 8138 48958 8154 48992
rect 8444 48958 8460 48992
rect 8636 48958 8652 48992
rect 7878 48898 7912 48914
rect 8695 48948 8729 48964
rect 7946 48870 7962 48904
rect 8138 48870 8154 48904
rect 8444 48870 8460 48904
rect 8636 48870 8652 48904
rect 8695 48898 8729 48914
rect 7790 48810 7820 48852
rect 7730 48680 7820 48810
rect 8790 48852 8798 49010
rect 8790 48810 8820 48852
rect 8860 48810 8880 49050
rect 8790 48680 8880 48810
rect 12720 49370 12810 49490
rect 12720 49110 12740 49370
rect 12780 49320 12810 49370
rect 12800 49162 12810 49320
rect 13780 49370 13870 49490
rect 13780 49320 13810 49370
rect 12868 49258 12902 49274
rect 12936 49268 12952 49302
rect 13128 49268 13144 49302
rect 13434 49268 13450 49302
rect 13626 49268 13642 49302
rect 12868 49208 12902 49224
rect 13685 49258 13719 49274
rect 12936 49180 12952 49214
rect 13128 49180 13144 49214
rect 13434 49180 13450 49214
rect 13626 49180 13642 49214
rect 13685 49208 13719 49224
rect 12780 49110 12810 49162
rect 12720 49050 12810 49110
rect 12720 48810 12740 49050
rect 12780 49010 12810 49050
rect 12800 48852 12810 49010
rect 13780 49162 13788 49320
rect 13780 49130 13810 49162
rect 13850 49130 13870 49370
rect 13780 49050 13870 49130
rect 13780 49010 13810 49050
rect 12868 48948 12902 48964
rect 12936 48958 12952 48992
rect 13128 48958 13144 48992
rect 13434 48958 13450 48992
rect 13626 48958 13642 48992
rect 12868 48898 12902 48914
rect 13685 48948 13719 48964
rect 12936 48870 12952 48904
rect 13128 48870 13144 48904
rect 13434 48870 13450 48904
rect 13626 48870 13642 48904
rect 13685 48898 13719 48914
rect 12780 48810 12810 48852
rect 12720 48680 12810 48810
rect 13780 48852 13788 49010
rect 13780 48810 13810 48852
rect 13850 48810 13870 49050
rect 13780 48680 13870 48810
rect 17710 49370 17800 49490
rect 17710 49110 17730 49370
rect 17770 49320 17800 49370
rect 17790 49162 17800 49320
rect 18770 49370 18860 49490
rect 18770 49320 18800 49370
rect 17858 49258 17892 49274
rect 17926 49268 17942 49302
rect 18118 49268 18134 49302
rect 18424 49268 18440 49302
rect 18616 49268 18632 49302
rect 17858 49208 17892 49224
rect 18675 49258 18709 49274
rect 17926 49180 17942 49214
rect 18118 49180 18134 49214
rect 18424 49180 18440 49214
rect 18616 49180 18632 49214
rect 18675 49208 18709 49224
rect 17770 49110 17800 49162
rect 17710 49050 17800 49110
rect 17710 48810 17730 49050
rect 17770 49010 17800 49050
rect 17790 48852 17800 49010
rect 18770 49162 18778 49320
rect 18770 49130 18800 49162
rect 18840 49130 18860 49370
rect 18770 49050 18860 49130
rect 18770 49010 18800 49050
rect 17858 48948 17892 48964
rect 17926 48958 17942 48992
rect 18118 48958 18134 48992
rect 18424 48958 18440 48992
rect 18616 48958 18632 48992
rect 17858 48898 17892 48914
rect 18675 48948 18709 48964
rect 17926 48870 17942 48904
rect 18118 48870 18134 48904
rect 18424 48870 18440 48904
rect 18616 48870 18632 48904
rect 18675 48898 18709 48914
rect 17770 48810 17800 48852
rect 17710 48680 17800 48810
rect 18770 48852 18778 49010
rect 18770 48810 18800 48852
rect 18840 48810 18860 49050
rect 18770 48680 18860 48810
rect 22700 49370 22790 49490
rect 22700 49110 22720 49370
rect 22760 49320 22790 49370
rect 22780 49162 22790 49320
rect 23760 49370 23850 49490
rect 23760 49320 23790 49370
rect 22848 49258 22882 49274
rect 22916 49268 22932 49302
rect 23108 49268 23124 49302
rect 23414 49268 23430 49302
rect 23606 49268 23622 49302
rect 22848 49208 22882 49224
rect 23665 49258 23699 49274
rect 22916 49180 22932 49214
rect 23108 49180 23124 49214
rect 23414 49180 23430 49214
rect 23606 49180 23622 49214
rect 23665 49208 23699 49224
rect 22760 49110 22790 49162
rect 22700 49050 22790 49110
rect 22700 48810 22720 49050
rect 22760 49010 22790 49050
rect 22780 48852 22790 49010
rect 23760 49162 23768 49320
rect 23760 49130 23790 49162
rect 23830 49130 23850 49370
rect 23760 49050 23850 49130
rect 23760 49010 23790 49050
rect 22848 48948 22882 48964
rect 22916 48958 22932 48992
rect 23108 48958 23124 48992
rect 23414 48958 23430 48992
rect 23606 48958 23622 48992
rect 22848 48898 22882 48914
rect 23665 48948 23699 48964
rect 22916 48870 22932 48904
rect 23108 48870 23124 48904
rect 23414 48870 23430 48904
rect 23606 48870 23622 48904
rect 23665 48898 23699 48914
rect 22760 48810 22790 48852
rect 22700 48680 22790 48810
rect 23760 48852 23768 49010
rect 23760 48810 23790 48852
rect 23830 48810 23850 49050
rect 23760 48680 23850 48810
rect 27690 49370 27780 49490
rect 27690 49110 27710 49370
rect 27750 49320 27780 49370
rect 27770 49162 27780 49320
rect 28750 49370 28840 49490
rect 28750 49320 28780 49370
rect 27838 49258 27872 49274
rect 27906 49268 27922 49302
rect 28098 49268 28114 49302
rect 28404 49268 28420 49302
rect 28596 49268 28612 49302
rect 27838 49208 27872 49224
rect 28655 49258 28689 49274
rect 27906 49180 27922 49214
rect 28098 49180 28114 49214
rect 28404 49180 28420 49214
rect 28596 49180 28612 49214
rect 28655 49208 28689 49224
rect 27750 49110 27780 49162
rect 27690 49050 27780 49110
rect 27690 48810 27710 49050
rect 27750 49010 27780 49050
rect 27770 48852 27780 49010
rect 28750 49162 28758 49320
rect 28750 49130 28780 49162
rect 28820 49130 28840 49370
rect 28750 49050 28840 49130
rect 28750 49010 28780 49050
rect 27838 48948 27872 48964
rect 27906 48958 27922 48992
rect 28098 48958 28114 48992
rect 28404 48958 28420 48992
rect 28596 48958 28612 48992
rect 27838 48898 27872 48914
rect 28655 48948 28689 48964
rect 27906 48870 27922 48904
rect 28098 48870 28114 48904
rect 28404 48870 28420 48904
rect 28596 48870 28612 48904
rect 28655 48898 28689 48914
rect 27750 48810 27780 48852
rect 27690 48680 27780 48810
rect 28750 48852 28758 49010
rect 28750 48810 28780 48852
rect 28820 48810 28840 49050
rect 28750 48680 28840 48810
rect 32680 49370 32770 49490
rect 32680 49110 32700 49370
rect 32740 49320 32770 49370
rect 32760 49162 32770 49320
rect 33740 49370 33830 49490
rect 33740 49320 33770 49370
rect 32828 49258 32862 49274
rect 32896 49268 32912 49302
rect 33088 49268 33104 49302
rect 33394 49268 33410 49302
rect 33586 49268 33602 49302
rect 32828 49208 32862 49224
rect 33645 49258 33679 49274
rect 32896 49180 32912 49214
rect 33088 49180 33104 49214
rect 33394 49180 33410 49214
rect 33586 49180 33602 49214
rect 33645 49208 33679 49224
rect 32740 49110 32770 49162
rect 32680 49050 32770 49110
rect 32680 48810 32700 49050
rect 32740 49010 32770 49050
rect 32760 48852 32770 49010
rect 33740 49162 33748 49320
rect 33740 49130 33770 49162
rect 33810 49130 33830 49370
rect 33740 49050 33830 49130
rect 33740 49010 33770 49050
rect 32828 48948 32862 48964
rect 32896 48958 32912 48992
rect 33088 48958 33104 48992
rect 33394 48958 33410 48992
rect 33586 48958 33602 48992
rect 32828 48898 32862 48914
rect 33645 48948 33679 48964
rect 32896 48870 32912 48904
rect 33088 48870 33104 48904
rect 33394 48870 33410 48904
rect 33586 48870 33602 48904
rect 33645 48898 33679 48914
rect 32740 48810 32770 48852
rect 32680 48680 32770 48810
rect 33740 48852 33748 49010
rect 33740 48810 33770 48852
rect 33810 48810 33830 49050
rect 33740 48680 33830 48810
rect 37670 49370 37760 49490
rect 37670 49110 37690 49370
rect 37730 49320 37760 49370
rect 37750 49162 37760 49320
rect 38730 49370 38820 49490
rect 38730 49320 38760 49370
rect 37818 49258 37852 49274
rect 37886 49268 37902 49302
rect 38078 49268 38094 49302
rect 38384 49268 38400 49302
rect 38576 49268 38592 49302
rect 37818 49208 37852 49224
rect 38635 49258 38669 49274
rect 37886 49180 37902 49214
rect 38078 49180 38094 49214
rect 38384 49180 38400 49214
rect 38576 49180 38592 49214
rect 38635 49208 38669 49224
rect 37730 49110 37760 49162
rect 37670 49050 37760 49110
rect 37670 48810 37690 49050
rect 37730 49010 37760 49050
rect 37750 48852 37760 49010
rect 38730 49162 38738 49320
rect 38730 49130 38760 49162
rect 38800 49130 38820 49370
rect 38730 49050 38820 49130
rect 38730 49010 38760 49050
rect 37818 48948 37852 48964
rect 37886 48958 37902 48992
rect 38078 48958 38094 48992
rect 38384 48958 38400 48992
rect 38576 48958 38592 48992
rect 37818 48898 37852 48914
rect 38635 48948 38669 48964
rect 37886 48870 37902 48904
rect 38078 48870 38094 48904
rect 38384 48870 38400 48904
rect 38576 48870 38592 48904
rect 38635 48898 38669 48914
rect 37730 48810 37760 48852
rect 37670 48680 37760 48810
rect 38730 48852 38738 49010
rect 38730 48810 38760 48852
rect 38800 48810 38820 49050
rect 38730 48680 38820 48810
rect 42660 49370 42750 49490
rect 42660 49110 42680 49370
rect 42720 49320 42750 49370
rect 42740 49162 42750 49320
rect 43720 49370 43810 49490
rect 43720 49320 43750 49370
rect 42808 49258 42842 49274
rect 42876 49268 42892 49302
rect 43068 49268 43084 49302
rect 43374 49268 43390 49302
rect 43566 49268 43582 49302
rect 42808 49208 42842 49224
rect 43625 49258 43659 49274
rect 42876 49180 42892 49214
rect 43068 49180 43084 49214
rect 43374 49180 43390 49214
rect 43566 49180 43582 49214
rect 43625 49208 43659 49224
rect 42720 49110 42750 49162
rect 42660 49050 42750 49110
rect 42660 48810 42680 49050
rect 42720 49010 42750 49050
rect 42740 48852 42750 49010
rect 43720 49162 43728 49320
rect 43720 49130 43750 49162
rect 43790 49130 43810 49370
rect 43720 49050 43810 49130
rect 43720 49010 43750 49050
rect 42808 48948 42842 48964
rect 42876 48958 42892 48992
rect 43068 48958 43084 48992
rect 43374 48958 43390 48992
rect 43566 48958 43582 48992
rect 42808 48898 42842 48914
rect 43625 48948 43659 48964
rect 42876 48870 42892 48904
rect 43068 48870 43084 48904
rect 43374 48870 43390 48904
rect 43566 48870 43582 48904
rect 43625 48898 43659 48914
rect 42720 48810 42750 48852
rect 42660 48680 42750 48810
rect 43720 48852 43728 49010
rect 43720 48810 43750 48852
rect 43790 48810 43810 49050
rect 43720 48680 43810 48810
rect 47650 49370 47740 49490
rect 47650 49110 47670 49370
rect 47710 49320 47740 49370
rect 47730 49162 47740 49320
rect 48710 49370 48800 49490
rect 48710 49320 48740 49370
rect 47798 49258 47832 49274
rect 47866 49268 47882 49302
rect 48058 49268 48074 49302
rect 48364 49268 48380 49302
rect 48556 49268 48572 49302
rect 47798 49208 47832 49224
rect 48615 49258 48649 49274
rect 47866 49180 47882 49214
rect 48058 49180 48074 49214
rect 48364 49180 48380 49214
rect 48556 49180 48572 49214
rect 48615 49208 48649 49224
rect 47710 49110 47740 49162
rect 47650 49050 47740 49110
rect 47650 48810 47670 49050
rect 47710 49010 47740 49050
rect 47730 48852 47740 49010
rect 48710 49162 48718 49320
rect 48710 49130 48740 49162
rect 48780 49130 48800 49370
rect 48710 49050 48800 49130
rect 48710 49010 48740 49050
rect 47798 48948 47832 48964
rect 47866 48958 47882 48992
rect 48058 48958 48074 48992
rect 48364 48958 48380 48992
rect 48556 48958 48572 48992
rect 47798 48898 47832 48914
rect 48615 48948 48649 48964
rect 47866 48870 47882 48904
rect 48058 48870 48074 48904
rect 48364 48870 48380 48904
rect 48556 48870 48572 48904
rect 48615 48898 48649 48914
rect 47710 48810 47740 48852
rect 47650 48680 47740 48810
rect 48710 48852 48718 49010
rect 48710 48810 48740 48852
rect 48780 48810 48800 49050
rect 48710 48680 48800 48810
rect 52640 49370 52730 49490
rect 52640 49110 52660 49370
rect 52700 49320 52730 49370
rect 52720 49162 52730 49320
rect 53700 49370 53790 49490
rect 53700 49320 53730 49370
rect 52788 49258 52822 49274
rect 52856 49268 52872 49302
rect 53048 49268 53064 49302
rect 53354 49268 53370 49302
rect 53546 49268 53562 49302
rect 52788 49208 52822 49224
rect 53605 49258 53639 49274
rect 52856 49180 52872 49214
rect 53048 49180 53064 49214
rect 53354 49180 53370 49214
rect 53546 49180 53562 49214
rect 53605 49208 53639 49224
rect 52700 49110 52730 49162
rect 52640 49050 52730 49110
rect 52640 48810 52660 49050
rect 52700 49010 52730 49050
rect 52720 48852 52730 49010
rect 53700 49162 53708 49320
rect 53700 49130 53730 49162
rect 53770 49130 53790 49370
rect 53700 49050 53790 49130
rect 53700 49010 53730 49050
rect 52788 48948 52822 48964
rect 52856 48958 52872 48992
rect 53048 48958 53064 48992
rect 53354 48958 53370 48992
rect 53546 48958 53562 48992
rect 52788 48898 52822 48914
rect 53605 48948 53639 48964
rect 52856 48870 52872 48904
rect 53048 48870 53064 48904
rect 53354 48870 53370 48904
rect 53546 48870 53562 48904
rect 53605 48898 53639 48914
rect 52700 48810 52730 48852
rect 52640 48680 52730 48810
rect 53700 48852 53708 49010
rect 53700 48810 53730 48852
rect 53770 48810 53790 49050
rect 53700 48680 53790 48810
rect 57630 49370 57720 49490
rect 57630 49110 57650 49370
rect 57690 49320 57720 49370
rect 57710 49162 57720 49320
rect 58690 49370 58780 49490
rect 58690 49320 58720 49370
rect 57778 49258 57812 49274
rect 57846 49268 57862 49302
rect 58038 49268 58054 49302
rect 58344 49268 58360 49302
rect 58536 49268 58552 49302
rect 57778 49208 57812 49224
rect 58595 49258 58629 49274
rect 57846 49180 57862 49214
rect 58038 49180 58054 49214
rect 58344 49180 58360 49214
rect 58536 49180 58552 49214
rect 58595 49208 58629 49224
rect 57690 49110 57720 49162
rect 57630 49050 57720 49110
rect 57630 48810 57650 49050
rect 57690 49010 57720 49050
rect 57710 48852 57720 49010
rect 58690 49162 58698 49320
rect 58690 49130 58720 49162
rect 58760 49130 58780 49370
rect 58690 49050 58780 49130
rect 58690 49010 58720 49050
rect 57778 48948 57812 48964
rect 57846 48958 57862 48992
rect 58038 48958 58054 48992
rect 58344 48958 58360 48992
rect 58536 48958 58552 48992
rect 57778 48898 57812 48914
rect 58595 48948 58629 48964
rect 57846 48870 57862 48904
rect 58038 48870 58054 48904
rect 58344 48870 58360 48904
rect 58536 48870 58552 48904
rect 58595 48898 58629 48914
rect 57690 48810 57720 48852
rect 57630 48680 57720 48810
rect 58690 48852 58698 49010
rect 58690 48810 58720 48852
rect 58760 48810 58780 49050
rect 58690 48680 58780 48810
rect 62620 49370 62710 49490
rect 62620 49110 62640 49370
rect 62680 49320 62710 49370
rect 62700 49162 62710 49320
rect 63680 49370 63770 49490
rect 63680 49320 63710 49370
rect 62768 49258 62802 49274
rect 62836 49268 62852 49302
rect 63028 49268 63044 49302
rect 63334 49268 63350 49302
rect 63526 49268 63542 49302
rect 62768 49208 62802 49224
rect 63585 49258 63619 49274
rect 62836 49180 62852 49214
rect 63028 49180 63044 49214
rect 63334 49180 63350 49214
rect 63526 49180 63542 49214
rect 63585 49208 63619 49224
rect 62680 49110 62710 49162
rect 62620 49050 62710 49110
rect 62620 48810 62640 49050
rect 62680 49010 62710 49050
rect 62700 48852 62710 49010
rect 63680 49162 63688 49320
rect 63680 49130 63710 49162
rect 63750 49130 63770 49370
rect 63680 49050 63770 49130
rect 63680 49010 63710 49050
rect 62768 48948 62802 48964
rect 62836 48958 62852 48992
rect 63028 48958 63044 48992
rect 63334 48958 63350 48992
rect 63526 48958 63542 48992
rect 62768 48898 62802 48914
rect 63585 48948 63619 48964
rect 62836 48870 62852 48904
rect 63028 48870 63044 48904
rect 63334 48870 63350 48904
rect 63526 48870 63542 48904
rect 63585 48898 63619 48914
rect 62680 48810 62710 48852
rect 62620 48680 62710 48810
rect 63680 48852 63688 49010
rect 63680 48810 63710 48852
rect 63750 48810 63770 49050
rect 63680 48680 63770 48810
rect 67610 49370 67700 49490
rect 67610 49110 67630 49370
rect 67670 49320 67700 49370
rect 67690 49162 67700 49320
rect 68670 49370 68760 49490
rect 68670 49320 68700 49370
rect 67758 49258 67792 49274
rect 67826 49268 67842 49302
rect 68018 49268 68034 49302
rect 68324 49268 68340 49302
rect 68516 49268 68532 49302
rect 67758 49208 67792 49224
rect 68575 49258 68609 49274
rect 67826 49180 67842 49214
rect 68018 49180 68034 49214
rect 68324 49180 68340 49214
rect 68516 49180 68532 49214
rect 68575 49208 68609 49224
rect 67670 49110 67700 49162
rect 67610 49050 67700 49110
rect 67610 48810 67630 49050
rect 67670 49010 67700 49050
rect 67690 48852 67700 49010
rect 68670 49162 68678 49320
rect 68670 49130 68700 49162
rect 68740 49130 68760 49370
rect 68670 49050 68760 49130
rect 68670 49010 68700 49050
rect 67758 48948 67792 48964
rect 67826 48958 67842 48992
rect 68018 48958 68034 48992
rect 68324 48958 68340 48992
rect 68516 48958 68532 48992
rect 67758 48898 67792 48914
rect 68575 48948 68609 48964
rect 67826 48870 67842 48904
rect 68018 48870 68034 48904
rect 68324 48870 68340 48904
rect 68516 48870 68532 48904
rect 68575 48898 68609 48914
rect 67670 48810 67700 48852
rect 67610 48680 67700 48810
rect 68670 48852 68678 49010
rect 68670 48810 68700 48852
rect 68740 48810 68760 49050
rect 68670 48680 68760 48810
rect 72600 49370 72690 49490
rect 72600 49110 72620 49370
rect 72660 49320 72690 49370
rect 72680 49162 72690 49320
rect 73660 49370 73750 49490
rect 73660 49320 73690 49370
rect 72748 49258 72782 49274
rect 72816 49268 72832 49302
rect 73008 49268 73024 49302
rect 73314 49268 73330 49302
rect 73506 49268 73522 49302
rect 72748 49208 72782 49224
rect 73565 49258 73599 49274
rect 72816 49180 72832 49214
rect 73008 49180 73024 49214
rect 73314 49180 73330 49214
rect 73506 49180 73522 49214
rect 73565 49208 73599 49224
rect 72660 49110 72690 49162
rect 72600 49050 72690 49110
rect 72600 48810 72620 49050
rect 72660 49010 72690 49050
rect 72680 48852 72690 49010
rect 73660 49162 73668 49320
rect 73660 49130 73690 49162
rect 73730 49130 73750 49370
rect 73660 49050 73750 49130
rect 73660 49010 73690 49050
rect 72748 48948 72782 48964
rect 72816 48958 72832 48992
rect 73008 48958 73024 48992
rect 73314 48958 73330 48992
rect 73506 48958 73522 48992
rect 72748 48898 72782 48914
rect 73565 48948 73599 48964
rect 72816 48870 72832 48904
rect 73008 48870 73024 48904
rect 73314 48870 73330 48904
rect 73506 48870 73522 48904
rect 73565 48898 73599 48914
rect 72660 48810 72690 48852
rect 72600 48680 72690 48810
rect 73660 48852 73668 49010
rect 73660 48810 73690 48852
rect 73730 48810 73750 49050
rect 73660 48680 73750 48810
rect 77590 49370 77680 49490
rect 77590 49110 77610 49370
rect 77650 49320 77680 49370
rect 77670 49162 77680 49320
rect 78650 49370 78740 49490
rect 78650 49320 78680 49370
rect 77738 49258 77772 49274
rect 77806 49268 77822 49302
rect 77998 49268 78014 49302
rect 78304 49268 78320 49302
rect 78496 49268 78512 49302
rect 77738 49208 77772 49224
rect 78555 49258 78589 49274
rect 77806 49180 77822 49214
rect 77998 49180 78014 49214
rect 78304 49180 78320 49214
rect 78496 49180 78512 49214
rect 78555 49208 78589 49224
rect 77650 49110 77680 49162
rect 77590 49050 77680 49110
rect 77590 48810 77610 49050
rect 77650 49010 77680 49050
rect 77670 48852 77680 49010
rect 78650 49162 78658 49320
rect 78650 49130 78680 49162
rect 78720 49130 78740 49370
rect 78650 49050 78740 49130
rect 78650 49010 78680 49050
rect 77738 48948 77772 48964
rect 77806 48958 77822 48992
rect 77998 48958 78014 48992
rect 78304 48958 78320 48992
rect 78496 48958 78512 48992
rect 77738 48898 77772 48914
rect 78555 48948 78589 48964
rect 77806 48870 77822 48904
rect 77998 48870 78014 48904
rect 78304 48870 78320 48904
rect 78496 48870 78512 48904
rect 78555 48898 78589 48914
rect 77650 48810 77680 48852
rect 77590 48680 77680 48810
rect 78650 48852 78658 49010
rect 78650 48810 78680 48852
rect 78720 48810 78740 49050
rect 78650 48680 78740 48810
rect 2740 47660 2830 47780
rect 2740 47400 2760 47660
rect 2800 47610 2830 47660
rect 2820 47452 2830 47610
rect 3800 47660 3890 47780
rect 3800 47610 3830 47660
rect 2888 47548 2922 47564
rect 2956 47558 2972 47592
rect 3148 47558 3164 47592
rect 3454 47558 3470 47592
rect 3646 47558 3662 47592
rect 2888 47498 2922 47514
rect 3705 47548 3739 47564
rect 2956 47470 2972 47504
rect 3148 47470 3164 47504
rect 3454 47470 3470 47504
rect 3646 47470 3662 47504
rect 3705 47498 3739 47514
rect 2800 47400 2830 47452
rect 2740 47340 2830 47400
rect 2740 47100 2760 47340
rect 2800 47300 2830 47340
rect 2820 47142 2830 47300
rect 3800 47452 3808 47610
rect 3800 47420 3830 47452
rect 3870 47420 3890 47660
rect 3800 47340 3890 47420
rect 3800 47300 3830 47340
rect 2888 47238 2922 47254
rect 2956 47248 2972 47282
rect 3148 47248 3164 47282
rect 3454 47248 3470 47282
rect 3646 47248 3662 47282
rect 2888 47188 2922 47204
rect 3705 47238 3739 47254
rect 2956 47160 2972 47194
rect 3148 47160 3164 47194
rect 3454 47160 3470 47194
rect 3646 47160 3662 47194
rect 3705 47188 3739 47204
rect 2800 47100 2830 47142
rect 2740 46970 2830 47100
rect 3800 47142 3808 47300
rect 3800 47100 3830 47142
rect 3870 47100 3890 47340
rect 3800 46970 3890 47100
rect 7730 47660 7820 47780
rect 7730 47400 7750 47660
rect 7790 47610 7820 47660
rect 7810 47452 7820 47610
rect 8790 47660 8880 47780
rect 8790 47610 8820 47660
rect 7878 47548 7912 47564
rect 7946 47558 7962 47592
rect 8138 47558 8154 47592
rect 8444 47558 8460 47592
rect 8636 47558 8652 47592
rect 7878 47498 7912 47514
rect 8695 47548 8729 47564
rect 7946 47470 7962 47504
rect 8138 47470 8154 47504
rect 8444 47470 8460 47504
rect 8636 47470 8652 47504
rect 8695 47498 8729 47514
rect 7790 47400 7820 47452
rect 7730 47340 7820 47400
rect 7730 47100 7750 47340
rect 7790 47300 7820 47340
rect 7810 47142 7820 47300
rect 8790 47452 8798 47610
rect 8790 47420 8820 47452
rect 8860 47420 8880 47660
rect 8790 47340 8880 47420
rect 8790 47300 8820 47340
rect 7878 47238 7912 47254
rect 7946 47248 7962 47282
rect 8138 47248 8154 47282
rect 8444 47248 8460 47282
rect 8636 47248 8652 47282
rect 7878 47188 7912 47204
rect 8695 47238 8729 47254
rect 7946 47160 7962 47194
rect 8138 47160 8154 47194
rect 8444 47160 8460 47194
rect 8636 47160 8652 47194
rect 8695 47188 8729 47204
rect 7790 47100 7820 47142
rect 7730 46970 7820 47100
rect 8790 47142 8798 47300
rect 8790 47100 8820 47142
rect 8860 47100 8880 47340
rect 8790 46970 8880 47100
rect 12720 47660 12810 47780
rect 12720 47400 12740 47660
rect 12780 47610 12810 47660
rect 12800 47452 12810 47610
rect 13780 47660 13870 47780
rect 13780 47610 13810 47660
rect 12868 47548 12902 47564
rect 12936 47558 12952 47592
rect 13128 47558 13144 47592
rect 13434 47558 13450 47592
rect 13626 47558 13642 47592
rect 12868 47498 12902 47514
rect 13685 47548 13719 47564
rect 12936 47470 12952 47504
rect 13128 47470 13144 47504
rect 13434 47470 13450 47504
rect 13626 47470 13642 47504
rect 13685 47498 13719 47514
rect 12780 47400 12810 47452
rect 12720 47340 12810 47400
rect 12720 47100 12740 47340
rect 12780 47300 12810 47340
rect 12800 47142 12810 47300
rect 13780 47452 13788 47610
rect 13780 47420 13810 47452
rect 13850 47420 13870 47660
rect 13780 47340 13870 47420
rect 13780 47300 13810 47340
rect 12868 47238 12902 47254
rect 12936 47248 12952 47282
rect 13128 47248 13144 47282
rect 13434 47248 13450 47282
rect 13626 47248 13642 47282
rect 12868 47188 12902 47204
rect 13685 47238 13719 47254
rect 12936 47160 12952 47194
rect 13128 47160 13144 47194
rect 13434 47160 13450 47194
rect 13626 47160 13642 47194
rect 13685 47188 13719 47204
rect 12780 47100 12810 47142
rect 12720 46970 12810 47100
rect 13780 47142 13788 47300
rect 13780 47100 13810 47142
rect 13850 47100 13870 47340
rect 13780 46970 13870 47100
rect 17710 47660 17800 47780
rect 17710 47400 17730 47660
rect 17770 47610 17800 47660
rect 17790 47452 17800 47610
rect 18770 47660 18860 47780
rect 18770 47610 18800 47660
rect 17858 47548 17892 47564
rect 17926 47558 17942 47592
rect 18118 47558 18134 47592
rect 18424 47558 18440 47592
rect 18616 47558 18632 47592
rect 17858 47498 17892 47514
rect 18675 47548 18709 47564
rect 17926 47470 17942 47504
rect 18118 47470 18134 47504
rect 18424 47470 18440 47504
rect 18616 47470 18632 47504
rect 18675 47498 18709 47514
rect 17770 47400 17800 47452
rect 17710 47340 17800 47400
rect 17710 47100 17730 47340
rect 17770 47300 17800 47340
rect 17790 47142 17800 47300
rect 18770 47452 18778 47610
rect 18770 47420 18800 47452
rect 18840 47420 18860 47660
rect 18770 47340 18860 47420
rect 18770 47300 18800 47340
rect 17858 47238 17892 47254
rect 17926 47248 17942 47282
rect 18118 47248 18134 47282
rect 18424 47248 18440 47282
rect 18616 47248 18632 47282
rect 17858 47188 17892 47204
rect 18675 47238 18709 47254
rect 17926 47160 17942 47194
rect 18118 47160 18134 47194
rect 18424 47160 18440 47194
rect 18616 47160 18632 47194
rect 18675 47188 18709 47204
rect 17770 47100 17800 47142
rect 17710 46970 17800 47100
rect 18770 47142 18778 47300
rect 18770 47100 18800 47142
rect 18840 47100 18860 47340
rect 18770 46970 18860 47100
rect 22700 47660 22790 47780
rect 22700 47400 22720 47660
rect 22760 47610 22790 47660
rect 22780 47452 22790 47610
rect 23760 47660 23850 47780
rect 23760 47610 23790 47660
rect 22848 47548 22882 47564
rect 22916 47558 22932 47592
rect 23108 47558 23124 47592
rect 23414 47558 23430 47592
rect 23606 47558 23622 47592
rect 22848 47498 22882 47514
rect 23665 47548 23699 47564
rect 22916 47470 22932 47504
rect 23108 47470 23124 47504
rect 23414 47470 23430 47504
rect 23606 47470 23622 47504
rect 23665 47498 23699 47514
rect 22760 47400 22790 47452
rect 22700 47340 22790 47400
rect 22700 47100 22720 47340
rect 22760 47300 22790 47340
rect 22780 47142 22790 47300
rect 23760 47452 23768 47610
rect 23760 47420 23790 47452
rect 23830 47420 23850 47660
rect 23760 47340 23850 47420
rect 23760 47300 23790 47340
rect 22848 47238 22882 47254
rect 22916 47248 22932 47282
rect 23108 47248 23124 47282
rect 23414 47248 23430 47282
rect 23606 47248 23622 47282
rect 22848 47188 22882 47204
rect 23665 47238 23699 47254
rect 22916 47160 22932 47194
rect 23108 47160 23124 47194
rect 23414 47160 23430 47194
rect 23606 47160 23622 47194
rect 23665 47188 23699 47204
rect 22760 47100 22790 47142
rect 22700 46970 22790 47100
rect 23760 47142 23768 47300
rect 23760 47100 23790 47142
rect 23830 47100 23850 47340
rect 23760 46970 23850 47100
rect 27690 47660 27780 47780
rect 27690 47400 27710 47660
rect 27750 47610 27780 47660
rect 27770 47452 27780 47610
rect 28750 47660 28840 47780
rect 28750 47610 28780 47660
rect 27838 47548 27872 47564
rect 27906 47558 27922 47592
rect 28098 47558 28114 47592
rect 28404 47558 28420 47592
rect 28596 47558 28612 47592
rect 27838 47498 27872 47514
rect 28655 47548 28689 47564
rect 27906 47470 27922 47504
rect 28098 47470 28114 47504
rect 28404 47470 28420 47504
rect 28596 47470 28612 47504
rect 28655 47498 28689 47514
rect 27750 47400 27780 47452
rect 27690 47340 27780 47400
rect 27690 47100 27710 47340
rect 27750 47300 27780 47340
rect 27770 47142 27780 47300
rect 28750 47452 28758 47610
rect 28750 47420 28780 47452
rect 28820 47420 28840 47660
rect 28750 47340 28840 47420
rect 28750 47300 28780 47340
rect 27838 47238 27872 47254
rect 27906 47248 27922 47282
rect 28098 47248 28114 47282
rect 28404 47248 28420 47282
rect 28596 47248 28612 47282
rect 27838 47188 27872 47204
rect 28655 47238 28689 47254
rect 27906 47160 27922 47194
rect 28098 47160 28114 47194
rect 28404 47160 28420 47194
rect 28596 47160 28612 47194
rect 28655 47188 28689 47204
rect 27750 47100 27780 47142
rect 27690 46970 27780 47100
rect 28750 47142 28758 47300
rect 28750 47100 28780 47142
rect 28820 47100 28840 47340
rect 28750 46970 28840 47100
rect 32680 47660 32770 47780
rect 32680 47400 32700 47660
rect 32740 47610 32770 47660
rect 32760 47452 32770 47610
rect 33740 47660 33830 47780
rect 33740 47610 33770 47660
rect 32828 47548 32862 47564
rect 32896 47558 32912 47592
rect 33088 47558 33104 47592
rect 33394 47558 33410 47592
rect 33586 47558 33602 47592
rect 32828 47498 32862 47514
rect 33645 47548 33679 47564
rect 32896 47470 32912 47504
rect 33088 47470 33104 47504
rect 33394 47470 33410 47504
rect 33586 47470 33602 47504
rect 33645 47498 33679 47514
rect 32740 47400 32770 47452
rect 32680 47340 32770 47400
rect 32680 47100 32700 47340
rect 32740 47300 32770 47340
rect 32760 47142 32770 47300
rect 33740 47452 33748 47610
rect 33740 47420 33770 47452
rect 33810 47420 33830 47660
rect 33740 47340 33830 47420
rect 33740 47300 33770 47340
rect 32828 47238 32862 47254
rect 32896 47248 32912 47282
rect 33088 47248 33104 47282
rect 33394 47248 33410 47282
rect 33586 47248 33602 47282
rect 32828 47188 32862 47204
rect 33645 47238 33679 47254
rect 32896 47160 32912 47194
rect 33088 47160 33104 47194
rect 33394 47160 33410 47194
rect 33586 47160 33602 47194
rect 33645 47188 33679 47204
rect 32740 47100 32770 47142
rect 32680 46970 32770 47100
rect 33740 47142 33748 47300
rect 33740 47100 33770 47142
rect 33810 47100 33830 47340
rect 33740 46970 33830 47100
rect 37670 47660 37760 47780
rect 37670 47400 37690 47660
rect 37730 47610 37760 47660
rect 37750 47452 37760 47610
rect 38730 47660 38820 47780
rect 38730 47610 38760 47660
rect 37818 47548 37852 47564
rect 37886 47558 37902 47592
rect 38078 47558 38094 47592
rect 38384 47558 38400 47592
rect 38576 47558 38592 47592
rect 37818 47498 37852 47514
rect 38635 47548 38669 47564
rect 37886 47470 37902 47504
rect 38078 47470 38094 47504
rect 38384 47470 38400 47504
rect 38576 47470 38592 47504
rect 38635 47498 38669 47514
rect 37730 47400 37760 47452
rect 37670 47340 37760 47400
rect 37670 47100 37690 47340
rect 37730 47300 37760 47340
rect 37750 47142 37760 47300
rect 38730 47452 38738 47610
rect 38730 47420 38760 47452
rect 38800 47420 38820 47660
rect 38730 47340 38820 47420
rect 38730 47300 38760 47340
rect 37818 47238 37852 47254
rect 37886 47248 37902 47282
rect 38078 47248 38094 47282
rect 38384 47248 38400 47282
rect 38576 47248 38592 47282
rect 37818 47188 37852 47204
rect 38635 47238 38669 47254
rect 37886 47160 37902 47194
rect 38078 47160 38094 47194
rect 38384 47160 38400 47194
rect 38576 47160 38592 47194
rect 38635 47188 38669 47204
rect 37730 47100 37760 47142
rect 37670 46970 37760 47100
rect 38730 47142 38738 47300
rect 38730 47100 38760 47142
rect 38800 47100 38820 47340
rect 38730 46970 38820 47100
rect 42660 47660 42750 47780
rect 42660 47400 42680 47660
rect 42720 47610 42750 47660
rect 42740 47452 42750 47610
rect 43720 47660 43810 47780
rect 43720 47610 43750 47660
rect 42808 47548 42842 47564
rect 42876 47558 42892 47592
rect 43068 47558 43084 47592
rect 43374 47558 43390 47592
rect 43566 47558 43582 47592
rect 42808 47498 42842 47514
rect 43625 47548 43659 47564
rect 42876 47470 42892 47504
rect 43068 47470 43084 47504
rect 43374 47470 43390 47504
rect 43566 47470 43582 47504
rect 43625 47498 43659 47514
rect 42720 47400 42750 47452
rect 42660 47340 42750 47400
rect 42660 47100 42680 47340
rect 42720 47300 42750 47340
rect 42740 47142 42750 47300
rect 43720 47452 43728 47610
rect 43720 47420 43750 47452
rect 43790 47420 43810 47660
rect 43720 47340 43810 47420
rect 43720 47300 43750 47340
rect 42808 47238 42842 47254
rect 42876 47248 42892 47282
rect 43068 47248 43084 47282
rect 43374 47248 43390 47282
rect 43566 47248 43582 47282
rect 42808 47188 42842 47204
rect 43625 47238 43659 47254
rect 42876 47160 42892 47194
rect 43068 47160 43084 47194
rect 43374 47160 43390 47194
rect 43566 47160 43582 47194
rect 43625 47188 43659 47204
rect 42720 47100 42750 47142
rect 42660 46970 42750 47100
rect 43720 47142 43728 47300
rect 43720 47100 43750 47142
rect 43790 47100 43810 47340
rect 43720 46970 43810 47100
rect 47650 47660 47740 47780
rect 47650 47400 47670 47660
rect 47710 47610 47740 47660
rect 47730 47452 47740 47610
rect 48710 47660 48800 47780
rect 48710 47610 48740 47660
rect 47798 47548 47832 47564
rect 47866 47558 47882 47592
rect 48058 47558 48074 47592
rect 48364 47558 48380 47592
rect 48556 47558 48572 47592
rect 47798 47498 47832 47514
rect 48615 47548 48649 47564
rect 47866 47470 47882 47504
rect 48058 47470 48074 47504
rect 48364 47470 48380 47504
rect 48556 47470 48572 47504
rect 48615 47498 48649 47514
rect 47710 47400 47740 47452
rect 47650 47340 47740 47400
rect 47650 47100 47670 47340
rect 47710 47300 47740 47340
rect 47730 47142 47740 47300
rect 48710 47452 48718 47610
rect 48710 47420 48740 47452
rect 48780 47420 48800 47660
rect 48710 47340 48800 47420
rect 48710 47300 48740 47340
rect 47798 47238 47832 47254
rect 47866 47248 47882 47282
rect 48058 47248 48074 47282
rect 48364 47248 48380 47282
rect 48556 47248 48572 47282
rect 47798 47188 47832 47204
rect 48615 47238 48649 47254
rect 47866 47160 47882 47194
rect 48058 47160 48074 47194
rect 48364 47160 48380 47194
rect 48556 47160 48572 47194
rect 48615 47188 48649 47204
rect 47710 47100 47740 47142
rect 47650 46970 47740 47100
rect 48710 47142 48718 47300
rect 48710 47100 48740 47142
rect 48780 47100 48800 47340
rect 48710 46970 48800 47100
rect 52640 47660 52730 47780
rect 52640 47400 52660 47660
rect 52700 47610 52730 47660
rect 52720 47452 52730 47610
rect 53700 47660 53790 47780
rect 53700 47610 53730 47660
rect 52788 47548 52822 47564
rect 52856 47558 52872 47592
rect 53048 47558 53064 47592
rect 53354 47558 53370 47592
rect 53546 47558 53562 47592
rect 52788 47498 52822 47514
rect 53605 47548 53639 47564
rect 52856 47470 52872 47504
rect 53048 47470 53064 47504
rect 53354 47470 53370 47504
rect 53546 47470 53562 47504
rect 53605 47498 53639 47514
rect 52700 47400 52730 47452
rect 52640 47340 52730 47400
rect 52640 47100 52660 47340
rect 52700 47300 52730 47340
rect 52720 47142 52730 47300
rect 53700 47452 53708 47610
rect 53700 47420 53730 47452
rect 53770 47420 53790 47660
rect 53700 47340 53790 47420
rect 53700 47300 53730 47340
rect 52788 47238 52822 47254
rect 52856 47248 52872 47282
rect 53048 47248 53064 47282
rect 53354 47248 53370 47282
rect 53546 47248 53562 47282
rect 52788 47188 52822 47204
rect 53605 47238 53639 47254
rect 52856 47160 52872 47194
rect 53048 47160 53064 47194
rect 53354 47160 53370 47194
rect 53546 47160 53562 47194
rect 53605 47188 53639 47204
rect 52700 47100 52730 47142
rect 52640 46970 52730 47100
rect 53700 47142 53708 47300
rect 53700 47100 53730 47142
rect 53770 47100 53790 47340
rect 53700 46970 53790 47100
rect 57630 47660 57720 47780
rect 57630 47400 57650 47660
rect 57690 47610 57720 47660
rect 57710 47452 57720 47610
rect 58690 47660 58780 47780
rect 58690 47610 58720 47660
rect 57778 47548 57812 47564
rect 57846 47558 57862 47592
rect 58038 47558 58054 47592
rect 58344 47558 58360 47592
rect 58536 47558 58552 47592
rect 57778 47498 57812 47514
rect 58595 47548 58629 47564
rect 57846 47470 57862 47504
rect 58038 47470 58054 47504
rect 58344 47470 58360 47504
rect 58536 47470 58552 47504
rect 58595 47498 58629 47514
rect 57690 47400 57720 47452
rect 57630 47340 57720 47400
rect 57630 47100 57650 47340
rect 57690 47300 57720 47340
rect 57710 47142 57720 47300
rect 58690 47452 58698 47610
rect 58690 47420 58720 47452
rect 58760 47420 58780 47660
rect 58690 47340 58780 47420
rect 58690 47300 58720 47340
rect 57778 47238 57812 47254
rect 57846 47248 57862 47282
rect 58038 47248 58054 47282
rect 58344 47248 58360 47282
rect 58536 47248 58552 47282
rect 57778 47188 57812 47204
rect 58595 47238 58629 47254
rect 57846 47160 57862 47194
rect 58038 47160 58054 47194
rect 58344 47160 58360 47194
rect 58536 47160 58552 47194
rect 58595 47188 58629 47204
rect 57690 47100 57720 47142
rect 57630 46970 57720 47100
rect 58690 47142 58698 47300
rect 58690 47100 58720 47142
rect 58760 47100 58780 47340
rect 58690 46970 58780 47100
rect 62620 47660 62710 47780
rect 62620 47400 62640 47660
rect 62680 47610 62710 47660
rect 62700 47452 62710 47610
rect 63680 47660 63770 47780
rect 63680 47610 63710 47660
rect 62768 47548 62802 47564
rect 62836 47558 62852 47592
rect 63028 47558 63044 47592
rect 63334 47558 63350 47592
rect 63526 47558 63542 47592
rect 62768 47498 62802 47514
rect 63585 47548 63619 47564
rect 62836 47470 62852 47504
rect 63028 47470 63044 47504
rect 63334 47470 63350 47504
rect 63526 47470 63542 47504
rect 63585 47498 63619 47514
rect 62680 47400 62710 47452
rect 62620 47340 62710 47400
rect 62620 47100 62640 47340
rect 62680 47300 62710 47340
rect 62700 47142 62710 47300
rect 63680 47452 63688 47610
rect 63680 47420 63710 47452
rect 63750 47420 63770 47660
rect 63680 47340 63770 47420
rect 63680 47300 63710 47340
rect 62768 47238 62802 47254
rect 62836 47248 62852 47282
rect 63028 47248 63044 47282
rect 63334 47248 63350 47282
rect 63526 47248 63542 47282
rect 62768 47188 62802 47204
rect 63585 47238 63619 47254
rect 62836 47160 62852 47194
rect 63028 47160 63044 47194
rect 63334 47160 63350 47194
rect 63526 47160 63542 47194
rect 63585 47188 63619 47204
rect 62680 47100 62710 47142
rect 62620 46970 62710 47100
rect 63680 47142 63688 47300
rect 63680 47100 63710 47142
rect 63750 47100 63770 47340
rect 63680 46970 63770 47100
rect 67610 47660 67700 47780
rect 67610 47400 67630 47660
rect 67670 47610 67700 47660
rect 67690 47452 67700 47610
rect 68670 47660 68760 47780
rect 68670 47610 68700 47660
rect 67758 47548 67792 47564
rect 67826 47558 67842 47592
rect 68018 47558 68034 47592
rect 68324 47558 68340 47592
rect 68516 47558 68532 47592
rect 67758 47498 67792 47514
rect 68575 47548 68609 47564
rect 67826 47470 67842 47504
rect 68018 47470 68034 47504
rect 68324 47470 68340 47504
rect 68516 47470 68532 47504
rect 68575 47498 68609 47514
rect 67670 47400 67700 47452
rect 67610 47340 67700 47400
rect 67610 47100 67630 47340
rect 67670 47300 67700 47340
rect 67690 47142 67700 47300
rect 68670 47452 68678 47610
rect 68670 47420 68700 47452
rect 68740 47420 68760 47660
rect 68670 47340 68760 47420
rect 68670 47300 68700 47340
rect 67758 47238 67792 47254
rect 67826 47248 67842 47282
rect 68018 47248 68034 47282
rect 68324 47248 68340 47282
rect 68516 47248 68532 47282
rect 67758 47188 67792 47204
rect 68575 47238 68609 47254
rect 67826 47160 67842 47194
rect 68018 47160 68034 47194
rect 68324 47160 68340 47194
rect 68516 47160 68532 47194
rect 68575 47188 68609 47204
rect 67670 47100 67700 47142
rect 67610 46970 67700 47100
rect 68670 47142 68678 47300
rect 68670 47100 68700 47142
rect 68740 47100 68760 47340
rect 68670 46970 68760 47100
rect 72600 47660 72690 47780
rect 72600 47400 72620 47660
rect 72660 47610 72690 47660
rect 72680 47452 72690 47610
rect 73660 47660 73750 47780
rect 73660 47610 73690 47660
rect 72748 47548 72782 47564
rect 72816 47558 72832 47592
rect 73008 47558 73024 47592
rect 73314 47558 73330 47592
rect 73506 47558 73522 47592
rect 72748 47498 72782 47514
rect 73565 47548 73599 47564
rect 72816 47470 72832 47504
rect 73008 47470 73024 47504
rect 73314 47470 73330 47504
rect 73506 47470 73522 47504
rect 73565 47498 73599 47514
rect 72660 47400 72690 47452
rect 72600 47340 72690 47400
rect 72600 47100 72620 47340
rect 72660 47300 72690 47340
rect 72680 47142 72690 47300
rect 73660 47452 73668 47610
rect 73660 47420 73690 47452
rect 73730 47420 73750 47660
rect 73660 47340 73750 47420
rect 73660 47300 73690 47340
rect 72748 47238 72782 47254
rect 72816 47248 72832 47282
rect 73008 47248 73024 47282
rect 73314 47248 73330 47282
rect 73506 47248 73522 47282
rect 72748 47188 72782 47204
rect 73565 47238 73599 47254
rect 72816 47160 72832 47194
rect 73008 47160 73024 47194
rect 73314 47160 73330 47194
rect 73506 47160 73522 47194
rect 73565 47188 73599 47204
rect 72660 47100 72690 47142
rect 72600 46970 72690 47100
rect 73660 47142 73668 47300
rect 73660 47100 73690 47142
rect 73730 47100 73750 47340
rect 73660 46970 73750 47100
rect 77590 47660 77680 47780
rect 77590 47400 77610 47660
rect 77650 47610 77680 47660
rect 77670 47452 77680 47610
rect 78650 47660 78740 47780
rect 78650 47610 78680 47660
rect 77738 47548 77772 47564
rect 77806 47558 77822 47592
rect 77998 47558 78014 47592
rect 78304 47558 78320 47592
rect 78496 47558 78512 47592
rect 77738 47498 77772 47514
rect 78555 47548 78589 47564
rect 77806 47470 77822 47504
rect 77998 47470 78014 47504
rect 78304 47470 78320 47504
rect 78496 47470 78512 47504
rect 78555 47498 78589 47514
rect 77650 47400 77680 47452
rect 77590 47340 77680 47400
rect 77590 47100 77610 47340
rect 77650 47300 77680 47340
rect 77670 47142 77680 47300
rect 78650 47452 78658 47610
rect 78650 47420 78680 47452
rect 78720 47420 78740 47660
rect 78650 47340 78740 47420
rect 78650 47300 78680 47340
rect 77738 47238 77772 47254
rect 77806 47248 77822 47282
rect 77998 47248 78014 47282
rect 78304 47248 78320 47282
rect 78496 47248 78512 47282
rect 77738 47188 77772 47204
rect 78555 47238 78589 47254
rect 77806 47160 77822 47194
rect 77998 47160 78014 47194
rect 78304 47160 78320 47194
rect 78496 47160 78512 47194
rect 78555 47188 78589 47204
rect 77650 47100 77680 47142
rect 77590 46970 77680 47100
rect 78650 47142 78658 47300
rect 78650 47100 78680 47142
rect 78720 47100 78740 47340
rect 78650 46970 78740 47100
rect 2740 45950 2830 46070
rect 2740 45690 2760 45950
rect 2800 45900 2830 45950
rect 2820 45742 2830 45900
rect 3800 45950 3890 46070
rect 3800 45900 3830 45950
rect 2888 45838 2922 45854
rect 2956 45848 2972 45882
rect 3148 45848 3164 45882
rect 3454 45848 3470 45882
rect 3646 45848 3662 45882
rect 2888 45788 2922 45804
rect 3705 45838 3739 45854
rect 2956 45760 2972 45794
rect 3148 45760 3164 45794
rect 3454 45760 3470 45794
rect 3646 45760 3662 45794
rect 3705 45788 3739 45804
rect 2800 45690 2830 45742
rect 2740 45630 2830 45690
rect 2740 45390 2760 45630
rect 2800 45590 2830 45630
rect 2820 45432 2830 45590
rect 3800 45742 3808 45900
rect 3800 45710 3830 45742
rect 3870 45710 3890 45950
rect 3800 45630 3890 45710
rect 3800 45590 3830 45630
rect 2888 45528 2922 45544
rect 2956 45538 2972 45572
rect 3148 45538 3164 45572
rect 3454 45538 3470 45572
rect 3646 45538 3662 45572
rect 2888 45478 2922 45494
rect 3705 45528 3739 45544
rect 2956 45450 2972 45484
rect 3148 45450 3164 45484
rect 3454 45450 3470 45484
rect 3646 45450 3662 45484
rect 3705 45478 3739 45494
rect 2800 45390 2830 45432
rect 2740 45260 2830 45390
rect 3800 45432 3808 45590
rect 3800 45390 3830 45432
rect 3870 45390 3890 45630
rect 3800 45260 3890 45390
rect 7730 45950 7820 46070
rect 7730 45690 7750 45950
rect 7790 45900 7820 45950
rect 7810 45742 7820 45900
rect 8790 45950 8880 46070
rect 8790 45900 8820 45950
rect 7878 45838 7912 45854
rect 7946 45848 7962 45882
rect 8138 45848 8154 45882
rect 8444 45848 8460 45882
rect 8636 45848 8652 45882
rect 7878 45788 7912 45804
rect 8695 45838 8729 45854
rect 7946 45760 7962 45794
rect 8138 45760 8154 45794
rect 8444 45760 8460 45794
rect 8636 45760 8652 45794
rect 8695 45788 8729 45804
rect 7790 45690 7820 45742
rect 7730 45630 7820 45690
rect 7730 45390 7750 45630
rect 7790 45590 7820 45630
rect 7810 45432 7820 45590
rect 8790 45742 8798 45900
rect 8790 45710 8820 45742
rect 8860 45710 8880 45950
rect 8790 45630 8880 45710
rect 8790 45590 8820 45630
rect 7878 45528 7912 45544
rect 7946 45538 7962 45572
rect 8138 45538 8154 45572
rect 8444 45538 8460 45572
rect 8636 45538 8652 45572
rect 7878 45478 7912 45494
rect 8695 45528 8729 45544
rect 7946 45450 7962 45484
rect 8138 45450 8154 45484
rect 8444 45450 8460 45484
rect 8636 45450 8652 45484
rect 8695 45478 8729 45494
rect 7790 45390 7820 45432
rect 7730 45260 7820 45390
rect 8790 45432 8798 45590
rect 8790 45390 8820 45432
rect 8860 45390 8880 45630
rect 8790 45260 8880 45390
rect 12720 45950 12810 46070
rect 12720 45690 12740 45950
rect 12780 45900 12810 45950
rect 12800 45742 12810 45900
rect 13780 45950 13870 46070
rect 13780 45900 13810 45950
rect 12868 45838 12902 45854
rect 12936 45848 12952 45882
rect 13128 45848 13144 45882
rect 13434 45848 13450 45882
rect 13626 45848 13642 45882
rect 12868 45788 12902 45804
rect 13685 45838 13719 45854
rect 12936 45760 12952 45794
rect 13128 45760 13144 45794
rect 13434 45760 13450 45794
rect 13626 45760 13642 45794
rect 13685 45788 13719 45804
rect 12780 45690 12810 45742
rect 12720 45630 12810 45690
rect 12720 45390 12740 45630
rect 12780 45590 12810 45630
rect 12800 45432 12810 45590
rect 13780 45742 13788 45900
rect 13780 45710 13810 45742
rect 13850 45710 13870 45950
rect 13780 45630 13870 45710
rect 13780 45590 13810 45630
rect 12868 45528 12902 45544
rect 12936 45538 12952 45572
rect 13128 45538 13144 45572
rect 13434 45538 13450 45572
rect 13626 45538 13642 45572
rect 12868 45478 12902 45494
rect 13685 45528 13719 45544
rect 12936 45450 12952 45484
rect 13128 45450 13144 45484
rect 13434 45450 13450 45484
rect 13626 45450 13642 45484
rect 13685 45478 13719 45494
rect 12780 45390 12810 45432
rect 12720 45260 12810 45390
rect 13780 45432 13788 45590
rect 13780 45390 13810 45432
rect 13850 45390 13870 45630
rect 13780 45260 13870 45390
rect 17710 45950 17800 46070
rect 17710 45690 17730 45950
rect 17770 45900 17800 45950
rect 17790 45742 17800 45900
rect 18770 45950 18860 46070
rect 18770 45900 18800 45950
rect 17858 45838 17892 45854
rect 17926 45848 17942 45882
rect 18118 45848 18134 45882
rect 18424 45848 18440 45882
rect 18616 45848 18632 45882
rect 17858 45788 17892 45804
rect 18675 45838 18709 45854
rect 17926 45760 17942 45794
rect 18118 45760 18134 45794
rect 18424 45760 18440 45794
rect 18616 45760 18632 45794
rect 18675 45788 18709 45804
rect 17770 45690 17800 45742
rect 17710 45630 17800 45690
rect 17710 45390 17730 45630
rect 17770 45590 17800 45630
rect 17790 45432 17800 45590
rect 18770 45742 18778 45900
rect 18770 45710 18800 45742
rect 18840 45710 18860 45950
rect 18770 45630 18860 45710
rect 18770 45590 18800 45630
rect 17858 45528 17892 45544
rect 17926 45538 17942 45572
rect 18118 45538 18134 45572
rect 18424 45538 18440 45572
rect 18616 45538 18632 45572
rect 17858 45478 17892 45494
rect 18675 45528 18709 45544
rect 17926 45450 17942 45484
rect 18118 45450 18134 45484
rect 18424 45450 18440 45484
rect 18616 45450 18632 45484
rect 18675 45478 18709 45494
rect 17770 45390 17800 45432
rect 17710 45260 17800 45390
rect 18770 45432 18778 45590
rect 18770 45390 18800 45432
rect 18840 45390 18860 45630
rect 18770 45260 18860 45390
rect 22700 45950 22790 46070
rect 22700 45690 22720 45950
rect 22760 45900 22790 45950
rect 22780 45742 22790 45900
rect 23760 45950 23850 46070
rect 23760 45900 23790 45950
rect 22848 45838 22882 45854
rect 22916 45848 22932 45882
rect 23108 45848 23124 45882
rect 23414 45848 23430 45882
rect 23606 45848 23622 45882
rect 22848 45788 22882 45804
rect 23665 45838 23699 45854
rect 22916 45760 22932 45794
rect 23108 45760 23124 45794
rect 23414 45760 23430 45794
rect 23606 45760 23622 45794
rect 23665 45788 23699 45804
rect 22760 45690 22790 45742
rect 22700 45630 22790 45690
rect 22700 45390 22720 45630
rect 22760 45590 22790 45630
rect 22780 45432 22790 45590
rect 23760 45742 23768 45900
rect 23760 45710 23790 45742
rect 23830 45710 23850 45950
rect 23760 45630 23850 45710
rect 23760 45590 23790 45630
rect 22848 45528 22882 45544
rect 22916 45538 22932 45572
rect 23108 45538 23124 45572
rect 23414 45538 23430 45572
rect 23606 45538 23622 45572
rect 22848 45478 22882 45494
rect 23665 45528 23699 45544
rect 22916 45450 22932 45484
rect 23108 45450 23124 45484
rect 23414 45450 23430 45484
rect 23606 45450 23622 45484
rect 23665 45478 23699 45494
rect 22760 45390 22790 45432
rect 22700 45260 22790 45390
rect 23760 45432 23768 45590
rect 23760 45390 23790 45432
rect 23830 45390 23850 45630
rect 23760 45260 23850 45390
rect 27690 45950 27780 46070
rect 27690 45690 27710 45950
rect 27750 45900 27780 45950
rect 27770 45742 27780 45900
rect 28750 45950 28840 46070
rect 28750 45900 28780 45950
rect 27838 45838 27872 45854
rect 27906 45848 27922 45882
rect 28098 45848 28114 45882
rect 28404 45848 28420 45882
rect 28596 45848 28612 45882
rect 27838 45788 27872 45804
rect 28655 45838 28689 45854
rect 27906 45760 27922 45794
rect 28098 45760 28114 45794
rect 28404 45760 28420 45794
rect 28596 45760 28612 45794
rect 28655 45788 28689 45804
rect 27750 45690 27780 45742
rect 27690 45630 27780 45690
rect 27690 45390 27710 45630
rect 27750 45590 27780 45630
rect 27770 45432 27780 45590
rect 28750 45742 28758 45900
rect 28750 45710 28780 45742
rect 28820 45710 28840 45950
rect 28750 45630 28840 45710
rect 28750 45590 28780 45630
rect 27838 45528 27872 45544
rect 27906 45538 27922 45572
rect 28098 45538 28114 45572
rect 28404 45538 28420 45572
rect 28596 45538 28612 45572
rect 27838 45478 27872 45494
rect 28655 45528 28689 45544
rect 27906 45450 27922 45484
rect 28098 45450 28114 45484
rect 28404 45450 28420 45484
rect 28596 45450 28612 45484
rect 28655 45478 28689 45494
rect 27750 45390 27780 45432
rect 27690 45260 27780 45390
rect 28750 45432 28758 45590
rect 28750 45390 28780 45432
rect 28820 45390 28840 45630
rect 28750 45260 28840 45390
rect 32680 45950 32770 46070
rect 32680 45690 32700 45950
rect 32740 45900 32770 45950
rect 32760 45742 32770 45900
rect 33740 45950 33830 46070
rect 33740 45900 33770 45950
rect 32828 45838 32862 45854
rect 32896 45848 32912 45882
rect 33088 45848 33104 45882
rect 33394 45848 33410 45882
rect 33586 45848 33602 45882
rect 32828 45788 32862 45804
rect 33645 45838 33679 45854
rect 32896 45760 32912 45794
rect 33088 45760 33104 45794
rect 33394 45760 33410 45794
rect 33586 45760 33602 45794
rect 33645 45788 33679 45804
rect 32740 45690 32770 45742
rect 32680 45630 32770 45690
rect 32680 45390 32700 45630
rect 32740 45590 32770 45630
rect 32760 45432 32770 45590
rect 33740 45742 33748 45900
rect 33740 45710 33770 45742
rect 33810 45710 33830 45950
rect 33740 45630 33830 45710
rect 33740 45590 33770 45630
rect 32828 45528 32862 45544
rect 32896 45538 32912 45572
rect 33088 45538 33104 45572
rect 33394 45538 33410 45572
rect 33586 45538 33602 45572
rect 32828 45478 32862 45494
rect 33645 45528 33679 45544
rect 32896 45450 32912 45484
rect 33088 45450 33104 45484
rect 33394 45450 33410 45484
rect 33586 45450 33602 45484
rect 33645 45478 33679 45494
rect 32740 45390 32770 45432
rect 32680 45260 32770 45390
rect 33740 45432 33748 45590
rect 33740 45390 33770 45432
rect 33810 45390 33830 45630
rect 33740 45260 33830 45390
rect 37670 45950 37760 46070
rect 37670 45690 37690 45950
rect 37730 45900 37760 45950
rect 37750 45742 37760 45900
rect 38730 45950 38820 46070
rect 38730 45900 38760 45950
rect 37818 45838 37852 45854
rect 37886 45848 37902 45882
rect 38078 45848 38094 45882
rect 38384 45848 38400 45882
rect 38576 45848 38592 45882
rect 37818 45788 37852 45804
rect 38635 45838 38669 45854
rect 37886 45760 37902 45794
rect 38078 45760 38094 45794
rect 38384 45760 38400 45794
rect 38576 45760 38592 45794
rect 38635 45788 38669 45804
rect 37730 45690 37760 45742
rect 37670 45630 37760 45690
rect 37670 45390 37690 45630
rect 37730 45590 37760 45630
rect 37750 45432 37760 45590
rect 38730 45742 38738 45900
rect 38730 45710 38760 45742
rect 38800 45710 38820 45950
rect 38730 45630 38820 45710
rect 38730 45590 38760 45630
rect 37818 45528 37852 45544
rect 37886 45538 37902 45572
rect 38078 45538 38094 45572
rect 38384 45538 38400 45572
rect 38576 45538 38592 45572
rect 37818 45478 37852 45494
rect 38635 45528 38669 45544
rect 37886 45450 37902 45484
rect 38078 45450 38094 45484
rect 38384 45450 38400 45484
rect 38576 45450 38592 45484
rect 38635 45478 38669 45494
rect 37730 45390 37760 45432
rect 37670 45260 37760 45390
rect 38730 45432 38738 45590
rect 38730 45390 38760 45432
rect 38800 45390 38820 45630
rect 38730 45260 38820 45390
rect 42660 45950 42750 46070
rect 42660 45690 42680 45950
rect 42720 45900 42750 45950
rect 42740 45742 42750 45900
rect 43720 45950 43810 46070
rect 43720 45900 43750 45950
rect 42808 45838 42842 45854
rect 42876 45848 42892 45882
rect 43068 45848 43084 45882
rect 43374 45848 43390 45882
rect 43566 45848 43582 45882
rect 42808 45788 42842 45804
rect 43625 45838 43659 45854
rect 42876 45760 42892 45794
rect 43068 45760 43084 45794
rect 43374 45760 43390 45794
rect 43566 45760 43582 45794
rect 43625 45788 43659 45804
rect 42720 45690 42750 45742
rect 42660 45630 42750 45690
rect 42660 45390 42680 45630
rect 42720 45590 42750 45630
rect 42740 45432 42750 45590
rect 43720 45742 43728 45900
rect 43720 45710 43750 45742
rect 43790 45710 43810 45950
rect 43720 45630 43810 45710
rect 43720 45590 43750 45630
rect 42808 45528 42842 45544
rect 42876 45538 42892 45572
rect 43068 45538 43084 45572
rect 43374 45538 43390 45572
rect 43566 45538 43582 45572
rect 42808 45478 42842 45494
rect 43625 45528 43659 45544
rect 42876 45450 42892 45484
rect 43068 45450 43084 45484
rect 43374 45450 43390 45484
rect 43566 45450 43582 45484
rect 43625 45478 43659 45494
rect 42720 45390 42750 45432
rect 42660 45260 42750 45390
rect 43720 45432 43728 45590
rect 43720 45390 43750 45432
rect 43790 45390 43810 45630
rect 43720 45260 43810 45390
rect 47650 45950 47740 46070
rect 47650 45690 47670 45950
rect 47710 45900 47740 45950
rect 47730 45742 47740 45900
rect 48710 45950 48800 46070
rect 48710 45900 48740 45950
rect 47798 45838 47832 45854
rect 47866 45848 47882 45882
rect 48058 45848 48074 45882
rect 48364 45848 48380 45882
rect 48556 45848 48572 45882
rect 47798 45788 47832 45804
rect 48615 45838 48649 45854
rect 47866 45760 47882 45794
rect 48058 45760 48074 45794
rect 48364 45760 48380 45794
rect 48556 45760 48572 45794
rect 48615 45788 48649 45804
rect 47710 45690 47740 45742
rect 47650 45630 47740 45690
rect 47650 45390 47670 45630
rect 47710 45590 47740 45630
rect 47730 45432 47740 45590
rect 48710 45742 48718 45900
rect 48710 45710 48740 45742
rect 48780 45710 48800 45950
rect 48710 45630 48800 45710
rect 48710 45590 48740 45630
rect 47798 45528 47832 45544
rect 47866 45538 47882 45572
rect 48058 45538 48074 45572
rect 48364 45538 48380 45572
rect 48556 45538 48572 45572
rect 47798 45478 47832 45494
rect 48615 45528 48649 45544
rect 47866 45450 47882 45484
rect 48058 45450 48074 45484
rect 48364 45450 48380 45484
rect 48556 45450 48572 45484
rect 48615 45478 48649 45494
rect 47710 45390 47740 45432
rect 47650 45260 47740 45390
rect 48710 45432 48718 45590
rect 48710 45390 48740 45432
rect 48780 45390 48800 45630
rect 48710 45260 48800 45390
rect 52640 45950 52730 46070
rect 52640 45690 52660 45950
rect 52700 45900 52730 45950
rect 52720 45742 52730 45900
rect 53700 45950 53790 46070
rect 53700 45900 53730 45950
rect 52788 45838 52822 45854
rect 52856 45848 52872 45882
rect 53048 45848 53064 45882
rect 53354 45848 53370 45882
rect 53546 45848 53562 45882
rect 52788 45788 52822 45804
rect 53605 45838 53639 45854
rect 52856 45760 52872 45794
rect 53048 45760 53064 45794
rect 53354 45760 53370 45794
rect 53546 45760 53562 45794
rect 53605 45788 53639 45804
rect 52700 45690 52730 45742
rect 52640 45630 52730 45690
rect 52640 45390 52660 45630
rect 52700 45590 52730 45630
rect 52720 45432 52730 45590
rect 53700 45742 53708 45900
rect 53700 45710 53730 45742
rect 53770 45710 53790 45950
rect 53700 45630 53790 45710
rect 53700 45590 53730 45630
rect 52788 45528 52822 45544
rect 52856 45538 52872 45572
rect 53048 45538 53064 45572
rect 53354 45538 53370 45572
rect 53546 45538 53562 45572
rect 52788 45478 52822 45494
rect 53605 45528 53639 45544
rect 52856 45450 52872 45484
rect 53048 45450 53064 45484
rect 53354 45450 53370 45484
rect 53546 45450 53562 45484
rect 53605 45478 53639 45494
rect 52700 45390 52730 45432
rect 52640 45260 52730 45390
rect 53700 45432 53708 45590
rect 53700 45390 53730 45432
rect 53770 45390 53790 45630
rect 53700 45260 53790 45390
rect 57630 45950 57720 46070
rect 57630 45690 57650 45950
rect 57690 45900 57720 45950
rect 57710 45742 57720 45900
rect 58690 45950 58780 46070
rect 58690 45900 58720 45950
rect 57778 45838 57812 45854
rect 57846 45848 57862 45882
rect 58038 45848 58054 45882
rect 58344 45848 58360 45882
rect 58536 45848 58552 45882
rect 57778 45788 57812 45804
rect 58595 45838 58629 45854
rect 57846 45760 57862 45794
rect 58038 45760 58054 45794
rect 58344 45760 58360 45794
rect 58536 45760 58552 45794
rect 58595 45788 58629 45804
rect 57690 45690 57720 45742
rect 57630 45630 57720 45690
rect 57630 45390 57650 45630
rect 57690 45590 57720 45630
rect 57710 45432 57720 45590
rect 58690 45742 58698 45900
rect 58690 45710 58720 45742
rect 58760 45710 58780 45950
rect 58690 45630 58780 45710
rect 58690 45590 58720 45630
rect 57778 45528 57812 45544
rect 57846 45538 57862 45572
rect 58038 45538 58054 45572
rect 58344 45538 58360 45572
rect 58536 45538 58552 45572
rect 57778 45478 57812 45494
rect 58595 45528 58629 45544
rect 57846 45450 57862 45484
rect 58038 45450 58054 45484
rect 58344 45450 58360 45484
rect 58536 45450 58552 45484
rect 58595 45478 58629 45494
rect 57690 45390 57720 45432
rect 57630 45260 57720 45390
rect 58690 45432 58698 45590
rect 58690 45390 58720 45432
rect 58760 45390 58780 45630
rect 58690 45260 58780 45390
rect 62620 45950 62710 46070
rect 62620 45690 62640 45950
rect 62680 45900 62710 45950
rect 62700 45742 62710 45900
rect 63680 45950 63770 46070
rect 63680 45900 63710 45950
rect 62768 45838 62802 45854
rect 62836 45848 62852 45882
rect 63028 45848 63044 45882
rect 63334 45848 63350 45882
rect 63526 45848 63542 45882
rect 62768 45788 62802 45804
rect 63585 45838 63619 45854
rect 62836 45760 62852 45794
rect 63028 45760 63044 45794
rect 63334 45760 63350 45794
rect 63526 45760 63542 45794
rect 63585 45788 63619 45804
rect 62680 45690 62710 45742
rect 62620 45630 62710 45690
rect 62620 45390 62640 45630
rect 62680 45590 62710 45630
rect 62700 45432 62710 45590
rect 63680 45742 63688 45900
rect 63680 45710 63710 45742
rect 63750 45710 63770 45950
rect 63680 45630 63770 45710
rect 63680 45590 63710 45630
rect 62768 45528 62802 45544
rect 62836 45538 62852 45572
rect 63028 45538 63044 45572
rect 63334 45538 63350 45572
rect 63526 45538 63542 45572
rect 62768 45478 62802 45494
rect 63585 45528 63619 45544
rect 62836 45450 62852 45484
rect 63028 45450 63044 45484
rect 63334 45450 63350 45484
rect 63526 45450 63542 45484
rect 63585 45478 63619 45494
rect 62680 45390 62710 45432
rect 62620 45260 62710 45390
rect 63680 45432 63688 45590
rect 63680 45390 63710 45432
rect 63750 45390 63770 45630
rect 63680 45260 63770 45390
rect 67610 45950 67700 46070
rect 67610 45690 67630 45950
rect 67670 45900 67700 45950
rect 67690 45742 67700 45900
rect 68670 45950 68760 46070
rect 68670 45900 68700 45950
rect 67758 45838 67792 45854
rect 67826 45848 67842 45882
rect 68018 45848 68034 45882
rect 68324 45848 68340 45882
rect 68516 45848 68532 45882
rect 67758 45788 67792 45804
rect 68575 45838 68609 45854
rect 67826 45760 67842 45794
rect 68018 45760 68034 45794
rect 68324 45760 68340 45794
rect 68516 45760 68532 45794
rect 68575 45788 68609 45804
rect 67670 45690 67700 45742
rect 67610 45630 67700 45690
rect 67610 45390 67630 45630
rect 67670 45590 67700 45630
rect 67690 45432 67700 45590
rect 68670 45742 68678 45900
rect 68670 45710 68700 45742
rect 68740 45710 68760 45950
rect 68670 45630 68760 45710
rect 68670 45590 68700 45630
rect 67758 45528 67792 45544
rect 67826 45538 67842 45572
rect 68018 45538 68034 45572
rect 68324 45538 68340 45572
rect 68516 45538 68532 45572
rect 67758 45478 67792 45494
rect 68575 45528 68609 45544
rect 67826 45450 67842 45484
rect 68018 45450 68034 45484
rect 68324 45450 68340 45484
rect 68516 45450 68532 45484
rect 68575 45478 68609 45494
rect 67670 45390 67700 45432
rect 67610 45260 67700 45390
rect 68670 45432 68678 45590
rect 68670 45390 68700 45432
rect 68740 45390 68760 45630
rect 68670 45260 68760 45390
rect 72600 45950 72690 46070
rect 72600 45690 72620 45950
rect 72660 45900 72690 45950
rect 72680 45742 72690 45900
rect 73660 45950 73750 46070
rect 73660 45900 73690 45950
rect 72748 45838 72782 45854
rect 72816 45848 72832 45882
rect 73008 45848 73024 45882
rect 73314 45848 73330 45882
rect 73506 45848 73522 45882
rect 72748 45788 72782 45804
rect 73565 45838 73599 45854
rect 72816 45760 72832 45794
rect 73008 45760 73024 45794
rect 73314 45760 73330 45794
rect 73506 45760 73522 45794
rect 73565 45788 73599 45804
rect 72660 45690 72690 45742
rect 72600 45630 72690 45690
rect 72600 45390 72620 45630
rect 72660 45590 72690 45630
rect 72680 45432 72690 45590
rect 73660 45742 73668 45900
rect 73660 45710 73690 45742
rect 73730 45710 73750 45950
rect 73660 45630 73750 45710
rect 73660 45590 73690 45630
rect 72748 45528 72782 45544
rect 72816 45538 72832 45572
rect 73008 45538 73024 45572
rect 73314 45538 73330 45572
rect 73506 45538 73522 45572
rect 72748 45478 72782 45494
rect 73565 45528 73599 45544
rect 72816 45450 72832 45484
rect 73008 45450 73024 45484
rect 73314 45450 73330 45484
rect 73506 45450 73522 45484
rect 73565 45478 73599 45494
rect 72660 45390 72690 45432
rect 72600 45260 72690 45390
rect 73660 45432 73668 45590
rect 73660 45390 73690 45432
rect 73730 45390 73750 45630
rect 73660 45260 73750 45390
rect 77590 45950 77680 46070
rect 77590 45690 77610 45950
rect 77650 45900 77680 45950
rect 77670 45742 77680 45900
rect 78650 45950 78740 46070
rect 78650 45900 78680 45950
rect 77738 45838 77772 45854
rect 77806 45848 77822 45882
rect 77998 45848 78014 45882
rect 78304 45848 78320 45882
rect 78496 45848 78512 45882
rect 77738 45788 77772 45804
rect 78555 45838 78589 45854
rect 77806 45760 77822 45794
rect 77998 45760 78014 45794
rect 78304 45760 78320 45794
rect 78496 45760 78512 45794
rect 78555 45788 78589 45804
rect 77650 45690 77680 45742
rect 77590 45630 77680 45690
rect 77590 45390 77610 45630
rect 77650 45590 77680 45630
rect 77670 45432 77680 45590
rect 78650 45742 78658 45900
rect 78650 45710 78680 45742
rect 78720 45710 78740 45950
rect 78650 45630 78740 45710
rect 78650 45590 78680 45630
rect 77738 45528 77772 45544
rect 77806 45538 77822 45572
rect 77998 45538 78014 45572
rect 78304 45538 78320 45572
rect 78496 45538 78512 45572
rect 77738 45478 77772 45494
rect 78555 45528 78589 45544
rect 77806 45450 77822 45484
rect 77998 45450 78014 45484
rect 78304 45450 78320 45484
rect 78496 45450 78512 45484
rect 78555 45478 78589 45494
rect 77650 45390 77680 45432
rect 77590 45260 77680 45390
rect 78650 45432 78658 45590
rect 78650 45390 78680 45432
rect 78720 45390 78740 45630
rect 78650 45260 78740 45390
rect 2740 44240 2830 44360
rect 2740 43980 2760 44240
rect 2800 44190 2830 44240
rect 2820 44032 2830 44190
rect 3800 44240 3890 44360
rect 3800 44190 3830 44240
rect 2888 44128 2922 44144
rect 2956 44138 2972 44172
rect 3148 44138 3164 44172
rect 3454 44138 3470 44172
rect 3646 44138 3662 44172
rect 2888 44078 2922 44094
rect 3705 44128 3739 44144
rect 2956 44050 2972 44084
rect 3148 44050 3164 44084
rect 3454 44050 3470 44084
rect 3646 44050 3662 44084
rect 3705 44078 3739 44094
rect 2800 43980 2830 44032
rect 2740 43920 2830 43980
rect 2740 43680 2760 43920
rect 2800 43880 2830 43920
rect 2820 43722 2830 43880
rect 3800 44032 3808 44190
rect 3800 44000 3830 44032
rect 3870 44000 3890 44240
rect 3800 43920 3890 44000
rect 3800 43880 3830 43920
rect 2888 43818 2922 43834
rect 2956 43828 2972 43862
rect 3148 43828 3164 43862
rect 3454 43828 3470 43862
rect 3646 43828 3662 43862
rect 2888 43768 2922 43784
rect 3705 43818 3739 43834
rect 2956 43740 2972 43774
rect 3148 43740 3164 43774
rect 3454 43740 3470 43774
rect 3646 43740 3662 43774
rect 3705 43768 3739 43784
rect 2800 43680 2830 43722
rect 2740 43550 2830 43680
rect 3800 43722 3808 43880
rect 3800 43680 3830 43722
rect 3870 43680 3890 43920
rect 3800 43550 3890 43680
rect 7730 44240 7820 44360
rect 7730 43980 7750 44240
rect 7790 44190 7820 44240
rect 7810 44032 7820 44190
rect 8790 44240 8880 44360
rect 8790 44190 8820 44240
rect 7878 44128 7912 44144
rect 7946 44138 7962 44172
rect 8138 44138 8154 44172
rect 8444 44138 8460 44172
rect 8636 44138 8652 44172
rect 7878 44078 7912 44094
rect 8695 44128 8729 44144
rect 7946 44050 7962 44084
rect 8138 44050 8154 44084
rect 8444 44050 8460 44084
rect 8636 44050 8652 44084
rect 8695 44078 8729 44094
rect 7790 43980 7820 44032
rect 7730 43920 7820 43980
rect 7730 43680 7750 43920
rect 7790 43880 7820 43920
rect 7810 43722 7820 43880
rect 8790 44032 8798 44190
rect 8790 44000 8820 44032
rect 8860 44000 8880 44240
rect 8790 43920 8880 44000
rect 8790 43880 8820 43920
rect 7878 43818 7912 43834
rect 7946 43828 7962 43862
rect 8138 43828 8154 43862
rect 8444 43828 8460 43862
rect 8636 43828 8652 43862
rect 7878 43768 7912 43784
rect 8695 43818 8729 43834
rect 7946 43740 7962 43774
rect 8138 43740 8154 43774
rect 8444 43740 8460 43774
rect 8636 43740 8652 43774
rect 8695 43768 8729 43784
rect 7790 43680 7820 43722
rect 7730 43550 7820 43680
rect 8790 43722 8798 43880
rect 8790 43680 8820 43722
rect 8860 43680 8880 43920
rect 8790 43550 8880 43680
rect 12720 44240 12810 44360
rect 12720 43980 12740 44240
rect 12780 44190 12810 44240
rect 12800 44032 12810 44190
rect 13780 44240 13870 44360
rect 13780 44190 13810 44240
rect 12868 44128 12902 44144
rect 12936 44138 12952 44172
rect 13128 44138 13144 44172
rect 13434 44138 13450 44172
rect 13626 44138 13642 44172
rect 12868 44078 12902 44094
rect 13685 44128 13719 44144
rect 12936 44050 12952 44084
rect 13128 44050 13144 44084
rect 13434 44050 13450 44084
rect 13626 44050 13642 44084
rect 13685 44078 13719 44094
rect 12780 43980 12810 44032
rect 12720 43920 12810 43980
rect 12720 43680 12740 43920
rect 12780 43880 12810 43920
rect 12800 43722 12810 43880
rect 13780 44032 13788 44190
rect 13780 44000 13810 44032
rect 13850 44000 13870 44240
rect 13780 43920 13870 44000
rect 13780 43880 13810 43920
rect 12868 43818 12902 43834
rect 12936 43828 12952 43862
rect 13128 43828 13144 43862
rect 13434 43828 13450 43862
rect 13626 43828 13642 43862
rect 12868 43768 12902 43784
rect 13685 43818 13719 43834
rect 12936 43740 12952 43774
rect 13128 43740 13144 43774
rect 13434 43740 13450 43774
rect 13626 43740 13642 43774
rect 13685 43768 13719 43784
rect 12780 43680 12810 43722
rect 12720 43550 12810 43680
rect 13780 43722 13788 43880
rect 13780 43680 13810 43722
rect 13850 43680 13870 43920
rect 13780 43550 13870 43680
rect 17710 44240 17800 44360
rect 17710 43980 17730 44240
rect 17770 44190 17800 44240
rect 17790 44032 17800 44190
rect 18770 44240 18860 44360
rect 18770 44190 18800 44240
rect 17858 44128 17892 44144
rect 17926 44138 17942 44172
rect 18118 44138 18134 44172
rect 18424 44138 18440 44172
rect 18616 44138 18632 44172
rect 17858 44078 17892 44094
rect 18675 44128 18709 44144
rect 17926 44050 17942 44084
rect 18118 44050 18134 44084
rect 18424 44050 18440 44084
rect 18616 44050 18632 44084
rect 18675 44078 18709 44094
rect 17770 43980 17800 44032
rect 17710 43920 17800 43980
rect 17710 43680 17730 43920
rect 17770 43880 17800 43920
rect 17790 43722 17800 43880
rect 18770 44032 18778 44190
rect 18770 44000 18800 44032
rect 18840 44000 18860 44240
rect 18770 43920 18860 44000
rect 18770 43880 18800 43920
rect 17858 43818 17892 43834
rect 17926 43828 17942 43862
rect 18118 43828 18134 43862
rect 18424 43828 18440 43862
rect 18616 43828 18632 43862
rect 17858 43768 17892 43784
rect 18675 43818 18709 43834
rect 17926 43740 17942 43774
rect 18118 43740 18134 43774
rect 18424 43740 18440 43774
rect 18616 43740 18632 43774
rect 18675 43768 18709 43784
rect 17770 43680 17800 43722
rect 17710 43550 17800 43680
rect 18770 43722 18778 43880
rect 18770 43680 18800 43722
rect 18840 43680 18860 43920
rect 18770 43550 18860 43680
rect 22700 44240 22790 44360
rect 22700 43980 22720 44240
rect 22760 44190 22790 44240
rect 22780 44032 22790 44190
rect 23760 44240 23850 44360
rect 23760 44190 23790 44240
rect 22848 44128 22882 44144
rect 22916 44138 22932 44172
rect 23108 44138 23124 44172
rect 23414 44138 23430 44172
rect 23606 44138 23622 44172
rect 22848 44078 22882 44094
rect 23665 44128 23699 44144
rect 22916 44050 22932 44084
rect 23108 44050 23124 44084
rect 23414 44050 23430 44084
rect 23606 44050 23622 44084
rect 23665 44078 23699 44094
rect 22760 43980 22790 44032
rect 22700 43920 22790 43980
rect 22700 43680 22720 43920
rect 22760 43880 22790 43920
rect 22780 43722 22790 43880
rect 23760 44032 23768 44190
rect 23760 44000 23790 44032
rect 23830 44000 23850 44240
rect 23760 43920 23850 44000
rect 23760 43880 23790 43920
rect 22848 43818 22882 43834
rect 22916 43828 22932 43862
rect 23108 43828 23124 43862
rect 23414 43828 23430 43862
rect 23606 43828 23622 43862
rect 22848 43768 22882 43784
rect 23665 43818 23699 43834
rect 22916 43740 22932 43774
rect 23108 43740 23124 43774
rect 23414 43740 23430 43774
rect 23606 43740 23622 43774
rect 23665 43768 23699 43784
rect 22760 43680 22790 43722
rect 22700 43550 22790 43680
rect 23760 43722 23768 43880
rect 23760 43680 23790 43722
rect 23830 43680 23850 43920
rect 23760 43550 23850 43680
rect 27690 44240 27780 44360
rect 27690 43980 27710 44240
rect 27750 44190 27780 44240
rect 27770 44032 27780 44190
rect 28750 44240 28840 44360
rect 28750 44190 28780 44240
rect 27838 44128 27872 44144
rect 27906 44138 27922 44172
rect 28098 44138 28114 44172
rect 28404 44138 28420 44172
rect 28596 44138 28612 44172
rect 27838 44078 27872 44094
rect 28655 44128 28689 44144
rect 27906 44050 27922 44084
rect 28098 44050 28114 44084
rect 28404 44050 28420 44084
rect 28596 44050 28612 44084
rect 28655 44078 28689 44094
rect 27750 43980 27780 44032
rect 27690 43920 27780 43980
rect 27690 43680 27710 43920
rect 27750 43880 27780 43920
rect 27770 43722 27780 43880
rect 28750 44032 28758 44190
rect 28750 44000 28780 44032
rect 28820 44000 28840 44240
rect 28750 43920 28840 44000
rect 28750 43880 28780 43920
rect 27838 43818 27872 43834
rect 27906 43828 27922 43862
rect 28098 43828 28114 43862
rect 28404 43828 28420 43862
rect 28596 43828 28612 43862
rect 27838 43768 27872 43784
rect 28655 43818 28689 43834
rect 27906 43740 27922 43774
rect 28098 43740 28114 43774
rect 28404 43740 28420 43774
rect 28596 43740 28612 43774
rect 28655 43768 28689 43784
rect 27750 43680 27780 43722
rect 27690 43550 27780 43680
rect 28750 43722 28758 43880
rect 28750 43680 28780 43722
rect 28820 43680 28840 43920
rect 28750 43550 28840 43680
rect 32680 44240 32770 44360
rect 32680 43980 32700 44240
rect 32740 44190 32770 44240
rect 32760 44032 32770 44190
rect 33740 44240 33830 44360
rect 33740 44190 33770 44240
rect 32828 44128 32862 44144
rect 32896 44138 32912 44172
rect 33088 44138 33104 44172
rect 33394 44138 33410 44172
rect 33586 44138 33602 44172
rect 32828 44078 32862 44094
rect 33645 44128 33679 44144
rect 32896 44050 32912 44084
rect 33088 44050 33104 44084
rect 33394 44050 33410 44084
rect 33586 44050 33602 44084
rect 33645 44078 33679 44094
rect 32740 43980 32770 44032
rect 32680 43920 32770 43980
rect 32680 43680 32700 43920
rect 32740 43880 32770 43920
rect 32760 43722 32770 43880
rect 33740 44032 33748 44190
rect 33740 44000 33770 44032
rect 33810 44000 33830 44240
rect 33740 43920 33830 44000
rect 33740 43880 33770 43920
rect 32828 43818 32862 43834
rect 32896 43828 32912 43862
rect 33088 43828 33104 43862
rect 33394 43828 33410 43862
rect 33586 43828 33602 43862
rect 32828 43768 32862 43784
rect 33645 43818 33679 43834
rect 32896 43740 32912 43774
rect 33088 43740 33104 43774
rect 33394 43740 33410 43774
rect 33586 43740 33602 43774
rect 33645 43768 33679 43784
rect 32740 43680 32770 43722
rect 32680 43550 32770 43680
rect 33740 43722 33748 43880
rect 33740 43680 33770 43722
rect 33810 43680 33830 43920
rect 33740 43550 33830 43680
rect 37670 44240 37760 44360
rect 37670 43980 37690 44240
rect 37730 44190 37760 44240
rect 37750 44032 37760 44190
rect 38730 44240 38820 44360
rect 38730 44190 38760 44240
rect 37818 44128 37852 44144
rect 37886 44138 37902 44172
rect 38078 44138 38094 44172
rect 38384 44138 38400 44172
rect 38576 44138 38592 44172
rect 37818 44078 37852 44094
rect 38635 44128 38669 44144
rect 37886 44050 37902 44084
rect 38078 44050 38094 44084
rect 38384 44050 38400 44084
rect 38576 44050 38592 44084
rect 38635 44078 38669 44094
rect 37730 43980 37760 44032
rect 37670 43920 37760 43980
rect 37670 43680 37690 43920
rect 37730 43880 37760 43920
rect 37750 43722 37760 43880
rect 38730 44032 38738 44190
rect 38730 44000 38760 44032
rect 38800 44000 38820 44240
rect 38730 43920 38820 44000
rect 38730 43880 38760 43920
rect 37818 43818 37852 43834
rect 37886 43828 37902 43862
rect 38078 43828 38094 43862
rect 38384 43828 38400 43862
rect 38576 43828 38592 43862
rect 37818 43768 37852 43784
rect 38635 43818 38669 43834
rect 37886 43740 37902 43774
rect 38078 43740 38094 43774
rect 38384 43740 38400 43774
rect 38576 43740 38592 43774
rect 38635 43768 38669 43784
rect 37730 43680 37760 43722
rect 37670 43550 37760 43680
rect 38730 43722 38738 43880
rect 38730 43680 38760 43722
rect 38800 43680 38820 43920
rect 38730 43550 38820 43680
rect 42660 44240 42750 44360
rect 42660 43980 42680 44240
rect 42720 44190 42750 44240
rect 42740 44032 42750 44190
rect 43720 44240 43810 44360
rect 43720 44190 43750 44240
rect 42808 44128 42842 44144
rect 42876 44138 42892 44172
rect 43068 44138 43084 44172
rect 43374 44138 43390 44172
rect 43566 44138 43582 44172
rect 42808 44078 42842 44094
rect 43625 44128 43659 44144
rect 42876 44050 42892 44084
rect 43068 44050 43084 44084
rect 43374 44050 43390 44084
rect 43566 44050 43582 44084
rect 43625 44078 43659 44094
rect 42720 43980 42750 44032
rect 42660 43920 42750 43980
rect 42660 43680 42680 43920
rect 42720 43880 42750 43920
rect 42740 43722 42750 43880
rect 43720 44032 43728 44190
rect 43720 44000 43750 44032
rect 43790 44000 43810 44240
rect 43720 43920 43810 44000
rect 43720 43880 43750 43920
rect 42808 43818 42842 43834
rect 42876 43828 42892 43862
rect 43068 43828 43084 43862
rect 43374 43828 43390 43862
rect 43566 43828 43582 43862
rect 42808 43768 42842 43784
rect 43625 43818 43659 43834
rect 42876 43740 42892 43774
rect 43068 43740 43084 43774
rect 43374 43740 43390 43774
rect 43566 43740 43582 43774
rect 43625 43768 43659 43784
rect 42720 43680 42750 43722
rect 42660 43550 42750 43680
rect 43720 43722 43728 43880
rect 43720 43680 43750 43722
rect 43790 43680 43810 43920
rect 43720 43550 43810 43680
rect 47650 44240 47740 44360
rect 47650 43980 47670 44240
rect 47710 44190 47740 44240
rect 47730 44032 47740 44190
rect 48710 44240 48800 44360
rect 48710 44190 48740 44240
rect 47798 44128 47832 44144
rect 47866 44138 47882 44172
rect 48058 44138 48074 44172
rect 48364 44138 48380 44172
rect 48556 44138 48572 44172
rect 47798 44078 47832 44094
rect 48615 44128 48649 44144
rect 47866 44050 47882 44084
rect 48058 44050 48074 44084
rect 48364 44050 48380 44084
rect 48556 44050 48572 44084
rect 48615 44078 48649 44094
rect 47710 43980 47740 44032
rect 47650 43920 47740 43980
rect 47650 43680 47670 43920
rect 47710 43880 47740 43920
rect 47730 43722 47740 43880
rect 48710 44032 48718 44190
rect 48710 44000 48740 44032
rect 48780 44000 48800 44240
rect 48710 43920 48800 44000
rect 48710 43880 48740 43920
rect 47798 43818 47832 43834
rect 47866 43828 47882 43862
rect 48058 43828 48074 43862
rect 48364 43828 48380 43862
rect 48556 43828 48572 43862
rect 47798 43768 47832 43784
rect 48615 43818 48649 43834
rect 47866 43740 47882 43774
rect 48058 43740 48074 43774
rect 48364 43740 48380 43774
rect 48556 43740 48572 43774
rect 48615 43768 48649 43784
rect 47710 43680 47740 43722
rect 47650 43550 47740 43680
rect 48710 43722 48718 43880
rect 48710 43680 48740 43722
rect 48780 43680 48800 43920
rect 48710 43550 48800 43680
rect 52640 44240 52730 44360
rect 52640 43980 52660 44240
rect 52700 44190 52730 44240
rect 52720 44032 52730 44190
rect 53700 44240 53790 44360
rect 53700 44190 53730 44240
rect 52788 44128 52822 44144
rect 52856 44138 52872 44172
rect 53048 44138 53064 44172
rect 53354 44138 53370 44172
rect 53546 44138 53562 44172
rect 52788 44078 52822 44094
rect 53605 44128 53639 44144
rect 52856 44050 52872 44084
rect 53048 44050 53064 44084
rect 53354 44050 53370 44084
rect 53546 44050 53562 44084
rect 53605 44078 53639 44094
rect 52700 43980 52730 44032
rect 52640 43920 52730 43980
rect 52640 43680 52660 43920
rect 52700 43880 52730 43920
rect 52720 43722 52730 43880
rect 53700 44032 53708 44190
rect 53700 44000 53730 44032
rect 53770 44000 53790 44240
rect 53700 43920 53790 44000
rect 53700 43880 53730 43920
rect 52788 43818 52822 43834
rect 52856 43828 52872 43862
rect 53048 43828 53064 43862
rect 53354 43828 53370 43862
rect 53546 43828 53562 43862
rect 52788 43768 52822 43784
rect 53605 43818 53639 43834
rect 52856 43740 52872 43774
rect 53048 43740 53064 43774
rect 53354 43740 53370 43774
rect 53546 43740 53562 43774
rect 53605 43768 53639 43784
rect 52700 43680 52730 43722
rect 52640 43550 52730 43680
rect 53700 43722 53708 43880
rect 53700 43680 53730 43722
rect 53770 43680 53790 43920
rect 53700 43550 53790 43680
rect 57630 44240 57720 44360
rect 57630 43980 57650 44240
rect 57690 44190 57720 44240
rect 57710 44032 57720 44190
rect 58690 44240 58780 44360
rect 58690 44190 58720 44240
rect 57778 44128 57812 44144
rect 57846 44138 57862 44172
rect 58038 44138 58054 44172
rect 58344 44138 58360 44172
rect 58536 44138 58552 44172
rect 57778 44078 57812 44094
rect 58595 44128 58629 44144
rect 57846 44050 57862 44084
rect 58038 44050 58054 44084
rect 58344 44050 58360 44084
rect 58536 44050 58552 44084
rect 58595 44078 58629 44094
rect 57690 43980 57720 44032
rect 57630 43920 57720 43980
rect 57630 43680 57650 43920
rect 57690 43880 57720 43920
rect 57710 43722 57720 43880
rect 58690 44032 58698 44190
rect 58690 44000 58720 44032
rect 58760 44000 58780 44240
rect 58690 43920 58780 44000
rect 58690 43880 58720 43920
rect 57778 43818 57812 43834
rect 57846 43828 57862 43862
rect 58038 43828 58054 43862
rect 58344 43828 58360 43862
rect 58536 43828 58552 43862
rect 57778 43768 57812 43784
rect 58595 43818 58629 43834
rect 57846 43740 57862 43774
rect 58038 43740 58054 43774
rect 58344 43740 58360 43774
rect 58536 43740 58552 43774
rect 58595 43768 58629 43784
rect 57690 43680 57720 43722
rect 57630 43550 57720 43680
rect 58690 43722 58698 43880
rect 58690 43680 58720 43722
rect 58760 43680 58780 43920
rect 58690 43550 58780 43680
rect 62620 44240 62710 44360
rect 62620 43980 62640 44240
rect 62680 44190 62710 44240
rect 62700 44032 62710 44190
rect 63680 44240 63770 44360
rect 63680 44190 63710 44240
rect 62768 44128 62802 44144
rect 62836 44138 62852 44172
rect 63028 44138 63044 44172
rect 63334 44138 63350 44172
rect 63526 44138 63542 44172
rect 62768 44078 62802 44094
rect 63585 44128 63619 44144
rect 62836 44050 62852 44084
rect 63028 44050 63044 44084
rect 63334 44050 63350 44084
rect 63526 44050 63542 44084
rect 63585 44078 63619 44094
rect 62680 43980 62710 44032
rect 62620 43920 62710 43980
rect 62620 43680 62640 43920
rect 62680 43880 62710 43920
rect 62700 43722 62710 43880
rect 63680 44032 63688 44190
rect 63680 44000 63710 44032
rect 63750 44000 63770 44240
rect 63680 43920 63770 44000
rect 63680 43880 63710 43920
rect 62768 43818 62802 43834
rect 62836 43828 62852 43862
rect 63028 43828 63044 43862
rect 63334 43828 63350 43862
rect 63526 43828 63542 43862
rect 62768 43768 62802 43784
rect 63585 43818 63619 43834
rect 62836 43740 62852 43774
rect 63028 43740 63044 43774
rect 63334 43740 63350 43774
rect 63526 43740 63542 43774
rect 63585 43768 63619 43784
rect 62680 43680 62710 43722
rect 62620 43550 62710 43680
rect 63680 43722 63688 43880
rect 63680 43680 63710 43722
rect 63750 43680 63770 43920
rect 63680 43550 63770 43680
rect 67610 44240 67700 44360
rect 67610 43980 67630 44240
rect 67670 44190 67700 44240
rect 67690 44032 67700 44190
rect 68670 44240 68760 44360
rect 68670 44190 68700 44240
rect 67758 44128 67792 44144
rect 67826 44138 67842 44172
rect 68018 44138 68034 44172
rect 68324 44138 68340 44172
rect 68516 44138 68532 44172
rect 67758 44078 67792 44094
rect 68575 44128 68609 44144
rect 67826 44050 67842 44084
rect 68018 44050 68034 44084
rect 68324 44050 68340 44084
rect 68516 44050 68532 44084
rect 68575 44078 68609 44094
rect 67670 43980 67700 44032
rect 67610 43920 67700 43980
rect 67610 43680 67630 43920
rect 67670 43880 67700 43920
rect 67690 43722 67700 43880
rect 68670 44032 68678 44190
rect 68670 44000 68700 44032
rect 68740 44000 68760 44240
rect 68670 43920 68760 44000
rect 68670 43880 68700 43920
rect 67758 43818 67792 43834
rect 67826 43828 67842 43862
rect 68018 43828 68034 43862
rect 68324 43828 68340 43862
rect 68516 43828 68532 43862
rect 67758 43768 67792 43784
rect 68575 43818 68609 43834
rect 67826 43740 67842 43774
rect 68018 43740 68034 43774
rect 68324 43740 68340 43774
rect 68516 43740 68532 43774
rect 68575 43768 68609 43784
rect 67670 43680 67700 43722
rect 67610 43550 67700 43680
rect 68670 43722 68678 43880
rect 68670 43680 68700 43722
rect 68740 43680 68760 43920
rect 68670 43550 68760 43680
rect 72600 44240 72690 44360
rect 72600 43980 72620 44240
rect 72660 44190 72690 44240
rect 72680 44032 72690 44190
rect 73660 44240 73750 44360
rect 73660 44190 73690 44240
rect 72748 44128 72782 44144
rect 72816 44138 72832 44172
rect 73008 44138 73024 44172
rect 73314 44138 73330 44172
rect 73506 44138 73522 44172
rect 72748 44078 72782 44094
rect 73565 44128 73599 44144
rect 72816 44050 72832 44084
rect 73008 44050 73024 44084
rect 73314 44050 73330 44084
rect 73506 44050 73522 44084
rect 73565 44078 73599 44094
rect 72660 43980 72690 44032
rect 72600 43920 72690 43980
rect 72600 43680 72620 43920
rect 72660 43880 72690 43920
rect 72680 43722 72690 43880
rect 73660 44032 73668 44190
rect 73660 44000 73690 44032
rect 73730 44000 73750 44240
rect 73660 43920 73750 44000
rect 73660 43880 73690 43920
rect 72748 43818 72782 43834
rect 72816 43828 72832 43862
rect 73008 43828 73024 43862
rect 73314 43828 73330 43862
rect 73506 43828 73522 43862
rect 72748 43768 72782 43784
rect 73565 43818 73599 43834
rect 72816 43740 72832 43774
rect 73008 43740 73024 43774
rect 73314 43740 73330 43774
rect 73506 43740 73522 43774
rect 73565 43768 73599 43784
rect 72660 43680 72690 43722
rect 72600 43550 72690 43680
rect 73660 43722 73668 43880
rect 73660 43680 73690 43722
rect 73730 43680 73750 43920
rect 73660 43550 73750 43680
rect 77590 44240 77680 44360
rect 77590 43980 77610 44240
rect 77650 44190 77680 44240
rect 77670 44032 77680 44190
rect 78650 44240 78740 44360
rect 78650 44190 78680 44240
rect 77738 44128 77772 44144
rect 77806 44138 77822 44172
rect 77998 44138 78014 44172
rect 78304 44138 78320 44172
rect 78496 44138 78512 44172
rect 77738 44078 77772 44094
rect 78555 44128 78589 44144
rect 77806 44050 77822 44084
rect 77998 44050 78014 44084
rect 78304 44050 78320 44084
rect 78496 44050 78512 44084
rect 78555 44078 78589 44094
rect 77650 43980 77680 44032
rect 77590 43920 77680 43980
rect 77590 43680 77610 43920
rect 77650 43880 77680 43920
rect 77670 43722 77680 43880
rect 78650 44032 78658 44190
rect 78650 44000 78680 44032
rect 78720 44000 78740 44240
rect 78650 43920 78740 44000
rect 78650 43880 78680 43920
rect 77738 43818 77772 43834
rect 77806 43828 77822 43862
rect 77998 43828 78014 43862
rect 78304 43828 78320 43862
rect 78496 43828 78512 43862
rect 77738 43768 77772 43784
rect 78555 43818 78589 43834
rect 77806 43740 77822 43774
rect 77998 43740 78014 43774
rect 78304 43740 78320 43774
rect 78496 43740 78512 43774
rect 78555 43768 78589 43784
rect 77650 43680 77680 43722
rect 77590 43550 77680 43680
rect 78650 43722 78658 43880
rect 78650 43680 78680 43722
rect 78720 43680 78740 43920
rect 78650 43550 78740 43680
rect 2740 42530 2830 42650
rect 2740 42270 2760 42530
rect 2800 42480 2830 42530
rect 2820 42322 2830 42480
rect 3800 42530 3890 42650
rect 3800 42480 3830 42530
rect 2888 42418 2922 42434
rect 2956 42428 2972 42462
rect 3148 42428 3164 42462
rect 3454 42428 3470 42462
rect 3646 42428 3662 42462
rect 2888 42368 2922 42384
rect 3705 42418 3739 42434
rect 2956 42340 2972 42374
rect 3148 42340 3164 42374
rect 3454 42340 3470 42374
rect 3646 42340 3662 42374
rect 3705 42368 3739 42384
rect 2800 42270 2830 42322
rect 2740 42210 2830 42270
rect 2740 41970 2760 42210
rect 2800 42170 2830 42210
rect 2820 42012 2830 42170
rect 3800 42322 3808 42480
rect 3800 42290 3830 42322
rect 3870 42290 3890 42530
rect 3800 42210 3890 42290
rect 3800 42170 3830 42210
rect 2888 42108 2922 42124
rect 2956 42118 2972 42152
rect 3148 42118 3164 42152
rect 3454 42118 3470 42152
rect 3646 42118 3662 42152
rect 2888 42058 2922 42074
rect 3705 42108 3739 42124
rect 2956 42030 2972 42064
rect 3148 42030 3164 42064
rect 3454 42030 3470 42064
rect 3646 42030 3662 42064
rect 3705 42058 3739 42074
rect 2800 41970 2830 42012
rect 2740 41840 2830 41970
rect 3800 42012 3808 42170
rect 3800 41970 3830 42012
rect 3870 41970 3890 42210
rect 3800 41840 3890 41970
rect 7730 42530 7820 42650
rect 7730 42270 7750 42530
rect 7790 42480 7820 42530
rect 7810 42322 7820 42480
rect 8790 42530 8880 42650
rect 8790 42480 8820 42530
rect 7878 42418 7912 42434
rect 7946 42428 7962 42462
rect 8138 42428 8154 42462
rect 8444 42428 8460 42462
rect 8636 42428 8652 42462
rect 7878 42368 7912 42384
rect 8695 42418 8729 42434
rect 7946 42340 7962 42374
rect 8138 42340 8154 42374
rect 8444 42340 8460 42374
rect 8636 42340 8652 42374
rect 8695 42368 8729 42384
rect 7790 42270 7820 42322
rect 7730 42210 7820 42270
rect 7730 41970 7750 42210
rect 7790 42170 7820 42210
rect 7810 42012 7820 42170
rect 8790 42322 8798 42480
rect 8790 42290 8820 42322
rect 8860 42290 8880 42530
rect 8790 42210 8880 42290
rect 8790 42170 8820 42210
rect 7878 42108 7912 42124
rect 7946 42118 7962 42152
rect 8138 42118 8154 42152
rect 8444 42118 8460 42152
rect 8636 42118 8652 42152
rect 7878 42058 7912 42074
rect 8695 42108 8729 42124
rect 7946 42030 7962 42064
rect 8138 42030 8154 42064
rect 8444 42030 8460 42064
rect 8636 42030 8652 42064
rect 8695 42058 8729 42074
rect 7790 41970 7820 42012
rect 7730 41840 7820 41970
rect 8790 42012 8798 42170
rect 8790 41970 8820 42012
rect 8860 41970 8880 42210
rect 8790 41840 8880 41970
rect 12720 42530 12810 42650
rect 12720 42270 12740 42530
rect 12780 42480 12810 42530
rect 12800 42322 12810 42480
rect 13780 42530 13870 42650
rect 13780 42480 13810 42530
rect 12868 42418 12902 42434
rect 12936 42428 12952 42462
rect 13128 42428 13144 42462
rect 13434 42428 13450 42462
rect 13626 42428 13642 42462
rect 12868 42368 12902 42384
rect 13685 42418 13719 42434
rect 12936 42340 12952 42374
rect 13128 42340 13144 42374
rect 13434 42340 13450 42374
rect 13626 42340 13642 42374
rect 13685 42368 13719 42384
rect 12780 42270 12810 42322
rect 12720 42210 12810 42270
rect 12720 41970 12740 42210
rect 12780 42170 12810 42210
rect 12800 42012 12810 42170
rect 13780 42322 13788 42480
rect 13780 42290 13810 42322
rect 13850 42290 13870 42530
rect 13780 42210 13870 42290
rect 13780 42170 13810 42210
rect 12868 42108 12902 42124
rect 12936 42118 12952 42152
rect 13128 42118 13144 42152
rect 13434 42118 13450 42152
rect 13626 42118 13642 42152
rect 12868 42058 12902 42074
rect 13685 42108 13719 42124
rect 12936 42030 12952 42064
rect 13128 42030 13144 42064
rect 13434 42030 13450 42064
rect 13626 42030 13642 42064
rect 13685 42058 13719 42074
rect 12780 41970 12810 42012
rect 12720 41840 12810 41970
rect 13780 42012 13788 42170
rect 13780 41970 13810 42012
rect 13850 41970 13870 42210
rect 13780 41840 13870 41970
rect 17710 42530 17800 42650
rect 17710 42270 17730 42530
rect 17770 42480 17800 42530
rect 17790 42322 17800 42480
rect 18770 42530 18860 42650
rect 18770 42480 18800 42530
rect 17858 42418 17892 42434
rect 17926 42428 17942 42462
rect 18118 42428 18134 42462
rect 18424 42428 18440 42462
rect 18616 42428 18632 42462
rect 17858 42368 17892 42384
rect 18675 42418 18709 42434
rect 17926 42340 17942 42374
rect 18118 42340 18134 42374
rect 18424 42340 18440 42374
rect 18616 42340 18632 42374
rect 18675 42368 18709 42384
rect 17770 42270 17800 42322
rect 17710 42210 17800 42270
rect 17710 41970 17730 42210
rect 17770 42170 17800 42210
rect 17790 42012 17800 42170
rect 18770 42322 18778 42480
rect 18770 42290 18800 42322
rect 18840 42290 18860 42530
rect 18770 42210 18860 42290
rect 18770 42170 18800 42210
rect 17858 42108 17892 42124
rect 17926 42118 17942 42152
rect 18118 42118 18134 42152
rect 18424 42118 18440 42152
rect 18616 42118 18632 42152
rect 17858 42058 17892 42074
rect 18675 42108 18709 42124
rect 17926 42030 17942 42064
rect 18118 42030 18134 42064
rect 18424 42030 18440 42064
rect 18616 42030 18632 42064
rect 18675 42058 18709 42074
rect 17770 41970 17800 42012
rect 17710 41840 17800 41970
rect 18770 42012 18778 42170
rect 18770 41970 18800 42012
rect 18840 41970 18860 42210
rect 18770 41840 18860 41970
rect 22700 42530 22790 42650
rect 22700 42270 22720 42530
rect 22760 42480 22790 42530
rect 22780 42322 22790 42480
rect 23760 42530 23850 42650
rect 23760 42480 23790 42530
rect 22848 42418 22882 42434
rect 22916 42428 22932 42462
rect 23108 42428 23124 42462
rect 23414 42428 23430 42462
rect 23606 42428 23622 42462
rect 22848 42368 22882 42384
rect 23665 42418 23699 42434
rect 22916 42340 22932 42374
rect 23108 42340 23124 42374
rect 23414 42340 23430 42374
rect 23606 42340 23622 42374
rect 23665 42368 23699 42384
rect 22760 42270 22790 42322
rect 22700 42210 22790 42270
rect 22700 41970 22720 42210
rect 22760 42170 22790 42210
rect 22780 42012 22790 42170
rect 23760 42322 23768 42480
rect 23760 42290 23790 42322
rect 23830 42290 23850 42530
rect 23760 42210 23850 42290
rect 23760 42170 23790 42210
rect 22848 42108 22882 42124
rect 22916 42118 22932 42152
rect 23108 42118 23124 42152
rect 23414 42118 23430 42152
rect 23606 42118 23622 42152
rect 22848 42058 22882 42074
rect 23665 42108 23699 42124
rect 22916 42030 22932 42064
rect 23108 42030 23124 42064
rect 23414 42030 23430 42064
rect 23606 42030 23622 42064
rect 23665 42058 23699 42074
rect 22760 41970 22790 42012
rect 22700 41840 22790 41970
rect 23760 42012 23768 42170
rect 23760 41970 23790 42012
rect 23830 41970 23850 42210
rect 23760 41840 23850 41970
rect 27690 42530 27780 42650
rect 27690 42270 27710 42530
rect 27750 42480 27780 42530
rect 27770 42322 27780 42480
rect 28750 42530 28840 42650
rect 28750 42480 28780 42530
rect 27838 42418 27872 42434
rect 27906 42428 27922 42462
rect 28098 42428 28114 42462
rect 28404 42428 28420 42462
rect 28596 42428 28612 42462
rect 27838 42368 27872 42384
rect 28655 42418 28689 42434
rect 27906 42340 27922 42374
rect 28098 42340 28114 42374
rect 28404 42340 28420 42374
rect 28596 42340 28612 42374
rect 28655 42368 28689 42384
rect 27750 42270 27780 42322
rect 27690 42210 27780 42270
rect 27690 41970 27710 42210
rect 27750 42170 27780 42210
rect 27770 42012 27780 42170
rect 28750 42322 28758 42480
rect 28750 42290 28780 42322
rect 28820 42290 28840 42530
rect 28750 42210 28840 42290
rect 28750 42170 28780 42210
rect 27838 42108 27872 42124
rect 27906 42118 27922 42152
rect 28098 42118 28114 42152
rect 28404 42118 28420 42152
rect 28596 42118 28612 42152
rect 27838 42058 27872 42074
rect 28655 42108 28689 42124
rect 27906 42030 27922 42064
rect 28098 42030 28114 42064
rect 28404 42030 28420 42064
rect 28596 42030 28612 42064
rect 28655 42058 28689 42074
rect 27750 41970 27780 42012
rect 27690 41840 27780 41970
rect 28750 42012 28758 42170
rect 28750 41970 28780 42012
rect 28820 41970 28840 42210
rect 28750 41840 28840 41970
rect 32680 42530 32770 42650
rect 32680 42270 32700 42530
rect 32740 42480 32770 42530
rect 32760 42322 32770 42480
rect 33740 42530 33830 42650
rect 33740 42480 33770 42530
rect 32828 42418 32862 42434
rect 32896 42428 32912 42462
rect 33088 42428 33104 42462
rect 33394 42428 33410 42462
rect 33586 42428 33602 42462
rect 32828 42368 32862 42384
rect 33645 42418 33679 42434
rect 32896 42340 32912 42374
rect 33088 42340 33104 42374
rect 33394 42340 33410 42374
rect 33586 42340 33602 42374
rect 33645 42368 33679 42384
rect 32740 42270 32770 42322
rect 32680 42210 32770 42270
rect 32680 41970 32700 42210
rect 32740 42170 32770 42210
rect 32760 42012 32770 42170
rect 33740 42322 33748 42480
rect 33740 42290 33770 42322
rect 33810 42290 33830 42530
rect 33740 42210 33830 42290
rect 33740 42170 33770 42210
rect 32828 42108 32862 42124
rect 32896 42118 32912 42152
rect 33088 42118 33104 42152
rect 33394 42118 33410 42152
rect 33586 42118 33602 42152
rect 32828 42058 32862 42074
rect 33645 42108 33679 42124
rect 32896 42030 32912 42064
rect 33088 42030 33104 42064
rect 33394 42030 33410 42064
rect 33586 42030 33602 42064
rect 33645 42058 33679 42074
rect 32740 41970 32770 42012
rect 32680 41840 32770 41970
rect 33740 42012 33748 42170
rect 33740 41970 33770 42012
rect 33810 41970 33830 42210
rect 33740 41840 33830 41970
rect 37670 42530 37760 42650
rect 37670 42270 37690 42530
rect 37730 42480 37760 42530
rect 37750 42322 37760 42480
rect 38730 42530 38820 42650
rect 38730 42480 38760 42530
rect 37818 42418 37852 42434
rect 37886 42428 37902 42462
rect 38078 42428 38094 42462
rect 38384 42428 38400 42462
rect 38576 42428 38592 42462
rect 37818 42368 37852 42384
rect 38635 42418 38669 42434
rect 37886 42340 37902 42374
rect 38078 42340 38094 42374
rect 38384 42340 38400 42374
rect 38576 42340 38592 42374
rect 38635 42368 38669 42384
rect 37730 42270 37760 42322
rect 37670 42210 37760 42270
rect 37670 41970 37690 42210
rect 37730 42170 37760 42210
rect 37750 42012 37760 42170
rect 38730 42322 38738 42480
rect 38730 42290 38760 42322
rect 38800 42290 38820 42530
rect 38730 42210 38820 42290
rect 38730 42170 38760 42210
rect 37818 42108 37852 42124
rect 37886 42118 37902 42152
rect 38078 42118 38094 42152
rect 38384 42118 38400 42152
rect 38576 42118 38592 42152
rect 37818 42058 37852 42074
rect 38635 42108 38669 42124
rect 37886 42030 37902 42064
rect 38078 42030 38094 42064
rect 38384 42030 38400 42064
rect 38576 42030 38592 42064
rect 38635 42058 38669 42074
rect 37730 41970 37760 42012
rect 37670 41840 37760 41970
rect 38730 42012 38738 42170
rect 38730 41970 38760 42012
rect 38800 41970 38820 42210
rect 38730 41840 38820 41970
rect 42660 42530 42750 42650
rect 42660 42270 42680 42530
rect 42720 42480 42750 42530
rect 42740 42322 42750 42480
rect 43720 42530 43810 42650
rect 43720 42480 43750 42530
rect 42808 42418 42842 42434
rect 42876 42428 42892 42462
rect 43068 42428 43084 42462
rect 43374 42428 43390 42462
rect 43566 42428 43582 42462
rect 42808 42368 42842 42384
rect 43625 42418 43659 42434
rect 42876 42340 42892 42374
rect 43068 42340 43084 42374
rect 43374 42340 43390 42374
rect 43566 42340 43582 42374
rect 43625 42368 43659 42384
rect 42720 42270 42750 42322
rect 42660 42210 42750 42270
rect 42660 41970 42680 42210
rect 42720 42170 42750 42210
rect 42740 42012 42750 42170
rect 43720 42322 43728 42480
rect 43720 42290 43750 42322
rect 43790 42290 43810 42530
rect 43720 42210 43810 42290
rect 43720 42170 43750 42210
rect 42808 42108 42842 42124
rect 42876 42118 42892 42152
rect 43068 42118 43084 42152
rect 43374 42118 43390 42152
rect 43566 42118 43582 42152
rect 42808 42058 42842 42074
rect 43625 42108 43659 42124
rect 42876 42030 42892 42064
rect 43068 42030 43084 42064
rect 43374 42030 43390 42064
rect 43566 42030 43582 42064
rect 43625 42058 43659 42074
rect 42720 41970 42750 42012
rect 42660 41840 42750 41970
rect 43720 42012 43728 42170
rect 43720 41970 43750 42012
rect 43790 41970 43810 42210
rect 43720 41840 43810 41970
rect 47650 42530 47740 42650
rect 47650 42270 47670 42530
rect 47710 42480 47740 42530
rect 47730 42322 47740 42480
rect 48710 42530 48800 42650
rect 48710 42480 48740 42530
rect 47798 42418 47832 42434
rect 47866 42428 47882 42462
rect 48058 42428 48074 42462
rect 48364 42428 48380 42462
rect 48556 42428 48572 42462
rect 47798 42368 47832 42384
rect 48615 42418 48649 42434
rect 47866 42340 47882 42374
rect 48058 42340 48074 42374
rect 48364 42340 48380 42374
rect 48556 42340 48572 42374
rect 48615 42368 48649 42384
rect 47710 42270 47740 42322
rect 47650 42210 47740 42270
rect 47650 41970 47670 42210
rect 47710 42170 47740 42210
rect 47730 42012 47740 42170
rect 48710 42322 48718 42480
rect 48710 42290 48740 42322
rect 48780 42290 48800 42530
rect 48710 42210 48800 42290
rect 48710 42170 48740 42210
rect 47798 42108 47832 42124
rect 47866 42118 47882 42152
rect 48058 42118 48074 42152
rect 48364 42118 48380 42152
rect 48556 42118 48572 42152
rect 47798 42058 47832 42074
rect 48615 42108 48649 42124
rect 47866 42030 47882 42064
rect 48058 42030 48074 42064
rect 48364 42030 48380 42064
rect 48556 42030 48572 42064
rect 48615 42058 48649 42074
rect 47710 41970 47740 42012
rect 47650 41840 47740 41970
rect 48710 42012 48718 42170
rect 48710 41970 48740 42012
rect 48780 41970 48800 42210
rect 48710 41840 48800 41970
rect 52640 42530 52730 42650
rect 52640 42270 52660 42530
rect 52700 42480 52730 42530
rect 52720 42322 52730 42480
rect 53700 42530 53790 42650
rect 53700 42480 53730 42530
rect 52788 42418 52822 42434
rect 52856 42428 52872 42462
rect 53048 42428 53064 42462
rect 53354 42428 53370 42462
rect 53546 42428 53562 42462
rect 52788 42368 52822 42384
rect 53605 42418 53639 42434
rect 52856 42340 52872 42374
rect 53048 42340 53064 42374
rect 53354 42340 53370 42374
rect 53546 42340 53562 42374
rect 53605 42368 53639 42384
rect 52700 42270 52730 42322
rect 52640 42210 52730 42270
rect 52640 41970 52660 42210
rect 52700 42170 52730 42210
rect 52720 42012 52730 42170
rect 53700 42322 53708 42480
rect 53700 42290 53730 42322
rect 53770 42290 53790 42530
rect 53700 42210 53790 42290
rect 53700 42170 53730 42210
rect 52788 42108 52822 42124
rect 52856 42118 52872 42152
rect 53048 42118 53064 42152
rect 53354 42118 53370 42152
rect 53546 42118 53562 42152
rect 52788 42058 52822 42074
rect 53605 42108 53639 42124
rect 52856 42030 52872 42064
rect 53048 42030 53064 42064
rect 53354 42030 53370 42064
rect 53546 42030 53562 42064
rect 53605 42058 53639 42074
rect 52700 41970 52730 42012
rect 52640 41840 52730 41970
rect 53700 42012 53708 42170
rect 53700 41970 53730 42012
rect 53770 41970 53790 42210
rect 53700 41840 53790 41970
rect 57630 42530 57720 42650
rect 57630 42270 57650 42530
rect 57690 42480 57720 42530
rect 57710 42322 57720 42480
rect 58690 42530 58780 42650
rect 58690 42480 58720 42530
rect 57778 42418 57812 42434
rect 57846 42428 57862 42462
rect 58038 42428 58054 42462
rect 58344 42428 58360 42462
rect 58536 42428 58552 42462
rect 57778 42368 57812 42384
rect 58595 42418 58629 42434
rect 57846 42340 57862 42374
rect 58038 42340 58054 42374
rect 58344 42340 58360 42374
rect 58536 42340 58552 42374
rect 58595 42368 58629 42384
rect 57690 42270 57720 42322
rect 57630 42210 57720 42270
rect 57630 41970 57650 42210
rect 57690 42170 57720 42210
rect 57710 42012 57720 42170
rect 58690 42322 58698 42480
rect 58690 42290 58720 42322
rect 58760 42290 58780 42530
rect 58690 42210 58780 42290
rect 58690 42170 58720 42210
rect 57778 42108 57812 42124
rect 57846 42118 57862 42152
rect 58038 42118 58054 42152
rect 58344 42118 58360 42152
rect 58536 42118 58552 42152
rect 57778 42058 57812 42074
rect 58595 42108 58629 42124
rect 57846 42030 57862 42064
rect 58038 42030 58054 42064
rect 58344 42030 58360 42064
rect 58536 42030 58552 42064
rect 58595 42058 58629 42074
rect 57690 41970 57720 42012
rect 57630 41840 57720 41970
rect 58690 42012 58698 42170
rect 58690 41970 58720 42012
rect 58760 41970 58780 42210
rect 58690 41840 58780 41970
rect 62620 42530 62710 42650
rect 62620 42270 62640 42530
rect 62680 42480 62710 42530
rect 62700 42322 62710 42480
rect 63680 42530 63770 42650
rect 63680 42480 63710 42530
rect 62768 42418 62802 42434
rect 62836 42428 62852 42462
rect 63028 42428 63044 42462
rect 63334 42428 63350 42462
rect 63526 42428 63542 42462
rect 62768 42368 62802 42384
rect 63585 42418 63619 42434
rect 62836 42340 62852 42374
rect 63028 42340 63044 42374
rect 63334 42340 63350 42374
rect 63526 42340 63542 42374
rect 63585 42368 63619 42384
rect 62680 42270 62710 42322
rect 62620 42210 62710 42270
rect 62620 41970 62640 42210
rect 62680 42170 62710 42210
rect 62700 42012 62710 42170
rect 63680 42322 63688 42480
rect 63680 42290 63710 42322
rect 63750 42290 63770 42530
rect 63680 42210 63770 42290
rect 63680 42170 63710 42210
rect 62768 42108 62802 42124
rect 62836 42118 62852 42152
rect 63028 42118 63044 42152
rect 63334 42118 63350 42152
rect 63526 42118 63542 42152
rect 62768 42058 62802 42074
rect 63585 42108 63619 42124
rect 62836 42030 62852 42064
rect 63028 42030 63044 42064
rect 63334 42030 63350 42064
rect 63526 42030 63542 42064
rect 63585 42058 63619 42074
rect 62680 41970 62710 42012
rect 62620 41840 62710 41970
rect 63680 42012 63688 42170
rect 63680 41970 63710 42012
rect 63750 41970 63770 42210
rect 63680 41840 63770 41970
rect 67610 42530 67700 42650
rect 67610 42270 67630 42530
rect 67670 42480 67700 42530
rect 67690 42322 67700 42480
rect 68670 42530 68760 42650
rect 68670 42480 68700 42530
rect 67758 42418 67792 42434
rect 67826 42428 67842 42462
rect 68018 42428 68034 42462
rect 68324 42428 68340 42462
rect 68516 42428 68532 42462
rect 67758 42368 67792 42384
rect 68575 42418 68609 42434
rect 67826 42340 67842 42374
rect 68018 42340 68034 42374
rect 68324 42340 68340 42374
rect 68516 42340 68532 42374
rect 68575 42368 68609 42384
rect 67670 42270 67700 42322
rect 67610 42210 67700 42270
rect 67610 41970 67630 42210
rect 67670 42170 67700 42210
rect 67690 42012 67700 42170
rect 68670 42322 68678 42480
rect 68670 42290 68700 42322
rect 68740 42290 68760 42530
rect 68670 42210 68760 42290
rect 68670 42170 68700 42210
rect 67758 42108 67792 42124
rect 67826 42118 67842 42152
rect 68018 42118 68034 42152
rect 68324 42118 68340 42152
rect 68516 42118 68532 42152
rect 67758 42058 67792 42074
rect 68575 42108 68609 42124
rect 67826 42030 67842 42064
rect 68018 42030 68034 42064
rect 68324 42030 68340 42064
rect 68516 42030 68532 42064
rect 68575 42058 68609 42074
rect 67670 41970 67700 42012
rect 67610 41840 67700 41970
rect 68670 42012 68678 42170
rect 68670 41970 68700 42012
rect 68740 41970 68760 42210
rect 68670 41840 68760 41970
rect 72600 42530 72690 42650
rect 72600 42270 72620 42530
rect 72660 42480 72690 42530
rect 72680 42322 72690 42480
rect 73660 42530 73750 42650
rect 73660 42480 73690 42530
rect 72748 42418 72782 42434
rect 72816 42428 72832 42462
rect 73008 42428 73024 42462
rect 73314 42428 73330 42462
rect 73506 42428 73522 42462
rect 72748 42368 72782 42384
rect 73565 42418 73599 42434
rect 72816 42340 72832 42374
rect 73008 42340 73024 42374
rect 73314 42340 73330 42374
rect 73506 42340 73522 42374
rect 73565 42368 73599 42384
rect 72660 42270 72690 42322
rect 72600 42210 72690 42270
rect 72600 41970 72620 42210
rect 72660 42170 72690 42210
rect 72680 42012 72690 42170
rect 73660 42322 73668 42480
rect 73660 42290 73690 42322
rect 73730 42290 73750 42530
rect 73660 42210 73750 42290
rect 73660 42170 73690 42210
rect 72748 42108 72782 42124
rect 72816 42118 72832 42152
rect 73008 42118 73024 42152
rect 73314 42118 73330 42152
rect 73506 42118 73522 42152
rect 72748 42058 72782 42074
rect 73565 42108 73599 42124
rect 72816 42030 72832 42064
rect 73008 42030 73024 42064
rect 73314 42030 73330 42064
rect 73506 42030 73522 42064
rect 73565 42058 73599 42074
rect 72660 41970 72690 42012
rect 72600 41840 72690 41970
rect 73660 42012 73668 42170
rect 73660 41970 73690 42012
rect 73730 41970 73750 42210
rect 73660 41840 73750 41970
rect 77590 42530 77680 42650
rect 77590 42270 77610 42530
rect 77650 42480 77680 42530
rect 77670 42322 77680 42480
rect 78650 42530 78740 42650
rect 78650 42480 78680 42530
rect 77738 42418 77772 42434
rect 77806 42428 77822 42462
rect 77998 42428 78014 42462
rect 78304 42428 78320 42462
rect 78496 42428 78512 42462
rect 77738 42368 77772 42384
rect 78555 42418 78589 42434
rect 77806 42340 77822 42374
rect 77998 42340 78014 42374
rect 78304 42340 78320 42374
rect 78496 42340 78512 42374
rect 78555 42368 78589 42384
rect 77650 42270 77680 42322
rect 77590 42210 77680 42270
rect 77590 41970 77610 42210
rect 77650 42170 77680 42210
rect 77670 42012 77680 42170
rect 78650 42322 78658 42480
rect 78650 42290 78680 42322
rect 78720 42290 78740 42530
rect 78650 42210 78740 42290
rect 78650 42170 78680 42210
rect 77738 42108 77772 42124
rect 77806 42118 77822 42152
rect 77998 42118 78014 42152
rect 78304 42118 78320 42152
rect 78496 42118 78512 42152
rect 77738 42058 77772 42074
rect 78555 42108 78589 42124
rect 77806 42030 77822 42064
rect 77998 42030 78014 42064
rect 78304 42030 78320 42064
rect 78496 42030 78512 42064
rect 78555 42058 78589 42074
rect 77650 41970 77680 42012
rect 77590 41840 77680 41970
rect 78650 42012 78658 42170
rect 78650 41970 78680 42012
rect 78720 41970 78740 42210
rect 78650 41840 78740 41970
rect 2740 40820 2830 40940
rect 2740 40560 2760 40820
rect 2800 40770 2830 40820
rect 2820 40612 2830 40770
rect 3800 40820 3890 40940
rect 3800 40770 3830 40820
rect 2888 40708 2922 40724
rect 2956 40718 2972 40752
rect 3148 40718 3164 40752
rect 3454 40718 3470 40752
rect 3646 40718 3662 40752
rect 2888 40658 2922 40674
rect 3705 40708 3739 40724
rect 2956 40630 2972 40664
rect 3148 40630 3164 40664
rect 3454 40630 3470 40664
rect 3646 40630 3662 40664
rect 3705 40658 3739 40674
rect 2800 40560 2830 40612
rect 2740 40500 2830 40560
rect 2740 40260 2760 40500
rect 2800 40460 2830 40500
rect 2820 40302 2830 40460
rect 3800 40612 3808 40770
rect 3800 40580 3830 40612
rect 3870 40580 3890 40820
rect 3800 40500 3890 40580
rect 3800 40460 3830 40500
rect 2888 40398 2922 40414
rect 2956 40408 2972 40442
rect 3148 40408 3164 40442
rect 3454 40408 3470 40442
rect 3646 40408 3662 40442
rect 2888 40348 2922 40364
rect 3705 40398 3739 40414
rect 2956 40320 2972 40354
rect 3148 40320 3164 40354
rect 3454 40320 3470 40354
rect 3646 40320 3662 40354
rect 3705 40348 3739 40364
rect 2800 40260 2830 40302
rect 2740 40130 2830 40260
rect 3800 40302 3808 40460
rect 3800 40260 3830 40302
rect 3870 40260 3890 40500
rect 3800 40130 3890 40260
rect 7730 40820 7820 40940
rect 7730 40560 7750 40820
rect 7790 40770 7820 40820
rect 7810 40612 7820 40770
rect 8790 40820 8880 40940
rect 8790 40770 8820 40820
rect 7878 40708 7912 40724
rect 7946 40718 7962 40752
rect 8138 40718 8154 40752
rect 8444 40718 8460 40752
rect 8636 40718 8652 40752
rect 7878 40658 7912 40674
rect 8695 40708 8729 40724
rect 7946 40630 7962 40664
rect 8138 40630 8154 40664
rect 8444 40630 8460 40664
rect 8636 40630 8652 40664
rect 8695 40658 8729 40674
rect 7790 40560 7820 40612
rect 7730 40500 7820 40560
rect 7730 40260 7750 40500
rect 7790 40460 7820 40500
rect 7810 40302 7820 40460
rect 8790 40612 8798 40770
rect 8790 40580 8820 40612
rect 8860 40580 8880 40820
rect 8790 40500 8880 40580
rect 8790 40460 8820 40500
rect 7878 40398 7912 40414
rect 7946 40408 7962 40442
rect 8138 40408 8154 40442
rect 8444 40408 8460 40442
rect 8636 40408 8652 40442
rect 7878 40348 7912 40364
rect 8695 40398 8729 40414
rect 7946 40320 7962 40354
rect 8138 40320 8154 40354
rect 8444 40320 8460 40354
rect 8636 40320 8652 40354
rect 8695 40348 8729 40364
rect 7790 40260 7820 40302
rect 7730 40130 7820 40260
rect 8790 40302 8798 40460
rect 8790 40260 8820 40302
rect 8860 40260 8880 40500
rect 8790 40130 8880 40260
rect 12720 40820 12810 40940
rect 12720 40560 12740 40820
rect 12780 40770 12810 40820
rect 12800 40612 12810 40770
rect 13780 40820 13870 40940
rect 13780 40770 13810 40820
rect 12868 40708 12902 40724
rect 12936 40718 12952 40752
rect 13128 40718 13144 40752
rect 13434 40718 13450 40752
rect 13626 40718 13642 40752
rect 12868 40658 12902 40674
rect 13685 40708 13719 40724
rect 12936 40630 12952 40664
rect 13128 40630 13144 40664
rect 13434 40630 13450 40664
rect 13626 40630 13642 40664
rect 13685 40658 13719 40674
rect 12780 40560 12810 40612
rect 12720 40500 12810 40560
rect 12720 40260 12740 40500
rect 12780 40460 12810 40500
rect 12800 40302 12810 40460
rect 13780 40612 13788 40770
rect 13780 40580 13810 40612
rect 13850 40580 13870 40820
rect 13780 40500 13870 40580
rect 13780 40460 13810 40500
rect 12868 40398 12902 40414
rect 12936 40408 12952 40442
rect 13128 40408 13144 40442
rect 13434 40408 13450 40442
rect 13626 40408 13642 40442
rect 12868 40348 12902 40364
rect 13685 40398 13719 40414
rect 12936 40320 12952 40354
rect 13128 40320 13144 40354
rect 13434 40320 13450 40354
rect 13626 40320 13642 40354
rect 13685 40348 13719 40364
rect 12780 40260 12810 40302
rect 12720 40130 12810 40260
rect 13780 40302 13788 40460
rect 13780 40260 13810 40302
rect 13850 40260 13870 40500
rect 13780 40130 13870 40260
rect 17710 40820 17800 40940
rect 17710 40560 17730 40820
rect 17770 40770 17800 40820
rect 17790 40612 17800 40770
rect 18770 40820 18860 40940
rect 18770 40770 18800 40820
rect 17858 40708 17892 40724
rect 17926 40718 17942 40752
rect 18118 40718 18134 40752
rect 18424 40718 18440 40752
rect 18616 40718 18632 40752
rect 17858 40658 17892 40674
rect 18675 40708 18709 40724
rect 17926 40630 17942 40664
rect 18118 40630 18134 40664
rect 18424 40630 18440 40664
rect 18616 40630 18632 40664
rect 18675 40658 18709 40674
rect 17770 40560 17800 40612
rect 17710 40500 17800 40560
rect 17710 40260 17730 40500
rect 17770 40460 17800 40500
rect 17790 40302 17800 40460
rect 18770 40612 18778 40770
rect 18770 40580 18800 40612
rect 18840 40580 18860 40820
rect 18770 40500 18860 40580
rect 18770 40460 18800 40500
rect 17858 40398 17892 40414
rect 17926 40408 17942 40442
rect 18118 40408 18134 40442
rect 18424 40408 18440 40442
rect 18616 40408 18632 40442
rect 17858 40348 17892 40364
rect 18675 40398 18709 40414
rect 17926 40320 17942 40354
rect 18118 40320 18134 40354
rect 18424 40320 18440 40354
rect 18616 40320 18632 40354
rect 18675 40348 18709 40364
rect 17770 40260 17800 40302
rect 17710 40130 17800 40260
rect 18770 40302 18778 40460
rect 18770 40260 18800 40302
rect 18840 40260 18860 40500
rect 18770 40130 18860 40260
rect 22700 40820 22790 40940
rect 22700 40560 22720 40820
rect 22760 40770 22790 40820
rect 22780 40612 22790 40770
rect 23760 40820 23850 40940
rect 23760 40770 23790 40820
rect 22848 40708 22882 40724
rect 22916 40718 22932 40752
rect 23108 40718 23124 40752
rect 23414 40718 23430 40752
rect 23606 40718 23622 40752
rect 22848 40658 22882 40674
rect 23665 40708 23699 40724
rect 22916 40630 22932 40664
rect 23108 40630 23124 40664
rect 23414 40630 23430 40664
rect 23606 40630 23622 40664
rect 23665 40658 23699 40674
rect 22760 40560 22790 40612
rect 22700 40500 22790 40560
rect 22700 40260 22720 40500
rect 22760 40460 22790 40500
rect 22780 40302 22790 40460
rect 23760 40612 23768 40770
rect 23760 40580 23790 40612
rect 23830 40580 23850 40820
rect 23760 40500 23850 40580
rect 23760 40460 23790 40500
rect 22848 40398 22882 40414
rect 22916 40408 22932 40442
rect 23108 40408 23124 40442
rect 23414 40408 23430 40442
rect 23606 40408 23622 40442
rect 22848 40348 22882 40364
rect 23665 40398 23699 40414
rect 22916 40320 22932 40354
rect 23108 40320 23124 40354
rect 23414 40320 23430 40354
rect 23606 40320 23622 40354
rect 23665 40348 23699 40364
rect 22760 40260 22790 40302
rect 22700 40130 22790 40260
rect 23760 40302 23768 40460
rect 23760 40260 23790 40302
rect 23830 40260 23850 40500
rect 23760 40130 23850 40260
rect 27690 40820 27780 40940
rect 27690 40560 27710 40820
rect 27750 40770 27780 40820
rect 27770 40612 27780 40770
rect 28750 40820 28840 40940
rect 28750 40770 28780 40820
rect 27838 40708 27872 40724
rect 27906 40718 27922 40752
rect 28098 40718 28114 40752
rect 28404 40718 28420 40752
rect 28596 40718 28612 40752
rect 27838 40658 27872 40674
rect 28655 40708 28689 40724
rect 27906 40630 27922 40664
rect 28098 40630 28114 40664
rect 28404 40630 28420 40664
rect 28596 40630 28612 40664
rect 28655 40658 28689 40674
rect 27750 40560 27780 40612
rect 27690 40500 27780 40560
rect 27690 40260 27710 40500
rect 27750 40460 27780 40500
rect 27770 40302 27780 40460
rect 28750 40612 28758 40770
rect 28750 40580 28780 40612
rect 28820 40580 28840 40820
rect 28750 40500 28840 40580
rect 28750 40460 28780 40500
rect 27838 40398 27872 40414
rect 27906 40408 27922 40442
rect 28098 40408 28114 40442
rect 28404 40408 28420 40442
rect 28596 40408 28612 40442
rect 27838 40348 27872 40364
rect 28655 40398 28689 40414
rect 27906 40320 27922 40354
rect 28098 40320 28114 40354
rect 28404 40320 28420 40354
rect 28596 40320 28612 40354
rect 28655 40348 28689 40364
rect 27750 40260 27780 40302
rect 27690 40130 27780 40260
rect 28750 40302 28758 40460
rect 28750 40260 28780 40302
rect 28820 40260 28840 40500
rect 28750 40130 28840 40260
rect 32680 40820 32770 40940
rect 32680 40560 32700 40820
rect 32740 40770 32770 40820
rect 32760 40612 32770 40770
rect 33740 40820 33830 40940
rect 33740 40770 33770 40820
rect 32828 40708 32862 40724
rect 32896 40718 32912 40752
rect 33088 40718 33104 40752
rect 33394 40718 33410 40752
rect 33586 40718 33602 40752
rect 32828 40658 32862 40674
rect 33645 40708 33679 40724
rect 32896 40630 32912 40664
rect 33088 40630 33104 40664
rect 33394 40630 33410 40664
rect 33586 40630 33602 40664
rect 33645 40658 33679 40674
rect 32740 40560 32770 40612
rect 32680 40500 32770 40560
rect 32680 40260 32700 40500
rect 32740 40460 32770 40500
rect 32760 40302 32770 40460
rect 33740 40612 33748 40770
rect 33740 40580 33770 40612
rect 33810 40580 33830 40820
rect 33740 40500 33830 40580
rect 33740 40460 33770 40500
rect 32828 40398 32862 40414
rect 32896 40408 32912 40442
rect 33088 40408 33104 40442
rect 33394 40408 33410 40442
rect 33586 40408 33602 40442
rect 32828 40348 32862 40364
rect 33645 40398 33679 40414
rect 32896 40320 32912 40354
rect 33088 40320 33104 40354
rect 33394 40320 33410 40354
rect 33586 40320 33602 40354
rect 33645 40348 33679 40364
rect 32740 40260 32770 40302
rect 32680 40130 32770 40260
rect 33740 40302 33748 40460
rect 33740 40260 33770 40302
rect 33810 40260 33830 40500
rect 33740 40130 33830 40260
rect 37670 40820 37760 40940
rect 37670 40560 37690 40820
rect 37730 40770 37760 40820
rect 37750 40612 37760 40770
rect 38730 40820 38820 40940
rect 38730 40770 38760 40820
rect 37818 40708 37852 40724
rect 37886 40718 37902 40752
rect 38078 40718 38094 40752
rect 38384 40718 38400 40752
rect 38576 40718 38592 40752
rect 37818 40658 37852 40674
rect 38635 40708 38669 40724
rect 37886 40630 37902 40664
rect 38078 40630 38094 40664
rect 38384 40630 38400 40664
rect 38576 40630 38592 40664
rect 38635 40658 38669 40674
rect 37730 40560 37760 40612
rect 37670 40500 37760 40560
rect 37670 40260 37690 40500
rect 37730 40460 37760 40500
rect 37750 40302 37760 40460
rect 38730 40612 38738 40770
rect 38730 40580 38760 40612
rect 38800 40580 38820 40820
rect 38730 40500 38820 40580
rect 38730 40460 38760 40500
rect 37818 40398 37852 40414
rect 37886 40408 37902 40442
rect 38078 40408 38094 40442
rect 38384 40408 38400 40442
rect 38576 40408 38592 40442
rect 37818 40348 37852 40364
rect 38635 40398 38669 40414
rect 37886 40320 37902 40354
rect 38078 40320 38094 40354
rect 38384 40320 38400 40354
rect 38576 40320 38592 40354
rect 38635 40348 38669 40364
rect 37730 40260 37760 40302
rect 37670 40130 37760 40260
rect 38730 40302 38738 40460
rect 38730 40260 38760 40302
rect 38800 40260 38820 40500
rect 38730 40130 38820 40260
rect 42660 40820 42750 40940
rect 42660 40560 42680 40820
rect 42720 40770 42750 40820
rect 42740 40612 42750 40770
rect 43720 40820 43810 40940
rect 43720 40770 43750 40820
rect 42808 40708 42842 40724
rect 42876 40718 42892 40752
rect 43068 40718 43084 40752
rect 43374 40718 43390 40752
rect 43566 40718 43582 40752
rect 42808 40658 42842 40674
rect 43625 40708 43659 40724
rect 42876 40630 42892 40664
rect 43068 40630 43084 40664
rect 43374 40630 43390 40664
rect 43566 40630 43582 40664
rect 43625 40658 43659 40674
rect 42720 40560 42750 40612
rect 42660 40500 42750 40560
rect 42660 40260 42680 40500
rect 42720 40460 42750 40500
rect 42740 40302 42750 40460
rect 43720 40612 43728 40770
rect 43720 40580 43750 40612
rect 43790 40580 43810 40820
rect 43720 40500 43810 40580
rect 43720 40460 43750 40500
rect 42808 40398 42842 40414
rect 42876 40408 42892 40442
rect 43068 40408 43084 40442
rect 43374 40408 43390 40442
rect 43566 40408 43582 40442
rect 42808 40348 42842 40364
rect 43625 40398 43659 40414
rect 42876 40320 42892 40354
rect 43068 40320 43084 40354
rect 43374 40320 43390 40354
rect 43566 40320 43582 40354
rect 43625 40348 43659 40364
rect 42720 40260 42750 40302
rect 42660 40130 42750 40260
rect 43720 40302 43728 40460
rect 43720 40260 43750 40302
rect 43790 40260 43810 40500
rect 43720 40130 43810 40260
rect 47650 40820 47740 40940
rect 47650 40560 47670 40820
rect 47710 40770 47740 40820
rect 47730 40612 47740 40770
rect 48710 40820 48800 40940
rect 48710 40770 48740 40820
rect 47798 40708 47832 40724
rect 47866 40718 47882 40752
rect 48058 40718 48074 40752
rect 48364 40718 48380 40752
rect 48556 40718 48572 40752
rect 47798 40658 47832 40674
rect 48615 40708 48649 40724
rect 47866 40630 47882 40664
rect 48058 40630 48074 40664
rect 48364 40630 48380 40664
rect 48556 40630 48572 40664
rect 48615 40658 48649 40674
rect 47710 40560 47740 40612
rect 47650 40500 47740 40560
rect 47650 40260 47670 40500
rect 47710 40460 47740 40500
rect 47730 40302 47740 40460
rect 48710 40612 48718 40770
rect 48710 40580 48740 40612
rect 48780 40580 48800 40820
rect 48710 40500 48800 40580
rect 48710 40460 48740 40500
rect 47798 40398 47832 40414
rect 47866 40408 47882 40442
rect 48058 40408 48074 40442
rect 48364 40408 48380 40442
rect 48556 40408 48572 40442
rect 47798 40348 47832 40364
rect 48615 40398 48649 40414
rect 47866 40320 47882 40354
rect 48058 40320 48074 40354
rect 48364 40320 48380 40354
rect 48556 40320 48572 40354
rect 48615 40348 48649 40364
rect 47710 40260 47740 40302
rect 47650 40130 47740 40260
rect 48710 40302 48718 40460
rect 48710 40260 48740 40302
rect 48780 40260 48800 40500
rect 48710 40130 48800 40260
rect 52640 40820 52730 40940
rect 52640 40560 52660 40820
rect 52700 40770 52730 40820
rect 52720 40612 52730 40770
rect 53700 40820 53790 40940
rect 53700 40770 53730 40820
rect 52788 40708 52822 40724
rect 52856 40718 52872 40752
rect 53048 40718 53064 40752
rect 53354 40718 53370 40752
rect 53546 40718 53562 40752
rect 52788 40658 52822 40674
rect 53605 40708 53639 40724
rect 52856 40630 52872 40664
rect 53048 40630 53064 40664
rect 53354 40630 53370 40664
rect 53546 40630 53562 40664
rect 53605 40658 53639 40674
rect 52700 40560 52730 40612
rect 52640 40500 52730 40560
rect 52640 40260 52660 40500
rect 52700 40460 52730 40500
rect 52720 40302 52730 40460
rect 53700 40612 53708 40770
rect 53700 40580 53730 40612
rect 53770 40580 53790 40820
rect 53700 40500 53790 40580
rect 53700 40460 53730 40500
rect 52788 40398 52822 40414
rect 52856 40408 52872 40442
rect 53048 40408 53064 40442
rect 53354 40408 53370 40442
rect 53546 40408 53562 40442
rect 52788 40348 52822 40364
rect 53605 40398 53639 40414
rect 52856 40320 52872 40354
rect 53048 40320 53064 40354
rect 53354 40320 53370 40354
rect 53546 40320 53562 40354
rect 53605 40348 53639 40364
rect 52700 40260 52730 40302
rect 52640 40130 52730 40260
rect 53700 40302 53708 40460
rect 53700 40260 53730 40302
rect 53770 40260 53790 40500
rect 53700 40130 53790 40260
rect 57630 40820 57720 40940
rect 57630 40560 57650 40820
rect 57690 40770 57720 40820
rect 57710 40612 57720 40770
rect 58690 40820 58780 40940
rect 58690 40770 58720 40820
rect 57778 40708 57812 40724
rect 57846 40718 57862 40752
rect 58038 40718 58054 40752
rect 58344 40718 58360 40752
rect 58536 40718 58552 40752
rect 57778 40658 57812 40674
rect 58595 40708 58629 40724
rect 57846 40630 57862 40664
rect 58038 40630 58054 40664
rect 58344 40630 58360 40664
rect 58536 40630 58552 40664
rect 58595 40658 58629 40674
rect 57690 40560 57720 40612
rect 57630 40500 57720 40560
rect 57630 40260 57650 40500
rect 57690 40460 57720 40500
rect 57710 40302 57720 40460
rect 58690 40612 58698 40770
rect 58690 40580 58720 40612
rect 58760 40580 58780 40820
rect 58690 40500 58780 40580
rect 58690 40460 58720 40500
rect 57778 40398 57812 40414
rect 57846 40408 57862 40442
rect 58038 40408 58054 40442
rect 58344 40408 58360 40442
rect 58536 40408 58552 40442
rect 57778 40348 57812 40364
rect 58595 40398 58629 40414
rect 57846 40320 57862 40354
rect 58038 40320 58054 40354
rect 58344 40320 58360 40354
rect 58536 40320 58552 40354
rect 58595 40348 58629 40364
rect 57690 40260 57720 40302
rect 57630 40130 57720 40260
rect 58690 40302 58698 40460
rect 58690 40260 58720 40302
rect 58760 40260 58780 40500
rect 58690 40130 58780 40260
rect 62620 40820 62710 40940
rect 62620 40560 62640 40820
rect 62680 40770 62710 40820
rect 62700 40612 62710 40770
rect 63680 40820 63770 40940
rect 63680 40770 63710 40820
rect 62768 40708 62802 40724
rect 62836 40718 62852 40752
rect 63028 40718 63044 40752
rect 63334 40718 63350 40752
rect 63526 40718 63542 40752
rect 62768 40658 62802 40674
rect 63585 40708 63619 40724
rect 62836 40630 62852 40664
rect 63028 40630 63044 40664
rect 63334 40630 63350 40664
rect 63526 40630 63542 40664
rect 63585 40658 63619 40674
rect 62680 40560 62710 40612
rect 62620 40500 62710 40560
rect 62620 40260 62640 40500
rect 62680 40460 62710 40500
rect 62700 40302 62710 40460
rect 63680 40612 63688 40770
rect 63680 40580 63710 40612
rect 63750 40580 63770 40820
rect 63680 40500 63770 40580
rect 63680 40460 63710 40500
rect 62768 40398 62802 40414
rect 62836 40408 62852 40442
rect 63028 40408 63044 40442
rect 63334 40408 63350 40442
rect 63526 40408 63542 40442
rect 62768 40348 62802 40364
rect 63585 40398 63619 40414
rect 62836 40320 62852 40354
rect 63028 40320 63044 40354
rect 63334 40320 63350 40354
rect 63526 40320 63542 40354
rect 63585 40348 63619 40364
rect 62680 40260 62710 40302
rect 62620 40130 62710 40260
rect 63680 40302 63688 40460
rect 63680 40260 63710 40302
rect 63750 40260 63770 40500
rect 63680 40130 63770 40260
rect 67610 40820 67700 40940
rect 67610 40560 67630 40820
rect 67670 40770 67700 40820
rect 67690 40612 67700 40770
rect 68670 40820 68760 40940
rect 68670 40770 68700 40820
rect 67758 40708 67792 40724
rect 67826 40718 67842 40752
rect 68018 40718 68034 40752
rect 68324 40718 68340 40752
rect 68516 40718 68532 40752
rect 67758 40658 67792 40674
rect 68575 40708 68609 40724
rect 67826 40630 67842 40664
rect 68018 40630 68034 40664
rect 68324 40630 68340 40664
rect 68516 40630 68532 40664
rect 68575 40658 68609 40674
rect 67670 40560 67700 40612
rect 67610 40500 67700 40560
rect 67610 40260 67630 40500
rect 67670 40460 67700 40500
rect 67690 40302 67700 40460
rect 68670 40612 68678 40770
rect 68670 40580 68700 40612
rect 68740 40580 68760 40820
rect 68670 40500 68760 40580
rect 68670 40460 68700 40500
rect 67758 40398 67792 40414
rect 67826 40408 67842 40442
rect 68018 40408 68034 40442
rect 68324 40408 68340 40442
rect 68516 40408 68532 40442
rect 67758 40348 67792 40364
rect 68575 40398 68609 40414
rect 67826 40320 67842 40354
rect 68018 40320 68034 40354
rect 68324 40320 68340 40354
rect 68516 40320 68532 40354
rect 68575 40348 68609 40364
rect 67670 40260 67700 40302
rect 67610 40130 67700 40260
rect 68670 40302 68678 40460
rect 68670 40260 68700 40302
rect 68740 40260 68760 40500
rect 68670 40130 68760 40260
rect 72600 40820 72690 40940
rect 72600 40560 72620 40820
rect 72660 40770 72690 40820
rect 72680 40612 72690 40770
rect 73660 40820 73750 40940
rect 73660 40770 73690 40820
rect 72748 40708 72782 40724
rect 72816 40718 72832 40752
rect 73008 40718 73024 40752
rect 73314 40718 73330 40752
rect 73506 40718 73522 40752
rect 72748 40658 72782 40674
rect 73565 40708 73599 40724
rect 72816 40630 72832 40664
rect 73008 40630 73024 40664
rect 73314 40630 73330 40664
rect 73506 40630 73522 40664
rect 73565 40658 73599 40674
rect 72660 40560 72690 40612
rect 72600 40500 72690 40560
rect 72600 40260 72620 40500
rect 72660 40460 72690 40500
rect 72680 40302 72690 40460
rect 73660 40612 73668 40770
rect 73660 40580 73690 40612
rect 73730 40580 73750 40820
rect 73660 40500 73750 40580
rect 73660 40460 73690 40500
rect 72748 40398 72782 40414
rect 72816 40408 72832 40442
rect 73008 40408 73024 40442
rect 73314 40408 73330 40442
rect 73506 40408 73522 40442
rect 72748 40348 72782 40364
rect 73565 40398 73599 40414
rect 72816 40320 72832 40354
rect 73008 40320 73024 40354
rect 73314 40320 73330 40354
rect 73506 40320 73522 40354
rect 73565 40348 73599 40364
rect 72660 40260 72690 40302
rect 72600 40130 72690 40260
rect 73660 40302 73668 40460
rect 73660 40260 73690 40302
rect 73730 40260 73750 40500
rect 73660 40130 73750 40260
rect 77590 40820 77680 40940
rect 77590 40560 77610 40820
rect 77650 40770 77680 40820
rect 77670 40612 77680 40770
rect 78650 40820 78740 40940
rect 78650 40770 78680 40820
rect 77738 40708 77772 40724
rect 77806 40718 77822 40752
rect 77998 40718 78014 40752
rect 78304 40718 78320 40752
rect 78496 40718 78512 40752
rect 77738 40658 77772 40674
rect 78555 40708 78589 40724
rect 77806 40630 77822 40664
rect 77998 40630 78014 40664
rect 78304 40630 78320 40664
rect 78496 40630 78512 40664
rect 78555 40658 78589 40674
rect 77650 40560 77680 40612
rect 77590 40500 77680 40560
rect 77590 40260 77610 40500
rect 77650 40460 77680 40500
rect 77670 40302 77680 40460
rect 78650 40612 78658 40770
rect 78650 40580 78680 40612
rect 78720 40580 78740 40820
rect 78650 40500 78740 40580
rect 78650 40460 78680 40500
rect 77738 40398 77772 40414
rect 77806 40408 77822 40442
rect 77998 40408 78014 40442
rect 78304 40408 78320 40442
rect 78496 40408 78512 40442
rect 77738 40348 77772 40364
rect 78555 40398 78589 40414
rect 77806 40320 77822 40354
rect 77998 40320 78014 40354
rect 78304 40320 78320 40354
rect 78496 40320 78512 40354
rect 78555 40348 78589 40364
rect 77650 40260 77680 40302
rect 77590 40130 77680 40260
rect 78650 40302 78658 40460
rect 78650 40260 78680 40302
rect 78720 40260 78740 40500
rect 78650 40130 78740 40260
<< viali >>
rect 2760 66420 2800 66470
rect 2760 66262 2786 66420
rect 2786 66262 2800 66420
rect 3830 66420 3870 66470
rect 2972 66368 3148 66402
rect 3470 66368 3646 66402
rect 2888 66324 2922 66358
rect 3705 66324 3739 66358
rect 2972 66280 3148 66314
rect 3470 66280 3646 66314
rect 2760 66210 2800 66262
rect 2760 66110 2800 66150
rect 2760 65952 2786 66110
rect 2786 65952 2800 66110
rect 3830 66262 3842 66420
rect 3842 66262 3870 66420
rect 3830 66230 3870 66262
rect 3830 66110 3870 66150
rect 2972 66058 3148 66092
rect 3470 66058 3646 66092
rect 2888 66014 2922 66048
rect 3705 66014 3739 66048
rect 2972 65970 3148 66004
rect 3470 65970 3646 66004
rect 2760 65910 2800 65952
rect 3830 65952 3842 66110
rect 3842 65952 3870 66110
rect 3830 65910 3870 65952
rect 7750 66420 7790 66470
rect 7750 66262 7776 66420
rect 7776 66262 7790 66420
rect 8820 66420 8860 66470
rect 7962 66368 8138 66402
rect 8460 66368 8636 66402
rect 7878 66324 7912 66358
rect 8695 66324 8729 66358
rect 7962 66280 8138 66314
rect 8460 66280 8636 66314
rect 7750 66210 7790 66262
rect 7750 66110 7790 66150
rect 7750 65952 7776 66110
rect 7776 65952 7790 66110
rect 8820 66262 8832 66420
rect 8832 66262 8860 66420
rect 8820 66230 8860 66262
rect 8820 66110 8860 66150
rect 7962 66058 8138 66092
rect 8460 66058 8636 66092
rect 7878 66014 7912 66048
rect 8695 66014 8729 66048
rect 7962 65970 8138 66004
rect 8460 65970 8636 66004
rect 7750 65910 7790 65952
rect 8820 65952 8832 66110
rect 8832 65952 8860 66110
rect 8820 65910 8860 65952
rect 12740 66420 12780 66470
rect 12740 66262 12766 66420
rect 12766 66262 12780 66420
rect 13810 66420 13850 66470
rect 12952 66368 13128 66402
rect 13450 66368 13626 66402
rect 12868 66324 12902 66358
rect 13685 66324 13719 66358
rect 12952 66280 13128 66314
rect 13450 66280 13626 66314
rect 12740 66210 12780 66262
rect 12740 66110 12780 66150
rect 12740 65952 12766 66110
rect 12766 65952 12780 66110
rect 13810 66262 13822 66420
rect 13822 66262 13850 66420
rect 13810 66230 13850 66262
rect 13810 66110 13850 66150
rect 12952 66058 13128 66092
rect 13450 66058 13626 66092
rect 12868 66014 12902 66048
rect 13685 66014 13719 66048
rect 12952 65970 13128 66004
rect 13450 65970 13626 66004
rect 12740 65910 12780 65952
rect 13810 65952 13822 66110
rect 13822 65952 13850 66110
rect 13810 65910 13850 65952
rect 17730 66420 17770 66470
rect 17730 66262 17756 66420
rect 17756 66262 17770 66420
rect 18800 66420 18840 66470
rect 17942 66368 18118 66402
rect 18440 66368 18616 66402
rect 17858 66324 17892 66358
rect 18675 66324 18709 66358
rect 17942 66280 18118 66314
rect 18440 66280 18616 66314
rect 17730 66210 17770 66262
rect 17730 66110 17770 66150
rect 17730 65952 17756 66110
rect 17756 65952 17770 66110
rect 18800 66262 18812 66420
rect 18812 66262 18840 66420
rect 18800 66230 18840 66262
rect 18800 66110 18840 66150
rect 17942 66058 18118 66092
rect 18440 66058 18616 66092
rect 17858 66014 17892 66048
rect 18675 66014 18709 66048
rect 17942 65970 18118 66004
rect 18440 65970 18616 66004
rect 17730 65910 17770 65952
rect 18800 65952 18812 66110
rect 18812 65952 18840 66110
rect 18800 65910 18840 65952
rect 22720 66420 22760 66470
rect 22720 66262 22746 66420
rect 22746 66262 22760 66420
rect 23790 66420 23830 66470
rect 22932 66368 23108 66402
rect 23430 66368 23606 66402
rect 22848 66324 22882 66358
rect 23665 66324 23699 66358
rect 22932 66280 23108 66314
rect 23430 66280 23606 66314
rect 22720 66210 22760 66262
rect 22720 66110 22760 66150
rect 22720 65952 22746 66110
rect 22746 65952 22760 66110
rect 23790 66262 23802 66420
rect 23802 66262 23830 66420
rect 23790 66230 23830 66262
rect 23790 66110 23830 66150
rect 22932 66058 23108 66092
rect 23430 66058 23606 66092
rect 22848 66014 22882 66048
rect 23665 66014 23699 66048
rect 22932 65970 23108 66004
rect 23430 65970 23606 66004
rect 22720 65910 22760 65952
rect 23790 65952 23802 66110
rect 23802 65952 23830 66110
rect 23790 65910 23830 65952
rect 27710 66420 27750 66470
rect 27710 66262 27736 66420
rect 27736 66262 27750 66420
rect 28780 66420 28820 66470
rect 27922 66368 28098 66402
rect 28420 66368 28596 66402
rect 27838 66324 27872 66358
rect 28655 66324 28689 66358
rect 27922 66280 28098 66314
rect 28420 66280 28596 66314
rect 27710 66210 27750 66262
rect 27710 66110 27750 66150
rect 27710 65952 27736 66110
rect 27736 65952 27750 66110
rect 28780 66262 28792 66420
rect 28792 66262 28820 66420
rect 28780 66230 28820 66262
rect 28780 66110 28820 66150
rect 27922 66058 28098 66092
rect 28420 66058 28596 66092
rect 27838 66014 27872 66048
rect 28655 66014 28689 66048
rect 27922 65970 28098 66004
rect 28420 65970 28596 66004
rect 27710 65910 27750 65952
rect 28780 65952 28792 66110
rect 28792 65952 28820 66110
rect 28780 65910 28820 65952
rect 32700 66420 32740 66470
rect 32700 66262 32726 66420
rect 32726 66262 32740 66420
rect 33770 66420 33810 66470
rect 32912 66368 33088 66402
rect 33410 66368 33586 66402
rect 32828 66324 32862 66358
rect 33645 66324 33679 66358
rect 32912 66280 33088 66314
rect 33410 66280 33586 66314
rect 32700 66210 32740 66262
rect 32700 66110 32740 66150
rect 32700 65952 32726 66110
rect 32726 65952 32740 66110
rect 33770 66262 33782 66420
rect 33782 66262 33810 66420
rect 33770 66230 33810 66262
rect 33770 66110 33810 66150
rect 32912 66058 33088 66092
rect 33410 66058 33586 66092
rect 32828 66014 32862 66048
rect 33645 66014 33679 66048
rect 32912 65970 33088 66004
rect 33410 65970 33586 66004
rect 32700 65910 32740 65952
rect 33770 65952 33782 66110
rect 33782 65952 33810 66110
rect 33770 65910 33810 65952
rect 37690 66420 37730 66470
rect 37690 66262 37716 66420
rect 37716 66262 37730 66420
rect 38760 66420 38800 66470
rect 37902 66368 38078 66402
rect 38400 66368 38576 66402
rect 37818 66324 37852 66358
rect 38635 66324 38669 66358
rect 37902 66280 38078 66314
rect 38400 66280 38576 66314
rect 37690 66210 37730 66262
rect 37690 66110 37730 66150
rect 37690 65952 37716 66110
rect 37716 65952 37730 66110
rect 38760 66262 38772 66420
rect 38772 66262 38800 66420
rect 38760 66230 38800 66262
rect 38760 66110 38800 66150
rect 37902 66058 38078 66092
rect 38400 66058 38576 66092
rect 37818 66014 37852 66048
rect 38635 66014 38669 66048
rect 37902 65970 38078 66004
rect 38400 65970 38576 66004
rect 37690 65910 37730 65952
rect 38760 65952 38772 66110
rect 38772 65952 38800 66110
rect 38760 65910 38800 65952
rect 42680 66420 42720 66470
rect 42680 66262 42706 66420
rect 42706 66262 42720 66420
rect 43750 66420 43790 66470
rect 42892 66368 43068 66402
rect 43390 66368 43566 66402
rect 42808 66324 42842 66358
rect 43625 66324 43659 66358
rect 42892 66280 43068 66314
rect 43390 66280 43566 66314
rect 42680 66210 42720 66262
rect 42680 66110 42720 66150
rect 42680 65952 42706 66110
rect 42706 65952 42720 66110
rect 43750 66262 43762 66420
rect 43762 66262 43790 66420
rect 43750 66230 43790 66262
rect 43750 66110 43790 66150
rect 42892 66058 43068 66092
rect 43390 66058 43566 66092
rect 42808 66014 42842 66048
rect 43625 66014 43659 66048
rect 42892 65970 43068 66004
rect 43390 65970 43566 66004
rect 42680 65910 42720 65952
rect 43750 65952 43762 66110
rect 43762 65952 43790 66110
rect 43750 65910 43790 65952
rect 47670 66420 47710 66470
rect 47670 66262 47696 66420
rect 47696 66262 47710 66420
rect 48740 66420 48780 66470
rect 47882 66368 48058 66402
rect 48380 66368 48556 66402
rect 47798 66324 47832 66358
rect 48615 66324 48649 66358
rect 47882 66280 48058 66314
rect 48380 66280 48556 66314
rect 47670 66210 47710 66262
rect 47670 66110 47710 66150
rect 47670 65952 47696 66110
rect 47696 65952 47710 66110
rect 48740 66262 48752 66420
rect 48752 66262 48780 66420
rect 48740 66230 48780 66262
rect 48740 66110 48780 66150
rect 47882 66058 48058 66092
rect 48380 66058 48556 66092
rect 47798 66014 47832 66048
rect 48615 66014 48649 66048
rect 47882 65970 48058 66004
rect 48380 65970 48556 66004
rect 47670 65910 47710 65952
rect 48740 65952 48752 66110
rect 48752 65952 48780 66110
rect 48740 65910 48780 65952
rect 52660 66420 52700 66470
rect 52660 66262 52686 66420
rect 52686 66262 52700 66420
rect 53730 66420 53770 66470
rect 52872 66368 53048 66402
rect 53370 66368 53546 66402
rect 52788 66324 52822 66358
rect 53605 66324 53639 66358
rect 52872 66280 53048 66314
rect 53370 66280 53546 66314
rect 52660 66210 52700 66262
rect 52660 66110 52700 66150
rect 52660 65952 52686 66110
rect 52686 65952 52700 66110
rect 53730 66262 53742 66420
rect 53742 66262 53770 66420
rect 53730 66230 53770 66262
rect 53730 66110 53770 66150
rect 52872 66058 53048 66092
rect 53370 66058 53546 66092
rect 52788 66014 52822 66048
rect 53605 66014 53639 66048
rect 52872 65970 53048 66004
rect 53370 65970 53546 66004
rect 52660 65910 52700 65952
rect 53730 65952 53742 66110
rect 53742 65952 53770 66110
rect 53730 65910 53770 65952
rect 57650 66420 57690 66470
rect 57650 66262 57676 66420
rect 57676 66262 57690 66420
rect 58720 66420 58760 66470
rect 57862 66368 58038 66402
rect 58360 66368 58536 66402
rect 57778 66324 57812 66358
rect 58595 66324 58629 66358
rect 57862 66280 58038 66314
rect 58360 66280 58536 66314
rect 57650 66210 57690 66262
rect 57650 66110 57690 66150
rect 57650 65952 57676 66110
rect 57676 65952 57690 66110
rect 58720 66262 58732 66420
rect 58732 66262 58760 66420
rect 58720 66230 58760 66262
rect 58720 66110 58760 66150
rect 57862 66058 58038 66092
rect 58360 66058 58536 66092
rect 57778 66014 57812 66048
rect 58595 66014 58629 66048
rect 57862 65970 58038 66004
rect 58360 65970 58536 66004
rect 57650 65910 57690 65952
rect 58720 65952 58732 66110
rect 58732 65952 58760 66110
rect 58720 65910 58760 65952
rect 62640 66420 62680 66470
rect 62640 66262 62666 66420
rect 62666 66262 62680 66420
rect 63710 66420 63750 66470
rect 62852 66368 63028 66402
rect 63350 66368 63526 66402
rect 62768 66324 62802 66358
rect 63585 66324 63619 66358
rect 62852 66280 63028 66314
rect 63350 66280 63526 66314
rect 62640 66210 62680 66262
rect 62640 66110 62680 66150
rect 62640 65952 62666 66110
rect 62666 65952 62680 66110
rect 63710 66262 63722 66420
rect 63722 66262 63750 66420
rect 63710 66230 63750 66262
rect 63710 66110 63750 66150
rect 62852 66058 63028 66092
rect 63350 66058 63526 66092
rect 62768 66014 62802 66048
rect 63585 66014 63619 66048
rect 62852 65970 63028 66004
rect 63350 65970 63526 66004
rect 62640 65910 62680 65952
rect 63710 65952 63722 66110
rect 63722 65952 63750 66110
rect 63710 65910 63750 65952
rect 67630 66420 67670 66470
rect 67630 66262 67656 66420
rect 67656 66262 67670 66420
rect 68700 66420 68740 66470
rect 67842 66368 68018 66402
rect 68340 66368 68516 66402
rect 67758 66324 67792 66358
rect 68575 66324 68609 66358
rect 67842 66280 68018 66314
rect 68340 66280 68516 66314
rect 67630 66210 67670 66262
rect 67630 66110 67670 66150
rect 67630 65952 67656 66110
rect 67656 65952 67670 66110
rect 68700 66262 68712 66420
rect 68712 66262 68740 66420
rect 68700 66230 68740 66262
rect 68700 66110 68740 66150
rect 67842 66058 68018 66092
rect 68340 66058 68516 66092
rect 67758 66014 67792 66048
rect 68575 66014 68609 66048
rect 67842 65970 68018 66004
rect 68340 65970 68516 66004
rect 67630 65910 67670 65952
rect 68700 65952 68712 66110
rect 68712 65952 68740 66110
rect 68700 65910 68740 65952
rect 72620 66420 72660 66470
rect 72620 66262 72646 66420
rect 72646 66262 72660 66420
rect 73690 66420 73730 66470
rect 72832 66368 73008 66402
rect 73330 66368 73506 66402
rect 72748 66324 72782 66358
rect 73565 66324 73599 66358
rect 72832 66280 73008 66314
rect 73330 66280 73506 66314
rect 72620 66210 72660 66262
rect 72620 66110 72660 66150
rect 72620 65952 72646 66110
rect 72646 65952 72660 66110
rect 73690 66262 73702 66420
rect 73702 66262 73730 66420
rect 73690 66230 73730 66262
rect 73690 66110 73730 66150
rect 72832 66058 73008 66092
rect 73330 66058 73506 66092
rect 72748 66014 72782 66048
rect 73565 66014 73599 66048
rect 72832 65970 73008 66004
rect 73330 65970 73506 66004
rect 72620 65910 72660 65952
rect 73690 65952 73702 66110
rect 73702 65952 73730 66110
rect 73690 65910 73730 65952
rect 77610 66420 77650 66470
rect 77610 66262 77636 66420
rect 77636 66262 77650 66420
rect 78680 66420 78720 66470
rect 77822 66368 77998 66402
rect 78320 66368 78496 66402
rect 77738 66324 77772 66358
rect 78555 66324 78589 66358
rect 77822 66280 77998 66314
rect 78320 66280 78496 66314
rect 77610 66210 77650 66262
rect 77610 66110 77650 66150
rect 77610 65952 77636 66110
rect 77636 65952 77650 66110
rect 78680 66262 78692 66420
rect 78692 66262 78720 66420
rect 78680 66230 78720 66262
rect 78680 66110 78720 66150
rect 77822 66058 77998 66092
rect 78320 66058 78496 66092
rect 77738 66014 77772 66048
rect 78555 66014 78589 66048
rect 77822 65970 77998 66004
rect 78320 65970 78496 66004
rect 77610 65910 77650 65952
rect 78680 65952 78692 66110
rect 78692 65952 78720 66110
rect 78680 65910 78720 65952
rect 2760 64710 2800 64760
rect 2760 64552 2786 64710
rect 2786 64552 2800 64710
rect 3830 64710 3870 64760
rect 2972 64658 3148 64692
rect 3470 64658 3646 64692
rect 2888 64614 2922 64648
rect 3705 64614 3739 64648
rect 2972 64570 3148 64604
rect 3470 64570 3646 64604
rect 2760 64500 2800 64552
rect 2760 64400 2800 64440
rect 2760 64242 2786 64400
rect 2786 64242 2800 64400
rect 3830 64552 3842 64710
rect 3842 64552 3870 64710
rect 3830 64520 3870 64552
rect 3830 64400 3870 64440
rect 2972 64348 3148 64382
rect 3470 64348 3646 64382
rect 2888 64304 2922 64338
rect 3705 64304 3739 64338
rect 2972 64260 3148 64294
rect 3470 64260 3646 64294
rect 2760 64200 2800 64242
rect 3830 64242 3842 64400
rect 3842 64242 3870 64400
rect 3830 64200 3870 64242
rect 7750 64710 7790 64760
rect 7750 64552 7776 64710
rect 7776 64552 7790 64710
rect 8820 64710 8860 64760
rect 7962 64658 8138 64692
rect 8460 64658 8636 64692
rect 7878 64614 7912 64648
rect 8695 64614 8729 64648
rect 7962 64570 8138 64604
rect 8460 64570 8636 64604
rect 7750 64500 7790 64552
rect 7750 64400 7790 64440
rect 7750 64242 7776 64400
rect 7776 64242 7790 64400
rect 8820 64552 8832 64710
rect 8832 64552 8860 64710
rect 8820 64520 8860 64552
rect 8820 64400 8860 64440
rect 7962 64348 8138 64382
rect 8460 64348 8636 64382
rect 7878 64304 7912 64338
rect 8695 64304 8729 64338
rect 7962 64260 8138 64294
rect 8460 64260 8636 64294
rect 7750 64200 7790 64242
rect 8820 64242 8832 64400
rect 8832 64242 8860 64400
rect 8820 64200 8860 64242
rect 12740 64710 12780 64760
rect 12740 64552 12766 64710
rect 12766 64552 12780 64710
rect 13810 64710 13850 64760
rect 12952 64658 13128 64692
rect 13450 64658 13626 64692
rect 12868 64614 12902 64648
rect 13685 64614 13719 64648
rect 12952 64570 13128 64604
rect 13450 64570 13626 64604
rect 12740 64500 12780 64552
rect 12740 64400 12780 64440
rect 12740 64242 12766 64400
rect 12766 64242 12780 64400
rect 13810 64552 13822 64710
rect 13822 64552 13850 64710
rect 13810 64520 13850 64552
rect 13810 64400 13850 64440
rect 12952 64348 13128 64382
rect 13450 64348 13626 64382
rect 12868 64304 12902 64338
rect 13685 64304 13719 64338
rect 12952 64260 13128 64294
rect 13450 64260 13626 64294
rect 12740 64200 12780 64242
rect 13810 64242 13822 64400
rect 13822 64242 13850 64400
rect 13810 64200 13850 64242
rect 17730 64710 17770 64760
rect 17730 64552 17756 64710
rect 17756 64552 17770 64710
rect 18800 64710 18840 64760
rect 17942 64658 18118 64692
rect 18440 64658 18616 64692
rect 17858 64614 17892 64648
rect 18675 64614 18709 64648
rect 17942 64570 18118 64604
rect 18440 64570 18616 64604
rect 17730 64500 17770 64552
rect 17730 64400 17770 64440
rect 17730 64242 17756 64400
rect 17756 64242 17770 64400
rect 18800 64552 18812 64710
rect 18812 64552 18840 64710
rect 18800 64520 18840 64552
rect 18800 64400 18840 64440
rect 17942 64348 18118 64382
rect 18440 64348 18616 64382
rect 17858 64304 17892 64338
rect 18675 64304 18709 64338
rect 17942 64260 18118 64294
rect 18440 64260 18616 64294
rect 17730 64200 17770 64242
rect 18800 64242 18812 64400
rect 18812 64242 18840 64400
rect 18800 64200 18840 64242
rect 22720 64710 22760 64760
rect 22720 64552 22746 64710
rect 22746 64552 22760 64710
rect 23790 64710 23830 64760
rect 22932 64658 23108 64692
rect 23430 64658 23606 64692
rect 22848 64614 22882 64648
rect 23665 64614 23699 64648
rect 22932 64570 23108 64604
rect 23430 64570 23606 64604
rect 22720 64500 22760 64552
rect 22720 64400 22760 64440
rect 22720 64242 22746 64400
rect 22746 64242 22760 64400
rect 23790 64552 23802 64710
rect 23802 64552 23830 64710
rect 23790 64520 23830 64552
rect 23790 64400 23830 64440
rect 22932 64348 23108 64382
rect 23430 64348 23606 64382
rect 22848 64304 22882 64338
rect 23665 64304 23699 64338
rect 22932 64260 23108 64294
rect 23430 64260 23606 64294
rect 22720 64200 22760 64242
rect 23790 64242 23802 64400
rect 23802 64242 23830 64400
rect 23790 64200 23830 64242
rect 27710 64710 27750 64760
rect 27710 64552 27736 64710
rect 27736 64552 27750 64710
rect 28780 64710 28820 64760
rect 27922 64658 28098 64692
rect 28420 64658 28596 64692
rect 27838 64614 27872 64648
rect 28655 64614 28689 64648
rect 27922 64570 28098 64604
rect 28420 64570 28596 64604
rect 27710 64500 27750 64552
rect 27710 64400 27750 64440
rect 27710 64242 27736 64400
rect 27736 64242 27750 64400
rect 28780 64552 28792 64710
rect 28792 64552 28820 64710
rect 28780 64520 28820 64552
rect 28780 64400 28820 64440
rect 27922 64348 28098 64382
rect 28420 64348 28596 64382
rect 27838 64304 27872 64338
rect 28655 64304 28689 64338
rect 27922 64260 28098 64294
rect 28420 64260 28596 64294
rect 27710 64200 27750 64242
rect 28780 64242 28792 64400
rect 28792 64242 28820 64400
rect 28780 64200 28820 64242
rect 32700 64710 32740 64760
rect 32700 64552 32726 64710
rect 32726 64552 32740 64710
rect 33770 64710 33810 64760
rect 32912 64658 33088 64692
rect 33410 64658 33586 64692
rect 32828 64614 32862 64648
rect 33645 64614 33679 64648
rect 32912 64570 33088 64604
rect 33410 64570 33586 64604
rect 32700 64500 32740 64552
rect 32700 64400 32740 64440
rect 32700 64242 32726 64400
rect 32726 64242 32740 64400
rect 33770 64552 33782 64710
rect 33782 64552 33810 64710
rect 33770 64520 33810 64552
rect 33770 64400 33810 64440
rect 32912 64348 33088 64382
rect 33410 64348 33586 64382
rect 32828 64304 32862 64338
rect 33645 64304 33679 64338
rect 32912 64260 33088 64294
rect 33410 64260 33586 64294
rect 32700 64200 32740 64242
rect 33770 64242 33782 64400
rect 33782 64242 33810 64400
rect 33770 64200 33810 64242
rect 37690 64710 37730 64760
rect 37690 64552 37716 64710
rect 37716 64552 37730 64710
rect 38760 64710 38800 64760
rect 37902 64658 38078 64692
rect 38400 64658 38576 64692
rect 37818 64614 37852 64648
rect 38635 64614 38669 64648
rect 37902 64570 38078 64604
rect 38400 64570 38576 64604
rect 37690 64500 37730 64552
rect 37690 64400 37730 64440
rect 37690 64242 37716 64400
rect 37716 64242 37730 64400
rect 38760 64552 38772 64710
rect 38772 64552 38800 64710
rect 38760 64520 38800 64552
rect 38760 64400 38800 64440
rect 37902 64348 38078 64382
rect 38400 64348 38576 64382
rect 37818 64304 37852 64338
rect 38635 64304 38669 64338
rect 37902 64260 38078 64294
rect 38400 64260 38576 64294
rect 37690 64200 37730 64242
rect 38760 64242 38772 64400
rect 38772 64242 38800 64400
rect 38760 64200 38800 64242
rect 42680 64710 42720 64760
rect 42680 64552 42706 64710
rect 42706 64552 42720 64710
rect 43750 64710 43790 64760
rect 42892 64658 43068 64692
rect 43390 64658 43566 64692
rect 42808 64614 42842 64648
rect 43625 64614 43659 64648
rect 42892 64570 43068 64604
rect 43390 64570 43566 64604
rect 42680 64500 42720 64552
rect 42680 64400 42720 64440
rect 42680 64242 42706 64400
rect 42706 64242 42720 64400
rect 43750 64552 43762 64710
rect 43762 64552 43790 64710
rect 43750 64520 43790 64552
rect 43750 64400 43790 64440
rect 42892 64348 43068 64382
rect 43390 64348 43566 64382
rect 42808 64304 42842 64338
rect 43625 64304 43659 64338
rect 42892 64260 43068 64294
rect 43390 64260 43566 64294
rect 42680 64200 42720 64242
rect 43750 64242 43762 64400
rect 43762 64242 43790 64400
rect 43750 64200 43790 64242
rect 47670 64710 47710 64760
rect 47670 64552 47696 64710
rect 47696 64552 47710 64710
rect 48740 64710 48780 64760
rect 47882 64658 48058 64692
rect 48380 64658 48556 64692
rect 47798 64614 47832 64648
rect 48615 64614 48649 64648
rect 47882 64570 48058 64604
rect 48380 64570 48556 64604
rect 47670 64500 47710 64552
rect 47670 64400 47710 64440
rect 47670 64242 47696 64400
rect 47696 64242 47710 64400
rect 48740 64552 48752 64710
rect 48752 64552 48780 64710
rect 48740 64520 48780 64552
rect 48740 64400 48780 64440
rect 47882 64348 48058 64382
rect 48380 64348 48556 64382
rect 47798 64304 47832 64338
rect 48615 64304 48649 64338
rect 47882 64260 48058 64294
rect 48380 64260 48556 64294
rect 47670 64200 47710 64242
rect 48740 64242 48752 64400
rect 48752 64242 48780 64400
rect 48740 64200 48780 64242
rect 52660 64710 52700 64760
rect 52660 64552 52686 64710
rect 52686 64552 52700 64710
rect 53730 64710 53770 64760
rect 52872 64658 53048 64692
rect 53370 64658 53546 64692
rect 52788 64614 52822 64648
rect 53605 64614 53639 64648
rect 52872 64570 53048 64604
rect 53370 64570 53546 64604
rect 52660 64500 52700 64552
rect 52660 64400 52700 64440
rect 52660 64242 52686 64400
rect 52686 64242 52700 64400
rect 53730 64552 53742 64710
rect 53742 64552 53770 64710
rect 53730 64520 53770 64552
rect 53730 64400 53770 64440
rect 52872 64348 53048 64382
rect 53370 64348 53546 64382
rect 52788 64304 52822 64338
rect 53605 64304 53639 64338
rect 52872 64260 53048 64294
rect 53370 64260 53546 64294
rect 52660 64200 52700 64242
rect 53730 64242 53742 64400
rect 53742 64242 53770 64400
rect 53730 64200 53770 64242
rect 57650 64710 57690 64760
rect 57650 64552 57676 64710
rect 57676 64552 57690 64710
rect 58720 64710 58760 64760
rect 57862 64658 58038 64692
rect 58360 64658 58536 64692
rect 57778 64614 57812 64648
rect 58595 64614 58629 64648
rect 57862 64570 58038 64604
rect 58360 64570 58536 64604
rect 57650 64500 57690 64552
rect 57650 64400 57690 64440
rect 57650 64242 57676 64400
rect 57676 64242 57690 64400
rect 58720 64552 58732 64710
rect 58732 64552 58760 64710
rect 58720 64520 58760 64552
rect 58720 64400 58760 64440
rect 57862 64348 58038 64382
rect 58360 64348 58536 64382
rect 57778 64304 57812 64338
rect 58595 64304 58629 64338
rect 57862 64260 58038 64294
rect 58360 64260 58536 64294
rect 57650 64200 57690 64242
rect 58720 64242 58732 64400
rect 58732 64242 58760 64400
rect 58720 64200 58760 64242
rect 62640 64710 62680 64760
rect 62640 64552 62666 64710
rect 62666 64552 62680 64710
rect 63710 64710 63750 64760
rect 62852 64658 63028 64692
rect 63350 64658 63526 64692
rect 62768 64614 62802 64648
rect 63585 64614 63619 64648
rect 62852 64570 63028 64604
rect 63350 64570 63526 64604
rect 62640 64500 62680 64552
rect 62640 64400 62680 64440
rect 62640 64242 62666 64400
rect 62666 64242 62680 64400
rect 63710 64552 63722 64710
rect 63722 64552 63750 64710
rect 63710 64520 63750 64552
rect 63710 64400 63750 64440
rect 62852 64348 63028 64382
rect 63350 64348 63526 64382
rect 62768 64304 62802 64338
rect 63585 64304 63619 64338
rect 62852 64260 63028 64294
rect 63350 64260 63526 64294
rect 62640 64200 62680 64242
rect 63710 64242 63722 64400
rect 63722 64242 63750 64400
rect 63710 64200 63750 64242
rect 67630 64710 67670 64760
rect 67630 64552 67656 64710
rect 67656 64552 67670 64710
rect 68700 64710 68740 64760
rect 67842 64658 68018 64692
rect 68340 64658 68516 64692
rect 67758 64614 67792 64648
rect 68575 64614 68609 64648
rect 67842 64570 68018 64604
rect 68340 64570 68516 64604
rect 67630 64500 67670 64552
rect 67630 64400 67670 64440
rect 67630 64242 67656 64400
rect 67656 64242 67670 64400
rect 68700 64552 68712 64710
rect 68712 64552 68740 64710
rect 68700 64520 68740 64552
rect 68700 64400 68740 64440
rect 67842 64348 68018 64382
rect 68340 64348 68516 64382
rect 67758 64304 67792 64338
rect 68575 64304 68609 64338
rect 67842 64260 68018 64294
rect 68340 64260 68516 64294
rect 67630 64200 67670 64242
rect 68700 64242 68712 64400
rect 68712 64242 68740 64400
rect 68700 64200 68740 64242
rect 72620 64710 72660 64760
rect 72620 64552 72646 64710
rect 72646 64552 72660 64710
rect 73690 64710 73730 64760
rect 72832 64658 73008 64692
rect 73330 64658 73506 64692
rect 72748 64614 72782 64648
rect 73565 64614 73599 64648
rect 72832 64570 73008 64604
rect 73330 64570 73506 64604
rect 72620 64500 72660 64552
rect 72620 64400 72660 64440
rect 72620 64242 72646 64400
rect 72646 64242 72660 64400
rect 73690 64552 73702 64710
rect 73702 64552 73730 64710
rect 73690 64520 73730 64552
rect 73690 64400 73730 64440
rect 72832 64348 73008 64382
rect 73330 64348 73506 64382
rect 72748 64304 72782 64338
rect 73565 64304 73599 64338
rect 72832 64260 73008 64294
rect 73330 64260 73506 64294
rect 72620 64200 72660 64242
rect 73690 64242 73702 64400
rect 73702 64242 73730 64400
rect 73690 64200 73730 64242
rect 77610 64710 77650 64760
rect 77610 64552 77636 64710
rect 77636 64552 77650 64710
rect 78680 64710 78720 64760
rect 77822 64658 77998 64692
rect 78320 64658 78496 64692
rect 77738 64614 77772 64648
rect 78555 64614 78589 64648
rect 77822 64570 77998 64604
rect 78320 64570 78496 64604
rect 77610 64500 77650 64552
rect 77610 64400 77650 64440
rect 77610 64242 77636 64400
rect 77636 64242 77650 64400
rect 78680 64552 78692 64710
rect 78692 64552 78720 64710
rect 78680 64520 78720 64552
rect 78680 64400 78720 64440
rect 77822 64348 77998 64382
rect 78320 64348 78496 64382
rect 77738 64304 77772 64338
rect 78555 64304 78589 64338
rect 77822 64260 77998 64294
rect 78320 64260 78496 64294
rect 77610 64200 77650 64242
rect 78680 64242 78692 64400
rect 78692 64242 78720 64400
rect 78680 64200 78720 64242
rect 2760 63000 2800 63050
rect 2760 62842 2786 63000
rect 2786 62842 2800 63000
rect 3830 63000 3870 63050
rect 2972 62948 3148 62982
rect 3470 62948 3646 62982
rect 2888 62904 2922 62938
rect 3705 62904 3739 62938
rect 2972 62860 3148 62894
rect 3470 62860 3646 62894
rect 2760 62790 2800 62842
rect 2760 62690 2800 62730
rect 2760 62532 2786 62690
rect 2786 62532 2800 62690
rect 3830 62842 3842 63000
rect 3842 62842 3870 63000
rect 3830 62810 3870 62842
rect 3830 62690 3870 62730
rect 2972 62638 3148 62672
rect 3470 62638 3646 62672
rect 2888 62594 2922 62628
rect 3705 62594 3739 62628
rect 2972 62550 3148 62584
rect 3470 62550 3646 62584
rect 2760 62490 2800 62532
rect 3830 62532 3842 62690
rect 3842 62532 3870 62690
rect 3830 62490 3870 62532
rect 7750 63000 7790 63050
rect 7750 62842 7776 63000
rect 7776 62842 7790 63000
rect 8820 63000 8860 63050
rect 7962 62948 8138 62982
rect 8460 62948 8636 62982
rect 7878 62904 7912 62938
rect 8695 62904 8729 62938
rect 7962 62860 8138 62894
rect 8460 62860 8636 62894
rect 7750 62790 7790 62842
rect 7750 62690 7790 62730
rect 7750 62532 7776 62690
rect 7776 62532 7790 62690
rect 8820 62842 8832 63000
rect 8832 62842 8860 63000
rect 8820 62810 8860 62842
rect 8820 62690 8860 62730
rect 7962 62638 8138 62672
rect 8460 62638 8636 62672
rect 7878 62594 7912 62628
rect 8695 62594 8729 62628
rect 7962 62550 8138 62584
rect 8460 62550 8636 62584
rect 7750 62490 7790 62532
rect 8820 62532 8832 62690
rect 8832 62532 8860 62690
rect 8820 62490 8860 62532
rect 12740 63000 12780 63050
rect 12740 62842 12766 63000
rect 12766 62842 12780 63000
rect 13810 63000 13850 63050
rect 12952 62948 13128 62982
rect 13450 62948 13626 62982
rect 12868 62904 12902 62938
rect 13685 62904 13719 62938
rect 12952 62860 13128 62894
rect 13450 62860 13626 62894
rect 12740 62790 12780 62842
rect 12740 62690 12780 62730
rect 12740 62532 12766 62690
rect 12766 62532 12780 62690
rect 13810 62842 13822 63000
rect 13822 62842 13850 63000
rect 13810 62810 13850 62842
rect 13810 62690 13850 62730
rect 12952 62638 13128 62672
rect 13450 62638 13626 62672
rect 12868 62594 12902 62628
rect 13685 62594 13719 62628
rect 12952 62550 13128 62584
rect 13450 62550 13626 62584
rect 12740 62490 12780 62532
rect 13810 62532 13822 62690
rect 13822 62532 13850 62690
rect 13810 62490 13850 62532
rect 17730 63000 17770 63050
rect 17730 62842 17756 63000
rect 17756 62842 17770 63000
rect 18800 63000 18840 63050
rect 17942 62948 18118 62982
rect 18440 62948 18616 62982
rect 17858 62904 17892 62938
rect 18675 62904 18709 62938
rect 17942 62860 18118 62894
rect 18440 62860 18616 62894
rect 17730 62790 17770 62842
rect 17730 62690 17770 62730
rect 17730 62532 17756 62690
rect 17756 62532 17770 62690
rect 18800 62842 18812 63000
rect 18812 62842 18840 63000
rect 18800 62810 18840 62842
rect 18800 62690 18840 62730
rect 17942 62638 18118 62672
rect 18440 62638 18616 62672
rect 17858 62594 17892 62628
rect 18675 62594 18709 62628
rect 17942 62550 18118 62584
rect 18440 62550 18616 62584
rect 17730 62490 17770 62532
rect 18800 62532 18812 62690
rect 18812 62532 18840 62690
rect 18800 62490 18840 62532
rect 22720 63000 22760 63050
rect 22720 62842 22746 63000
rect 22746 62842 22760 63000
rect 23790 63000 23830 63050
rect 22932 62948 23108 62982
rect 23430 62948 23606 62982
rect 22848 62904 22882 62938
rect 23665 62904 23699 62938
rect 22932 62860 23108 62894
rect 23430 62860 23606 62894
rect 22720 62790 22760 62842
rect 22720 62690 22760 62730
rect 22720 62532 22746 62690
rect 22746 62532 22760 62690
rect 23790 62842 23802 63000
rect 23802 62842 23830 63000
rect 23790 62810 23830 62842
rect 23790 62690 23830 62730
rect 22932 62638 23108 62672
rect 23430 62638 23606 62672
rect 22848 62594 22882 62628
rect 23665 62594 23699 62628
rect 22932 62550 23108 62584
rect 23430 62550 23606 62584
rect 22720 62490 22760 62532
rect 23790 62532 23802 62690
rect 23802 62532 23830 62690
rect 23790 62490 23830 62532
rect 27710 63000 27750 63050
rect 27710 62842 27736 63000
rect 27736 62842 27750 63000
rect 28780 63000 28820 63050
rect 27922 62948 28098 62982
rect 28420 62948 28596 62982
rect 27838 62904 27872 62938
rect 28655 62904 28689 62938
rect 27922 62860 28098 62894
rect 28420 62860 28596 62894
rect 27710 62790 27750 62842
rect 27710 62690 27750 62730
rect 27710 62532 27736 62690
rect 27736 62532 27750 62690
rect 28780 62842 28792 63000
rect 28792 62842 28820 63000
rect 28780 62810 28820 62842
rect 28780 62690 28820 62730
rect 27922 62638 28098 62672
rect 28420 62638 28596 62672
rect 27838 62594 27872 62628
rect 28655 62594 28689 62628
rect 27922 62550 28098 62584
rect 28420 62550 28596 62584
rect 27710 62490 27750 62532
rect 28780 62532 28792 62690
rect 28792 62532 28820 62690
rect 28780 62490 28820 62532
rect 32700 63000 32740 63050
rect 32700 62842 32726 63000
rect 32726 62842 32740 63000
rect 33770 63000 33810 63050
rect 32912 62948 33088 62982
rect 33410 62948 33586 62982
rect 32828 62904 32862 62938
rect 33645 62904 33679 62938
rect 32912 62860 33088 62894
rect 33410 62860 33586 62894
rect 32700 62790 32740 62842
rect 32700 62690 32740 62730
rect 32700 62532 32726 62690
rect 32726 62532 32740 62690
rect 33770 62842 33782 63000
rect 33782 62842 33810 63000
rect 33770 62810 33810 62842
rect 33770 62690 33810 62730
rect 32912 62638 33088 62672
rect 33410 62638 33586 62672
rect 32828 62594 32862 62628
rect 33645 62594 33679 62628
rect 32912 62550 33088 62584
rect 33410 62550 33586 62584
rect 32700 62490 32740 62532
rect 33770 62532 33782 62690
rect 33782 62532 33810 62690
rect 33770 62490 33810 62532
rect 37690 63000 37730 63050
rect 37690 62842 37716 63000
rect 37716 62842 37730 63000
rect 38760 63000 38800 63050
rect 37902 62948 38078 62982
rect 38400 62948 38576 62982
rect 37818 62904 37852 62938
rect 38635 62904 38669 62938
rect 37902 62860 38078 62894
rect 38400 62860 38576 62894
rect 37690 62790 37730 62842
rect 37690 62690 37730 62730
rect 37690 62532 37716 62690
rect 37716 62532 37730 62690
rect 38760 62842 38772 63000
rect 38772 62842 38800 63000
rect 38760 62810 38800 62842
rect 38760 62690 38800 62730
rect 37902 62638 38078 62672
rect 38400 62638 38576 62672
rect 37818 62594 37852 62628
rect 38635 62594 38669 62628
rect 37902 62550 38078 62584
rect 38400 62550 38576 62584
rect 37690 62490 37730 62532
rect 38760 62532 38772 62690
rect 38772 62532 38800 62690
rect 38760 62490 38800 62532
rect 42680 63000 42720 63050
rect 42680 62842 42706 63000
rect 42706 62842 42720 63000
rect 43750 63000 43790 63050
rect 42892 62948 43068 62982
rect 43390 62948 43566 62982
rect 42808 62904 42842 62938
rect 43625 62904 43659 62938
rect 42892 62860 43068 62894
rect 43390 62860 43566 62894
rect 42680 62790 42720 62842
rect 42680 62690 42720 62730
rect 42680 62532 42706 62690
rect 42706 62532 42720 62690
rect 43750 62842 43762 63000
rect 43762 62842 43790 63000
rect 43750 62810 43790 62842
rect 43750 62690 43790 62730
rect 42892 62638 43068 62672
rect 43390 62638 43566 62672
rect 42808 62594 42842 62628
rect 43625 62594 43659 62628
rect 42892 62550 43068 62584
rect 43390 62550 43566 62584
rect 42680 62490 42720 62532
rect 43750 62532 43762 62690
rect 43762 62532 43790 62690
rect 43750 62490 43790 62532
rect 47670 63000 47710 63050
rect 47670 62842 47696 63000
rect 47696 62842 47710 63000
rect 48740 63000 48780 63050
rect 47882 62948 48058 62982
rect 48380 62948 48556 62982
rect 47798 62904 47832 62938
rect 48615 62904 48649 62938
rect 47882 62860 48058 62894
rect 48380 62860 48556 62894
rect 47670 62790 47710 62842
rect 47670 62690 47710 62730
rect 47670 62532 47696 62690
rect 47696 62532 47710 62690
rect 48740 62842 48752 63000
rect 48752 62842 48780 63000
rect 48740 62810 48780 62842
rect 48740 62690 48780 62730
rect 47882 62638 48058 62672
rect 48380 62638 48556 62672
rect 47798 62594 47832 62628
rect 48615 62594 48649 62628
rect 47882 62550 48058 62584
rect 48380 62550 48556 62584
rect 47670 62490 47710 62532
rect 48740 62532 48752 62690
rect 48752 62532 48780 62690
rect 48740 62490 48780 62532
rect 52660 63000 52700 63050
rect 52660 62842 52686 63000
rect 52686 62842 52700 63000
rect 53730 63000 53770 63050
rect 52872 62948 53048 62982
rect 53370 62948 53546 62982
rect 52788 62904 52822 62938
rect 53605 62904 53639 62938
rect 52872 62860 53048 62894
rect 53370 62860 53546 62894
rect 52660 62790 52700 62842
rect 52660 62690 52700 62730
rect 52660 62532 52686 62690
rect 52686 62532 52700 62690
rect 53730 62842 53742 63000
rect 53742 62842 53770 63000
rect 53730 62810 53770 62842
rect 53730 62690 53770 62730
rect 52872 62638 53048 62672
rect 53370 62638 53546 62672
rect 52788 62594 52822 62628
rect 53605 62594 53639 62628
rect 52872 62550 53048 62584
rect 53370 62550 53546 62584
rect 52660 62490 52700 62532
rect 53730 62532 53742 62690
rect 53742 62532 53770 62690
rect 53730 62490 53770 62532
rect 57650 63000 57690 63050
rect 57650 62842 57676 63000
rect 57676 62842 57690 63000
rect 58720 63000 58760 63050
rect 57862 62948 58038 62982
rect 58360 62948 58536 62982
rect 57778 62904 57812 62938
rect 58595 62904 58629 62938
rect 57862 62860 58038 62894
rect 58360 62860 58536 62894
rect 57650 62790 57690 62842
rect 57650 62690 57690 62730
rect 57650 62532 57676 62690
rect 57676 62532 57690 62690
rect 58720 62842 58732 63000
rect 58732 62842 58760 63000
rect 58720 62810 58760 62842
rect 58720 62690 58760 62730
rect 57862 62638 58038 62672
rect 58360 62638 58536 62672
rect 57778 62594 57812 62628
rect 58595 62594 58629 62628
rect 57862 62550 58038 62584
rect 58360 62550 58536 62584
rect 57650 62490 57690 62532
rect 58720 62532 58732 62690
rect 58732 62532 58760 62690
rect 58720 62490 58760 62532
rect 62640 63000 62680 63050
rect 62640 62842 62666 63000
rect 62666 62842 62680 63000
rect 63710 63000 63750 63050
rect 62852 62948 63028 62982
rect 63350 62948 63526 62982
rect 62768 62904 62802 62938
rect 63585 62904 63619 62938
rect 62852 62860 63028 62894
rect 63350 62860 63526 62894
rect 62640 62790 62680 62842
rect 62640 62690 62680 62730
rect 62640 62532 62666 62690
rect 62666 62532 62680 62690
rect 63710 62842 63722 63000
rect 63722 62842 63750 63000
rect 63710 62810 63750 62842
rect 63710 62690 63750 62730
rect 62852 62638 63028 62672
rect 63350 62638 63526 62672
rect 62768 62594 62802 62628
rect 63585 62594 63619 62628
rect 62852 62550 63028 62584
rect 63350 62550 63526 62584
rect 62640 62490 62680 62532
rect 63710 62532 63722 62690
rect 63722 62532 63750 62690
rect 63710 62490 63750 62532
rect 67630 63000 67670 63050
rect 67630 62842 67656 63000
rect 67656 62842 67670 63000
rect 68700 63000 68740 63050
rect 67842 62948 68018 62982
rect 68340 62948 68516 62982
rect 67758 62904 67792 62938
rect 68575 62904 68609 62938
rect 67842 62860 68018 62894
rect 68340 62860 68516 62894
rect 67630 62790 67670 62842
rect 67630 62690 67670 62730
rect 67630 62532 67656 62690
rect 67656 62532 67670 62690
rect 68700 62842 68712 63000
rect 68712 62842 68740 63000
rect 68700 62810 68740 62842
rect 68700 62690 68740 62730
rect 67842 62638 68018 62672
rect 68340 62638 68516 62672
rect 67758 62594 67792 62628
rect 68575 62594 68609 62628
rect 67842 62550 68018 62584
rect 68340 62550 68516 62584
rect 67630 62490 67670 62532
rect 68700 62532 68712 62690
rect 68712 62532 68740 62690
rect 68700 62490 68740 62532
rect 72620 63000 72660 63050
rect 72620 62842 72646 63000
rect 72646 62842 72660 63000
rect 73690 63000 73730 63050
rect 72832 62948 73008 62982
rect 73330 62948 73506 62982
rect 72748 62904 72782 62938
rect 73565 62904 73599 62938
rect 72832 62860 73008 62894
rect 73330 62860 73506 62894
rect 72620 62790 72660 62842
rect 72620 62690 72660 62730
rect 72620 62532 72646 62690
rect 72646 62532 72660 62690
rect 73690 62842 73702 63000
rect 73702 62842 73730 63000
rect 73690 62810 73730 62842
rect 73690 62690 73730 62730
rect 72832 62638 73008 62672
rect 73330 62638 73506 62672
rect 72748 62594 72782 62628
rect 73565 62594 73599 62628
rect 72832 62550 73008 62584
rect 73330 62550 73506 62584
rect 72620 62490 72660 62532
rect 73690 62532 73702 62690
rect 73702 62532 73730 62690
rect 73690 62490 73730 62532
rect 77610 63000 77650 63050
rect 77610 62842 77636 63000
rect 77636 62842 77650 63000
rect 78680 63000 78720 63050
rect 77822 62948 77998 62982
rect 78320 62948 78496 62982
rect 77738 62904 77772 62938
rect 78555 62904 78589 62938
rect 77822 62860 77998 62894
rect 78320 62860 78496 62894
rect 77610 62790 77650 62842
rect 77610 62690 77650 62730
rect 77610 62532 77636 62690
rect 77636 62532 77650 62690
rect 78680 62842 78692 63000
rect 78692 62842 78720 63000
rect 78680 62810 78720 62842
rect 78680 62690 78720 62730
rect 77822 62638 77998 62672
rect 78320 62638 78496 62672
rect 77738 62594 77772 62628
rect 78555 62594 78589 62628
rect 77822 62550 77998 62584
rect 78320 62550 78496 62584
rect 77610 62490 77650 62532
rect 78680 62532 78692 62690
rect 78692 62532 78720 62690
rect 78680 62490 78720 62532
rect 2760 61290 2800 61340
rect 2760 61132 2786 61290
rect 2786 61132 2800 61290
rect 3830 61290 3870 61340
rect 2972 61238 3148 61272
rect 3470 61238 3646 61272
rect 2888 61194 2922 61228
rect 3705 61194 3739 61228
rect 2972 61150 3148 61184
rect 3470 61150 3646 61184
rect 2760 61080 2800 61132
rect 2760 60980 2800 61020
rect 2760 60822 2786 60980
rect 2786 60822 2800 60980
rect 3830 61132 3842 61290
rect 3842 61132 3870 61290
rect 3830 61100 3870 61132
rect 3830 60980 3870 61020
rect 2972 60928 3148 60962
rect 3470 60928 3646 60962
rect 2888 60884 2922 60918
rect 3705 60884 3739 60918
rect 2972 60840 3148 60874
rect 3470 60840 3646 60874
rect 2760 60780 2800 60822
rect 3830 60822 3842 60980
rect 3842 60822 3870 60980
rect 3830 60780 3870 60822
rect 7750 61290 7790 61340
rect 7750 61132 7776 61290
rect 7776 61132 7790 61290
rect 8820 61290 8860 61340
rect 7962 61238 8138 61272
rect 8460 61238 8636 61272
rect 7878 61194 7912 61228
rect 8695 61194 8729 61228
rect 7962 61150 8138 61184
rect 8460 61150 8636 61184
rect 7750 61080 7790 61132
rect 7750 60980 7790 61020
rect 7750 60822 7776 60980
rect 7776 60822 7790 60980
rect 8820 61132 8832 61290
rect 8832 61132 8860 61290
rect 8820 61100 8860 61132
rect 8820 60980 8860 61020
rect 7962 60928 8138 60962
rect 8460 60928 8636 60962
rect 7878 60884 7912 60918
rect 8695 60884 8729 60918
rect 7962 60840 8138 60874
rect 8460 60840 8636 60874
rect 7750 60780 7790 60822
rect 8820 60822 8832 60980
rect 8832 60822 8860 60980
rect 8820 60780 8860 60822
rect 12740 61290 12780 61340
rect 12740 61132 12766 61290
rect 12766 61132 12780 61290
rect 13810 61290 13850 61340
rect 12952 61238 13128 61272
rect 13450 61238 13626 61272
rect 12868 61194 12902 61228
rect 13685 61194 13719 61228
rect 12952 61150 13128 61184
rect 13450 61150 13626 61184
rect 12740 61080 12780 61132
rect 12740 60980 12780 61020
rect 12740 60822 12766 60980
rect 12766 60822 12780 60980
rect 13810 61132 13822 61290
rect 13822 61132 13850 61290
rect 13810 61100 13850 61132
rect 13810 60980 13850 61020
rect 12952 60928 13128 60962
rect 13450 60928 13626 60962
rect 12868 60884 12902 60918
rect 13685 60884 13719 60918
rect 12952 60840 13128 60874
rect 13450 60840 13626 60874
rect 12740 60780 12780 60822
rect 13810 60822 13822 60980
rect 13822 60822 13850 60980
rect 13810 60780 13850 60822
rect 17730 61290 17770 61340
rect 17730 61132 17756 61290
rect 17756 61132 17770 61290
rect 18800 61290 18840 61340
rect 17942 61238 18118 61272
rect 18440 61238 18616 61272
rect 17858 61194 17892 61228
rect 18675 61194 18709 61228
rect 17942 61150 18118 61184
rect 18440 61150 18616 61184
rect 17730 61080 17770 61132
rect 17730 60980 17770 61020
rect 17730 60822 17756 60980
rect 17756 60822 17770 60980
rect 18800 61132 18812 61290
rect 18812 61132 18840 61290
rect 18800 61100 18840 61132
rect 18800 60980 18840 61020
rect 17942 60928 18118 60962
rect 18440 60928 18616 60962
rect 17858 60884 17892 60918
rect 18675 60884 18709 60918
rect 17942 60840 18118 60874
rect 18440 60840 18616 60874
rect 17730 60780 17770 60822
rect 18800 60822 18812 60980
rect 18812 60822 18840 60980
rect 18800 60780 18840 60822
rect 22720 61290 22760 61340
rect 22720 61132 22746 61290
rect 22746 61132 22760 61290
rect 23790 61290 23830 61340
rect 22932 61238 23108 61272
rect 23430 61238 23606 61272
rect 22848 61194 22882 61228
rect 23665 61194 23699 61228
rect 22932 61150 23108 61184
rect 23430 61150 23606 61184
rect 22720 61080 22760 61132
rect 22720 60980 22760 61020
rect 22720 60822 22746 60980
rect 22746 60822 22760 60980
rect 23790 61132 23802 61290
rect 23802 61132 23830 61290
rect 23790 61100 23830 61132
rect 23790 60980 23830 61020
rect 22932 60928 23108 60962
rect 23430 60928 23606 60962
rect 22848 60884 22882 60918
rect 23665 60884 23699 60918
rect 22932 60840 23108 60874
rect 23430 60840 23606 60874
rect 22720 60780 22760 60822
rect 23790 60822 23802 60980
rect 23802 60822 23830 60980
rect 23790 60780 23830 60822
rect 27710 61290 27750 61340
rect 27710 61132 27736 61290
rect 27736 61132 27750 61290
rect 28780 61290 28820 61340
rect 27922 61238 28098 61272
rect 28420 61238 28596 61272
rect 27838 61194 27872 61228
rect 28655 61194 28689 61228
rect 27922 61150 28098 61184
rect 28420 61150 28596 61184
rect 27710 61080 27750 61132
rect 27710 60980 27750 61020
rect 27710 60822 27736 60980
rect 27736 60822 27750 60980
rect 28780 61132 28792 61290
rect 28792 61132 28820 61290
rect 28780 61100 28820 61132
rect 28780 60980 28820 61020
rect 27922 60928 28098 60962
rect 28420 60928 28596 60962
rect 27838 60884 27872 60918
rect 28655 60884 28689 60918
rect 27922 60840 28098 60874
rect 28420 60840 28596 60874
rect 27710 60780 27750 60822
rect 28780 60822 28792 60980
rect 28792 60822 28820 60980
rect 28780 60780 28820 60822
rect 32700 61290 32740 61340
rect 32700 61132 32726 61290
rect 32726 61132 32740 61290
rect 33770 61290 33810 61340
rect 32912 61238 33088 61272
rect 33410 61238 33586 61272
rect 32828 61194 32862 61228
rect 33645 61194 33679 61228
rect 32912 61150 33088 61184
rect 33410 61150 33586 61184
rect 32700 61080 32740 61132
rect 32700 60980 32740 61020
rect 32700 60822 32726 60980
rect 32726 60822 32740 60980
rect 33770 61132 33782 61290
rect 33782 61132 33810 61290
rect 33770 61100 33810 61132
rect 33770 60980 33810 61020
rect 32912 60928 33088 60962
rect 33410 60928 33586 60962
rect 32828 60884 32862 60918
rect 33645 60884 33679 60918
rect 32912 60840 33088 60874
rect 33410 60840 33586 60874
rect 32700 60780 32740 60822
rect 33770 60822 33782 60980
rect 33782 60822 33810 60980
rect 33770 60780 33810 60822
rect 37690 61290 37730 61340
rect 37690 61132 37716 61290
rect 37716 61132 37730 61290
rect 38760 61290 38800 61340
rect 37902 61238 38078 61272
rect 38400 61238 38576 61272
rect 37818 61194 37852 61228
rect 38635 61194 38669 61228
rect 37902 61150 38078 61184
rect 38400 61150 38576 61184
rect 37690 61080 37730 61132
rect 37690 60980 37730 61020
rect 37690 60822 37716 60980
rect 37716 60822 37730 60980
rect 38760 61132 38772 61290
rect 38772 61132 38800 61290
rect 38760 61100 38800 61132
rect 38760 60980 38800 61020
rect 37902 60928 38078 60962
rect 38400 60928 38576 60962
rect 37818 60884 37852 60918
rect 38635 60884 38669 60918
rect 37902 60840 38078 60874
rect 38400 60840 38576 60874
rect 37690 60780 37730 60822
rect 38760 60822 38772 60980
rect 38772 60822 38800 60980
rect 38760 60780 38800 60822
rect 42680 61290 42720 61340
rect 42680 61132 42706 61290
rect 42706 61132 42720 61290
rect 43750 61290 43790 61340
rect 42892 61238 43068 61272
rect 43390 61238 43566 61272
rect 42808 61194 42842 61228
rect 43625 61194 43659 61228
rect 42892 61150 43068 61184
rect 43390 61150 43566 61184
rect 42680 61080 42720 61132
rect 42680 60980 42720 61020
rect 42680 60822 42706 60980
rect 42706 60822 42720 60980
rect 43750 61132 43762 61290
rect 43762 61132 43790 61290
rect 43750 61100 43790 61132
rect 43750 60980 43790 61020
rect 42892 60928 43068 60962
rect 43390 60928 43566 60962
rect 42808 60884 42842 60918
rect 43625 60884 43659 60918
rect 42892 60840 43068 60874
rect 43390 60840 43566 60874
rect 42680 60780 42720 60822
rect 43750 60822 43762 60980
rect 43762 60822 43790 60980
rect 43750 60780 43790 60822
rect 47670 61290 47710 61340
rect 47670 61132 47696 61290
rect 47696 61132 47710 61290
rect 48740 61290 48780 61340
rect 47882 61238 48058 61272
rect 48380 61238 48556 61272
rect 47798 61194 47832 61228
rect 48615 61194 48649 61228
rect 47882 61150 48058 61184
rect 48380 61150 48556 61184
rect 47670 61080 47710 61132
rect 47670 60980 47710 61020
rect 47670 60822 47696 60980
rect 47696 60822 47710 60980
rect 48740 61132 48752 61290
rect 48752 61132 48780 61290
rect 48740 61100 48780 61132
rect 48740 60980 48780 61020
rect 47882 60928 48058 60962
rect 48380 60928 48556 60962
rect 47798 60884 47832 60918
rect 48615 60884 48649 60918
rect 47882 60840 48058 60874
rect 48380 60840 48556 60874
rect 47670 60780 47710 60822
rect 48740 60822 48752 60980
rect 48752 60822 48780 60980
rect 48740 60780 48780 60822
rect 52660 61290 52700 61340
rect 52660 61132 52686 61290
rect 52686 61132 52700 61290
rect 53730 61290 53770 61340
rect 52872 61238 53048 61272
rect 53370 61238 53546 61272
rect 52788 61194 52822 61228
rect 53605 61194 53639 61228
rect 52872 61150 53048 61184
rect 53370 61150 53546 61184
rect 52660 61080 52700 61132
rect 52660 60980 52700 61020
rect 52660 60822 52686 60980
rect 52686 60822 52700 60980
rect 53730 61132 53742 61290
rect 53742 61132 53770 61290
rect 53730 61100 53770 61132
rect 53730 60980 53770 61020
rect 52872 60928 53048 60962
rect 53370 60928 53546 60962
rect 52788 60884 52822 60918
rect 53605 60884 53639 60918
rect 52872 60840 53048 60874
rect 53370 60840 53546 60874
rect 52660 60780 52700 60822
rect 53730 60822 53742 60980
rect 53742 60822 53770 60980
rect 53730 60780 53770 60822
rect 57650 61290 57690 61340
rect 57650 61132 57676 61290
rect 57676 61132 57690 61290
rect 58720 61290 58760 61340
rect 57862 61238 58038 61272
rect 58360 61238 58536 61272
rect 57778 61194 57812 61228
rect 58595 61194 58629 61228
rect 57862 61150 58038 61184
rect 58360 61150 58536 61184
rect 57650 61080 57690 61132
rect 57650 60980 57690 61020
rect 57650 60822 57676 60980
rect 57676 60822 57690 60980
rect 58720 61132 58732 61290
rect 58732 61132 58760 61290
rect 58720 61100 58760 61132
rect 58720 60980 58760 61020
rect 57862 60928 58038 60962
rect 58360 60928 58536 60962
rect 57778 60884 57812 60918
rect 58595 60884 58629 60918
rect 57862 60840 58038 60874
rect 58360 60840 58536 60874
rect 57650 60780 57690 60822
rect 58720 60822 58732 60980
rect 58732 60822 58760 60980
rect 58720 60780 58760 60822
rect 62640 61290 62680 61340
rect 62640 61132 62666 61290
rect 62666 61132 62680 61290
rect 63710 61290 63750 61340
rect 62852 61238 63028 61272
rect 63350 61238 63526 61272
rect 62768 61194 62802 61228
rect 63585 61194 63619 61228
rect 62852 61150 63028 61184
rect 63350 61150 63526 61184
rect 62640 61080 62680 61132
rect 62640 60980 62680 61020
rect 62640 60822 62666 60980
rect 62666 60822 62680 60980
rect 63710 61132 63722 61290
rect 63722 61132 63750 61290
rect 63710 61100 63750 61132
rect 63710 60980 63750 61020
rect 62852 60928 63028 60962
rect 63350 60928 63526 60962
rect 62768 60884 62802 60918
rect 63585 60884 63619 60918
rect 62852 60840 63028 60874
rect 63350 60840 63526 60874
rect 62640 60780 62680 60822
rect 63710 60822 63722 60980
rect 63722 60822 63750 60980
rect 63710 60780 63750 60822
rect 67630 61290 67670 61340
rect 67630 61132 67656 61290
rect 67656 61132 67670 61290
rect 68700 61290 68740 61340
rect 67842 61238 68018 61272
rect 68340 61238 68516 61272
rect 67758 61194 67792 61228
rect 68575 61194 68609 61228
rect 67842 61150 68018 61184
rect 68340 61150 68516 61184
rect 67630 61080 67670 61132
rect 67630 60980 67670 61020
rect 67630 60822 67656 60980
rect 67656 60822 67670 60980
rect 68700 61132 68712 61290
rect 68712 61132 68740 61290
rect 68700 61100 68740 61132
rect 68700 60980 68740 61020
rect 67842 60928 68018 60962
rect 68340 60928 68516 60962
rect 67758 60884 67792 60918
rect 68575 60884 68609 60918
rect 67842 60840 68018 60874
rect 68340 60840 68516 60874
rect 67630 60780 67670 60822
rect 68700 60822 68712 60980
rect 68712 60822 68740 60980
rect 68700 60780 68740 60822
rect 72620 61290 72660 61340
rect 72620 61132 72646 61290
rect 72646 61132 72660 61290
rect 73690 61290 73730 61340
rect 72832 61238 73008 61272
rect 73330 61238 73506 61272
rect 72748 61194 72782 61228
rect 73565 61194 73599 61228
rect 72832 61150 73008 61184
rect 73330 61150 73506 61184
rect 72620 61080 72660 61132
rect 72620 60980 72660 61020
rect 72620 60822 72646 60980
rect 72646 60822 72660 60980
rect 73690 61132 73702 61290
rect 73702 61132 73730 61290
rect 73690 61100 73730 61132
rect 73690 60980 73730 61020
rect 72832 60928 73008 60962
rect 73330 60928 73506 60962
rect 72748 60884 72782 60918
rect 73565 60884 73599 60918
rect 72832 60840 73008 60874
rect 73330 60840 73506 60874
rect 72620 60780 72660 60822
rect 73690 60822 73702 60980
rect 73702 60822 73730 60980
rect 73690 60780 73730 60822
rect 77610 61290 77650 61340
rect 77610 61132 77636 61290
rect 77636 61132 77650 61290
rect 78680 61290 78720 61340
rect 77822 61238 77998 61272
rect 78320 61238 78496 61272
rect 77738 61194 77772 61228
rect 78555 61194 78589 61228
rect 77822 61150 77998 61184
rect 78320 61150 78496 61184
rect 77610 61080 77650 61132
rect 77610 60980 77650 61020
rect 77610 60822 77636 60980
rect 77636 60822 77650 60980
rect 78680 61132 78692 61290
rect 78692 61132 78720 61290
rect 78680 61100 78720 61132
rect 78680 60980 78720 61020
rect 77822 60928 77998 60962
rect 78320 60928 78496 60962
rect 77738 60884 77772 60918
rect 78555 60884 78589 60918
rect 77822 60840 77998 60874
rect 78320 60840 78496 60874
rect 77610 60780 77650 60822
rect 78680 60822 78692 60980
rect 78692 60822 78720 60980
rect 78680 60780 78720 60822
rect 2760 59580 2800 59630
rect 2760 59422 2786 59580
rect 2786 59422 2800 59580
rect 3830 59580 3870 59630
rect 2972 59528 3148 59562
rect 3470 59528 3646 59562
rect 2888 59484 2922 59518
rect 3705 59484 3739 59518
rect 2972 59440 3148 59474
rect 3470 59440 3646 59474
rect 2760 59370 2800 59422
rect 2760 59270 2800 59310
rect 2760 59112 2786 59270
rect 2786 59112 2800 59270
rect 3830 59422 3842 59580
rect 3842 59422 3870 59580
rect 3830 59390 3870 59422
rect 3830 59270 3870 59310
rect 2972 59218 3148 59252
rect 3470 59218 3646 59252
rect 2888 59174 2922 59208
rect 3705 59174 3739 59208
rect 2972 59130 3148 59164
rect 3470 59130 3646 59164
rect 2760 59070 2800 59112
rect 3830 59112 3842 59270
rect 3842 59112 3870 59270
rect 3830 59070 3870 59112
rect 7750 59580 7790 59630
rect 7750 59422 7776 59580
rect 7776 59422 7790 59580
rect 8820 59580 8860 59630
rect 7962 59528 8138 59562
rect 8460 59528 8636 59562
rect 7878 59484 7912 59518
rect 8695 59484 8729 59518
rect 7962 59440 8138 59474
rect 8460 59440 8636 59474
rect 7750 59370 7790 59422
rect 7750 59270 7790 59310
rect 7750 59112 7776 59270
rect 7776 59112 7790 59270
rect 8820 59422 8832 59580
rect 8832 59422 8860 59580
rect 8820 59390 8860 59422
rect 8820 59270 8860 59310
rect 7962 59218 8138 59252
rect 8460 59218 8636 59252
rect 7878 59174 7912 59208
rect 8695 59174 8729 59208
rect 7962 59130 8138 59164
rect 8460 59130 8636 59164
rect 7750 59070 7790 59112
rect 8820 59112 8832 59270
rect 8832 59112 8860 59270
rect 8820 59070 8860 59112
rect 12740 59580 12780 59630
rect 12740 59422 12766 59580
rect 12766 59422 12780 59580
rect 13810 59580 13850 59630
rect 12952 59528 13128 59562
rect 13450 59528 13626 59562
rect 12868 59484 12902 59518
rect 13685 59484 13719 59518
rect 12952 59440 13128 59474
rect 13450 59440 13626 59474
rect 12740 59370 12780 59422
rect 12740 59270 12780 59310
rect 12740 59112 12766 59270
rect 12766 59112 12780 59270
rect 13810 59422 13822 59580
rect 13822 59422 13850 59580
rect 13810 59390 13850 59422
rect 13810 59270 13850 59310
rect 12952 59218 13128 59252
rect 13450 59218 13626 59252
rect 12868 59174 12902 59208
rect 13685 59174 13719 59208
rect 12952 59130 13128 59164
rect 13450 59130 13626 59164
rect 12740 59070 12780 59112
rect 13810 59112 13822 59270
rect 13822 59112 13850 59270
rect 13810 59070 13850 59112
rect 17730 59580 17770 59630
rect 17730 59422 17756 59580
rect 17756 59422 17770 59580
rect 18800 59580 18840 59630
rect 17942 59528 18118 59562
rect 18440 59528 18616 59562
rect 17858 59484 17892 59518
rect 18675 59484 18709 59518
rect 17942 59440 18118 59474
rect 18440 59440 18616 59474
rect 17730 59370 17770 59422
rect 17730 59270 17770 59310
rect 17730 59112 17756 59270
rect 17756 59112 17770 59270
rect 18800 59422 18812 59580
rect 18812 59422 18840 59580
rect 18800 59390 18840 59422
rect 18800 59270 18840 59310
rect 17942 59218 18118 59252
rect 18440 59218 18616 59252
rect 17858 59174 17892 59208
rect 18675 59174 18709 59208
rect 17942 59130 18118 59164
rect 18440 59130 18616 59164
rect 17730 59070 17770 59112
rect 18800 59112 18812 59270
rect 18812 59112 18840 59270
rect 18800 59070 18840 59112
rect 22720 59580 22760 59630
rect 22720 59422 22746 59580
rect 22746 59422 22760 59580
rect 23790 59580 23830 59630
rect 22932 59528 23108 59562
rect 23430 59528 23606 59562
rect 22848 59484 22882 59518
rect 23665 59484 23699 59518
rect 22932 59440 23108 59474
rect 23430 59440 23606 59474
rect 22720 59370 22760 59422
rect 22720 59270 22760 59310
rect 22720 59112 22746 59270
rect 22746 59112 22760 59270
rect 23790 59422 23802 59580
rect 23802 59422 23830 59580
rect 23790 59390 23830 59422
rect 23790 59270 23830 59310
rect 22932 59218 23108 59252
rect 23430 59218 23606 59252
rect 22848 59174 22882 59208
rect 23665 59174 23699 59208
rect 22932 59130 23108 59164
rect 23430 59130 23606 59164
rect 22720 59070 22760 59112
rect 23790 59112 23802 59270
rect 23802 59112 23830 59270
rect 23790 59070 23830 59112
rect 27710 59580 27750 59630
rect 27710 59422 27736 59580
rect 27736 59422 27750 59580
rect 28780 59580 28820 59630
rect 27922 59528 28098 59562
rect 28420 59528 28596 59562
rect 27838 59484 27872 59518
rect 28655 59484 28689 59518
rect 27922 59440 28098 59474
rect 28420 59440 28596 59474
rect 27710 59370 27750 59422
rect 27710 59270 27750 59310
rect 27710 59112 27736 59270
rect 27736 59112 27750 59270
rect 28780 59422 28792 59580
rect 28792 59422 28820 59580
rect 28780 59390 28820 59422
rect 28780 59270 28820 59310
rect 27922 59218 28098 59252
rect 28420 59218 28596 59252
rect 27838 59174 27872 59208
rect 28655 59174 28689 59208
rect 27922 59130 28098 59164
rect 28420 59130 28596 59164
rect 27710 59070 27750 59112
rect 28780 59112 28792 59270
rect 28792 59112 28820 59270
rect 28780 59070 28820 59112
rect 32700 59580 32740 59630
rect 32700 59422 32726 59580
rect 32726 59422 32740 59580
rect 33770 59580 33810 59630
rect 32912 59528 33088 59562
rect 33410 59528 33586 59562
rect 32828 59484 32862 59518
rect 33645 59484 33679 59518
rect 32912 59440 33088 59474
rect 33410 59440 33586 59474
rect 32700 59370 32740 59422
rect 32700 59270 32740 59310
rect 32700 59112 32726 59270
rect 32726 59112 32740 59270
rect 33770 59422 33782 59580
rect 33782 59422 33810 59580
rect 33770 59390 33810 59422
rect 33770 59270 33810 59310
rect 32912 59218 33088 59252
rect 33410 59218 33586 59252
rect 32828 59174 32862 59208
rect 33645 59174 33679 59208
rect 32912 59130 33088 59164
rect 33410 59130 33586 59164
rect 32700 59070 32740 59112
rect 33770 59112 33782 59270
rect 33782 59112 33810 59270
rect 33770 59070 33810 59112
rect 37690 59580 37730 59630
rect 37690 59422 37716 59580
rect 37716 59422 37730 59580
rect 38760 59580 38800 59630
rect 37902 59528 38078 59562
rect 38400 59528 38576 59562
rect 37818 59484 37852 59518
rect 38635 59484 38669 59518
rect 37902 59440 38078 59474
rect 38400 59440 38576 59474
rect 37690 59370 37730 59422
rect 37690 59270 37730 59310
rect 37690 59112 37716 59270
rect 37716 59112 37730 59270
rect 38760 59422 38772 59580
rect 38772 59422 38800 59580
rect 38760 59390 38800 59422
rect 38760 59270 38800 59310
rect 37902 59218 38078 59252
rect 38400 59218 38576 59252
rect 37818 59174 37852 59208
rect 38635 59174 38669 59208
rect 37902 59130 38078 59164
rect 38400 59130 38576 59164
rect 37690 59070 37730 59112
rect 38760 59112 38772 59270
rect 38772 59112 38800 59270
rect 38760 59070 38800 59112
rect 42680 59580 42720 59630
rect 42680 59422 42706 59580
rect 42706 59422 42720 59580
rect 43750 59580 43790 59630
rect 42892 59528 43068 59562
rect 43390 59528 43566 59562
rect 42808 59484 42842 59518
rect 43625 59484 43659 59518
rect 42892 59440 43068 59474
rect 43390 59440 43566 59474
rect 42680 59370 42720 59422
rect 42680 59270 42720 59310
rect 42680 59112 42706 59270
rect 42706 59112 42720 59270
rect 43750 59422 43762 59580
rect 43762 59422 43790 59580
rect 43750 59390 43790 59422
rect 43750 59270 43790 59310
rect 42892 59218 43068 59252
rect 43390 59218 43566 59252
rect 42808 59174 42842 59208
rect 43625 59174 43659 59208
rect 42892 59130 43068 59164
rect 43390 59130 43566 59164
rect 42680 59070 42720 59112
rect 43750 59112 43762 59270
rect 43762 59112 43790 59270
rect 43750 59070 43790 59112
rect 47670 59580 47710 59630
rect 47670 59422 47696 59580
rect 47696 59422 47710 59580
rect 48740 59580 48780 59630
rect 47882 59528 48058 59562
rect 48380 59528 48556 59562
rect 47798 59484 47832 59518
rect 48615 59484 48649 59518
rect 47882 59440 48058 59474
rect 48380 59440 48556 59474
rect 47670 59370 47710 59422
rect 47670 59270 47710 59310
rect 47670 59112 47696 59270
rect 47696 59112 47710 59270
rect 48740 59422 48752 59580
rect 48752 59422 48780 59580
rect 48740 59390 48780 59422
rect 48740 59270 48780 59310
rect 47882 59218 48058 59252
rect 48380 59218 48556 59252
rect 47798 59174 47832 59208
rect 48615 59174 48649 59208
rect 47882 59130 48058 59164
rect 48380 59130 48556 59164
rect 47670 59070 47710 59112
rect 48740 59112 48752 59270
rect 48752 59112 48780 59270
rect 48740 59070 48780 59112
rect 52660 59580 52700 59630
rect 52660 59422 52686 59580
rect 52686 59422 52700 59580
rect 53730 59580 53770 59630
rect 52872 59528 53048 59562
rect 53370 59528 53546 59562
rect 52788 59484 52822 59518
rect 53605 59484 53639 59518
rect 52872 59440 53048 59474
rect 53370 59440 53546 59474
rect 52660 59370 52700 59422
rect 52660 59270 52700 59310
rect 52660 59112 52686 59270
rect 52686 59112 52700 59270
rect 53730 59422 53742 59580
rect 53742 59422 53770 59580
rect 53730 59390 53770 59422
rect 53730 59270 53770 59310
rect 52872 59218 53048 59252
rect 53370 59218 53546 59252
rect 52788 59174 52822 59208
rect 53605 59174 53639 59208
rect 52872 59130 53048 59164
rect 53370 59130 53546 59164
rect 52660 59070 52700 59112
rect 53730 59112 53742 59270
rect 53742 59112 53770 59270
rect 53730 59070 53770 59112
rect 57650 59580 57690 59630
rect 57650 59422 57676 59580
rect 57676 59422 57690 59580
rect 58720 59580 58760 59630
rect 57862 59528 58038 59562
rect 58360 59528 58536 59562
rect 57778 59484 57812 59518
rect 58595 59484 58629 59518
rect 57862 59440 58038 59474
rect 58360 59440 58536 59474
rect 57650 59370 57690 59422
rect 57650 59270 57690 59310
rect 57650 59112 57676 59270
rect 57676 59112 57690 59270
rect 58720 59422 58732 59580
rect 58732 59422 58760 59580
rect 58720 59390 58760 59422
rect 58720 59270 58760 59310
rect 57862 59218 58038 59252
rect 58360 59218 58536 59252
rect 57778 59174 57812 59208
rect 58595 59174 58629 59208
rect 57862 59130 58038 59164
rect 58360 59130 58536 59164
rect 57650 59070 57690 59112
rect 58720 59112 58732 59270
rect 58732 59112 58760 59270
rect 58720 59070 58760 59112
rect 62640 59580 62680 59630
rect 62640 59422 62666 59580
rect 62666 59422 62680 59580
rect 63710 59580 63750 59630
rect 62852 59528 63028 59562
rect 63350 59528 63526 59562
rect 62768 59484 62802 59518
rect 63585 59484 63619 59518
rect 62852 59440 63028 59474
rect 63350 59440 63526 59474
rect 62640 59370 62680 59422
rect 62640 59270 62680 59310
rect 62640 59112 62666 59270
rect 62666 59112 62680 59270
rect 63710 59422 63722 59580
rect 63722 59422 63750 59580
rect 63710 59390 63750 59422
rect 63710 59270 63750 59310
rect 62852 59218 63028 59252
rect 63350 59218 63526 59252
rect 62768 59174 62802 59208
rect 63585 59174 63619 59208
rect 62852 59130 63028 59164
rect 63350 59130 63526 59164
rect 62640 59070 62680 59112
rect 63710 59112 63722 59270
rect 63722 59112 63750 59270
rect 63710 59070 63750 59112
rect 67630 59580 67670 59630
rect 67630 59422 67656 59580
rect 67656 59422 67670 59580
rect 68700 59580 68740 59630
rect 67842 59528 68018 59562
rect 68340 59528 68516 59562
rect 67758 59484 67792 59518
rect 68575 59484 68609 59518
rect 67842 59440 68018 59474
rect 68340 59440 68516 59474
rect 67630 59370 67670 59422
rect 67630 59270 67670 59310
rect 67630 59112 67656 59270
rect 67656 59112 67670 59270
rect 68700 59422 68712 59580
rect 68712 59422 68740 59580
rect 68700 59390 68740 59422
rect 68700 59270 68740 59310
rect 67842 59218 68018 59252
rect 68340 59218 68516 59252
rect 67758 59174 67792 59208
rect 68575 59174 68609 59208
rect 67842 59130 68018 59164
rect 68340 59130 68516 59164
rect 67630 59070 67670 59112
rect 68700 59112 68712 59270
rect 68712 59112 68740 59270
rect 68700 59070 68740 59112
rect 72620 59580 72660 59630
rect 72620 59422 72646 59580
rect 72646 59422 72660 59580
rect 73690 59580 73730 59630
rect 72832 59528 73008 59562
rect 73330 59528 73506 59562
rect 72748 59484 72782 59518
rect 73565 59484 73599 59518
rect 72832 59440 73008 59474
rect 73330 59440 73506 59474
rect 72620 59370 72660 59422
rect 72620 59270 72660 59310
rect 72620 59112 72646 59270
rect 72646 59112 72660 59270
rect 73690 59422 73702 59580
rect 73702 59422 73730 59580
rect 73690 59390 73730 59422
rect 73690 59270 73730 59310
rect 72832 59218 73008 59252
rect 73330 59218 73506 59252
rect 72748 59174 72782 59208
rect 73565 59174 73599 59208
rect 72832 59130 73008 59164
rect 73330 59130 73506 59164
rect 72620 59070 72660 59112
rect 73690 59112 73702 59270
rect 73702 59112 73730 59270
rect 73690 59070 73730 59112
rect 77610 59580 77650 59630
rect 77610 59422 77636 59580
rect 77636 59422 77650 59580
rect 78680 59580 78720 59630
rect 77822 59528 77998 59562
rect 78320 59528 78496 59562
rect 77738 59484 77772 59518
rect 78555 59484 78589 59518
rect 77822 59440 77998 59474
rect 78320 59440 78496 59474
rect 77610 59370 77650 59422
rect 77610 59270 77650 59310
rect 77610 59112 77636 59270
rect 77636 59112 77650 59270
rect 78680 59422 78692 59580
rect 78692 59422 78720 59580
rect 78680 59390 78720 59422
rect 78680 59270 78720 59310
rect 77822 59218 77998 59252
rect 78320 59218 78496 59252
rect 77738 59174 77772 59208
rect 78555 59174 78589 59208
rect 77822 59130 77998 59164
rect 78320 59130 78496 59164
rect 77610 59070 77650 59112
rect 78680 59112 78692 59270
rect 78692 59112 78720 59270
rect 78680 59070 78720 59112
rect 2760 57870 2800 57920
rect 2760 57712 2786 57870
rect 2786 57712 2800 57870
rect 3830 57870 3870 57920
rect 2972 57818 3148 57852
rect 3470 57818 3646 57852
rect 2888 57774 2922 57808
rect 3705 57774 3739 57808
rect 2972 57730 3148 57764
rect 3470 57730 3646 57764
rect 2760 57660 2800 57712
rect 2760 57560 2800 57600
rect 2760 57402 2786 57560
rect 2786 57402 2800 57560
rect 3830 57712 3842 57870
rect 3842 57712 3870 57870
rect 3830 57680 3870 57712
rect 3830 57560 3870 57600
rect 2972 57508 3148 57542
rect 3470 57508 3646 57542
rect 2888 57464 2922 57498
rect 3705 57464 3739 57498
rect 2972 57420 3148 57454
rect 3470 57420 3646 57454
rect 2760 57360 2800 57402
rect 3830 57402 3842 57560
rect 3842 57402 3870 57560
rect 3830 57360 3870 57402
rect 7750 57870 7790 57920
rect 7750 57712 7776 57870
rect 7776 57712 7790 57870
rect 8820 57870 8860 57920
rect 7962 57818 8138 57852
rect 8460 57818 8636 57852
rect 7878 57774 7912 57808
rect 8695 57774 8729 57808
rect 7962 57730 8138 57764
rect 8460 57730 8636 57764
rect 7750 57660 7790 57712
rect 7750 57560 7790 57600
rect 7750 57402 7776 57560
rect 7776 57402 7790 57560
rect 8820 57712 8832 57870
rect 8832 57712 8860 57870
rect 8820 57680 8860 57712
rect 8820 57560 8860 57600
rect 7962 57508 8138 57542
rect 8460 57508 8636 57542
rect 7878 57464 7912 57498
rect 8695 57464 8729 57498
rect 7962 57420 8138 57454
rect 8460 57420 8636 57454
rect 7750 57360 7790 57402
rect 8820 57402 8832 57560
rect 8832 57402 8860 57560
rect 8820 57360 8860 57402
rect 12740 57870 12780 57920
rect 12740 57712 12766 57870
rect 12766 57712 12780 57870
rect 13810 57870 13850 57920
rect 12952 57818 13128 57852
rect 13450 57818 13626 57852
rect 12868 57774 12902 57808
rect 13685 57774 13719 57808
rect 12952 57730 13128 57764
rect 13450 57730 13626 57764
rect 12740 57660 12780 57712
rect 12740 57560 12780 57600
rect 12740 57402 12766 57560
rect 12766 57402 12780 57560
rect 13810 57712 13822 57870
rect 13822 57712 13850 57870
rect 13810 57680 13850 57712
rect 13810 57560 13850 57600
rect 12952 57508 13128 57542
rect 13450 57508 13626 57542
rect 12868 57464 12902 57498
rect 13685 57464 13719 57498
rect 12952 57420 13128 57454
rect 13450 57420 13626 57454
rect 12740 57360 12780 57402
rect 13810 57402 13822 57560
rect 13822 57402 13850 57560
rect 13810 57360 13850 57402
rect 17730 57870 17770 57920
rect 17730 57712 17756 57870
rect 17756 57712 17770 57870
rect 18800 57870 18840 57920
rect 17942 57818 18118 57852
rect 18440 57818 18616 57852
rect 17858 57774 17892 57808
rect 18675 57774 18709 57808
rect 17942 57730 18118 57764
rect 18440 57730 18616 57764
rect 17730 57660 17770 57712
rect 17730 57560 17770 57600
rect 17730 57402 17756 57560
rect 17756 57402 17770 57560
rect 18800 57712 18812 57870
rect 18812 57712 18840 57870
rect 18800 57680 18840 57712
rect 18800 57560 18840 57600
rect 17942 57508 18118 57542
rect 18440 57508 18616 57542
rect 17858 57464 17892 57498
rect 18675 57464 18709 57498
rect 17942 57420 18118 57454
rect 18440 57420 18616 57454
rect 17730 57360 17770 57402
rect 18800 57402 18812 57560
rect 18812 57402 18840 57560
rect 18800 57360 18840 57402
rect 22720 57870 22760 57920
rect 22720 57712 22746 57870
rect 22746 57712 22760 57870
rect 23790 57870 23830 57920
rect 22932 57818 23108 57852
rect 23430 57818 23606 57852
rect 22848 57774 22882 57808
rect 23665 57774 23699 57808
rect 22932 57730 23108 57764
rect 23430 57730 23606 57764
rect 22720 57660 22760 57712
rect 22720 57560 22760 57600
rect 22720 57402 22746 57560
rect 22746 57402 22760 57560
rect 23790 57712 23802 57870
rect 23802 57712 23830 57870
rect 23790 57680 23830 57712
rect 23790 57560 23830 57600
rect 22932 57508 23108 57542
rect 23430 57508 23606 57542
rect 22848 57464 22882 57498
rect 23665 57464 23699 57498
rect 22932 57420 23108 57454
rect 23430 57420 23606 57454
rect 22720 57360 22760 57402
rect 23790 57402 23802 57560
rect 23802 57402 23830 57560
rect 23790 57360 23830 57402
rect 27710 57870 27750 57920
rect 27710 57712 27736 57870
rect 27736 57712 27750 57870
rect 28780 57870 28820 57920
rect 27922 57818 28098 57852
rect 28420 57818 28596 57852
rect 27838 57774 27872 57808
rect 28655 57774 28689 57808
rect 27922 57730 28098 57764
rect 28420 57730 28596 57764
rect 27710 57660 27750 57712
rect 27710 57560 27750 57600
rect 27710 57402 27736 57560
rect 27736 57402 27750 57560
rect 28780 57712 28792 57870
rect 28792 57712 28820 57870
rect 28780 57680 28820 57712
rect 28780 57560 28820 57600
rect 27922 57508 28098 57542
rect 28420 57508 28596 57542
rect 27838 57464 27872 57498
rect 28655 57464 28689 57498
rect 27922 57420 28098 57454
rect 28420 57420 28596 57454
rect 27710 57360 27750 57402
rect 28780 57402 28792 57560
rect 28792 57402 28820 57560
rect 28780 57360 28820 57402
rect 32700 57870 32740 57920
rect 32700 57712 32726 57870
rect 32726 57712 32740 57870
rect 33770 57870 33810 57920
rect 32912 57818 33088 57852
rect 33410 57818 33586 57852
rect 32828 57774 32862 57808
rect 33645 57774 33679 57808
rect 32912 57730 33088 57764
rect 33410 57730 33586 57764
rect 32700 57660 32740 57712
rect 32700 57560 32740 57600
rect 32700 57402 32726 57560
rect 32726 57402 32740 57560
rect 33770 57712 33782 57870
rect 33782 57712 33810 57870
rect 33770 57680 33810 57712
rect 33770 57560 33810 57600
rect 32912 57508 33088 57542
rect 33410 57508 33586 57542
rect 32828 57464 32862 57498
rect 33645 57464 33679 57498
rect 32912 57420 33088 57454
rect 33410 57420 33586 57454
rect 32700 57360 32740 57402
rect 33770 57402 33782 57560
rect 33782 57402 33810 57560
rect 33770 57360 33810 57402
rect 37690 57870 37730 57920
rect 37690 57712 37716 57870
rect 37716 57712 37730 57870
rect 38760 57870 38800 57920
rect 37902 57818 38078 57852
rect 38400 57818 38576 57852
rect 37818 57774 37852 57808
rect 38635 57774 38669 57808
rect 37902 57730 38078 57764
rect 38400 57730 38576 57764
rect 37690 57660 37730 57712
rect 37690 57560 37730 57600
rect 37690 57402 37716 57560
rect 37716 57402 37730 57560
rect 38760 57712 38772 57870
rect 38772 57712 38800 57870
rect 38760 57680 38800 57712
rect 38760 57560 38800 57600
rect 37902 57508 38078 57542
rect 38400 57508 38576 57542
rect 37818 57464 37852 57498
rect 38635 57464 38669 57498
rect 37902 57420 38078 57454
rect 38400 57420 38576 57454
rect 37690 57360 37730 57402
rect 38760 57402 38772 57560
rect 38772 57402 38800 57560
rect 38760 57360 38800 57402
rect 42680 57870 42720 57920
rect 42680 57712 42706 57870
rect 42706 57712 42720 57870
rect 43750 57870 43790 57920
rect 42892 57818 43068 57852
rect 43390 57818 43566 57852
rect 42808 57774 42842 57808
rect 43625 57774 43659 57808
rect 42892 57730 43068 57764
rect 43390 57730 43566 57764
rect 42680 57660 42720 57712
rect 42680 57560 42720 57600
rect 42680 57402 42706 57560
rect 42706 57402 42720 57560
rect 43750 57712 43762 57870
rect 43762 57712 43790 57870
rect 43750 57680 43790 57712
rect 43750 57560 43790 57600
rect 42892 57508 43068 57542
rect 43390 57508 43566 57542
rect 42808 57464 42842 57498
rect 43625 57464 43659 57498
rect 42892 57420 43068 57454
rect 43390 57420 43566 57454
rect 42680 57360 42720 57402
rect 43750 57402 43762 57560
rect 43762 57402 43790 57560
rect 43750 57360 43790 57402
rect 47670 57870 47710 57920
rect 47670 57712 47696 57870
rect 47696 57712 47710 57870
rect 48740 57870 48780 57920
rect 47882 57818 48058 57852
rect 48380 57818 48556 57852
rect 47798 57774 47832 57808
rect 48615 57774 48649 57808
rect 47882 57730 48058 57764
rect 48380 57730 48556 57764
rect 47670 57660 47710 57712
rect 47670 57560 47710 57600
rect 47670 57402 47696 57560
rect 47696 57402 47710 57560
rect 48740 57712 48752 57870
rect 48752 57712 48780 57870
rect 48740 57680 48780 57712
rect 48740 57560 48780 57600
rect 47882 57508 48058 57542
rect 48380 57508 48556 57542
rect 47798 57464 47832 57498
rect 48615 57464 48649 57498
rect 47882 57420 48058 57454
rect 48380 57420 48556 57454
rect 47670 57360 47710 57402
rect 48740 57402 48752 57560
rect 48752 57402 48780 57560
rect 48740 57360 48780 57402
rect 52660 57870 52700 57920
rect 52660 57712 52686 57870
rect 52686 57712 52700 57870
rect 53730 57870 53770 57920
rect 52872 57818 53048 57852
rect 53370 57818 53546 57852
rect 52788 57774 52822 57808
rect 53605 57774 53639 57808
rect 52872 57730 53048 57764
rect 53370 57730 53546 57764
rect 52660 57660 52700 57712
rect 52660 57560 52700 57600
rect 52660 57402 52686 57560
rect 52686 57402 52700 57560
rect 53730 57712 53742 57870
rect 53742 57712 53770 57870
rect 53730 57680 53770 57712
rect 53730 57560 53770 57600
rect 52872 57508 53048 57542
rect 53370 57508 53546 57542
rect 52788 57464 52822 57498
rect 53605 57464 53639 57498
rect 52872 57420 53048 57454
rect 53370 57420 53546 57454
rect 52660 57360 52700 57402
rect 53730 57402 53742 57560
rect 53742 57402 53770 57560
rect 53730 57360 53770 57402
rect 57650 57870 57690 57920
rect 57650 57712 57676 57870
rect 57676 57712 57690 57870
rect 58720 57870 58760 57920
rect 57862 57818 58038 57852
rect 58360 57818 58536 57852
rect 57778 57774 57812 57808
rect 58595 57774 58629 57808
rect 57862 57730 58038 57764
rect 58360 57730 58536 57764
rect 57650 57660 57690 57712
rect 57650 57560 57690 57600
rect 57650 57402 57676 57560
rect 57676 57402 57690 57560
rect 58720 57712 58732 57870
rect 58732 57712 58760 57870
rect 58720 57680 58760 57712
rect 58720 57560 58760 57600
rect 57862 57508 58038 57542
rect 58360 57508 58536 57542
rect 57778 57464 57812 57498
rect 58595 57464 58629 57498
rect 57862 57420 58038 57454
rect 58360 57420 58536 57454
rect 57650 57360 57690 57402
rect 58720 57402 58732 57560
rect 58732 57402 58760 57560
rect 58720 57360 58760 57402
rect 62640 57870 62680 57920
rect 62640 57712 62666 57870
rect 62666 57712 62680 57870
rect 63710 57870 63750 57920
rect 62852 57818 63028 57852
rect 63350 57818 63526 57852
rect 62768 57774 62802 57808
rect 63585 57774 63619 57808
rect 62852 57730 63028 57764
rect 63350 57730 63526 57764
rect 62640 57660 62680 57712
rect 62640 57560 62680 57600
rect 62640 57402 62666 57560
rect 62666 57402 62680 57560
rect 63710 57712 63722 57870
rect 63722 57712 63750 57870
rect 63710 57680 63750 57712
rect 63710 57560 63750 57600
rect 62852 57508 63028 57542
rect 63350 57508 63526 57542
rect 62768 57464 62802 57498
rect 63585 57464 63619 57498
rect 62852 57420 63028 57454
rect 63350 57420 63526 57454
rect 62640 57360 62680 57402
rect 63710 57402 63722 57560
rect 63722 57402 63750 57560
rect 63710 57360 63750 57402
rect 67630 57870 67670 57920
rect 67630 57712 67656 57870
rect 67656 57712 67670 57870
rect 68700 57870 68740 57920
rect 67842 57818 68018 57852
rect 68340 57818 68516 57852
rect 67758 57774 67792 57808
rect 68575 57774 68609 57808
rect 67842 57730 68018 57764
rect 68340 57730 68516 57764
rect 67630 57660 67670 57712
rect 67630 57560 67670 57600
rect 67630 57402 67656 57560
rect 67656 57402 67670 57560
rect 68700 57712 68712 57870
rect 68712 57712 68740 57870
rect 68700 57680 68740 57712
rect 68700 57560 68740 57600
rect 67842 57508 68018 57542
rect 68340 57508 68516 57542
rect 67758 57464 67792 57498
rect 68575 57464 68609 57498
rect 67842 57420 68018 57454
rect 68340 57420 68516 57454
rect 67630 57360 67670 57402
rect 68700 57402 68712 57560
rect 68712 57402 68740 57560
rect 68700 57360 68740 57402
rect 72620 57870 72660 57920
rect 72620 57712 72646 57870
rect 72646 57712 72660 57870
rect 73690 57870 73730 57920
rect 72832 57818 73008 57852
rect 73330 57818 73506 57852
rect 72748 57774 72782 57808
rect 73565 57774 73599 57808
rect 72832 57730 73008 57764
rect 73330 57730 73506 57764
rect 72620 57660 72660 57712
rect 72620 57560 72660 57600
rect 72620 57402 72646 57560
rect 72646 57402 72660 57560
rect 73690 57712 73702 57870
rect 73702 57712 73730 57870
rect 73690 57680 73730 57712
rect 73690 57560 73730 57600
rect 72832 57508 73008 57542
rect 73330 57508 73506 57542
rect 72748 57464 72782 57498
rect 73565 57464 73599 57498
rect 72832 57420 73008 57454
rect 73330 57420 73506 57454
rect 72620 57360 72660 57402
rect 73690 57402 73702 57560
rect 73702 57402 73730 57560
rect 73690 57360 73730 57402
rect 77610 57870 77650 57920
rect 77610 57712 77636 57870
rect 77636 57712 77650 57870
rect 78680 57870 78720 57920
rect 77822 57818 77998 57852
rect 78320 57818 78496 57852
rect 77738 57774 77772 57808
rect 78555 57774 78589 57808
rect 77822 57730 77998 57764
rect 78320 57730 78496 57764
rect 77610 57660 77650 57712
rect 77610 57560 77650 57600
rect 77610 57402 77636 57560
rect 77636 57402 77650 57560
rect 78680 57712 78692 57870
rect 78692 57712 78720 57870
rect 78680 57680 78720 57712
rect 78680 57560 78720 57600
rect 77822 57508 77998 57542
rect 78320 57508 78496 57542
rect 77738 57464 77772 57498
rect 78555 57464 78589 57498
rect 77822 57420 77998 57454
rect 78320 57420 78496 57454
rect 77610 57360 77650 57402
rect 78680 57402 78692 57560
rect 78692 57402 78720 57560
rect 78680 57360 78720 57402
rect 2760 56160 2800 56210
rect 2760 56002 2786 56160
rect 2786 56002 2800 56160
rect 3830 56160 3870 56210
rect 2972 56108 3148 56142
rect 3470 56108 3646 56142
rect 2888 56064 2922 56098
rect 3705 56064 3739 56098
rect 2972 56020 3148 56054
rect 3470 56020 3646 56054
rect 2760 55950 2800 56002
rect 2760 55850 2800 55890
rect 2760 55692 2786 55850
rect 2786 55692 2800 55850
rect 3830 56002 3842 56160
rect 3842 56002 3870 56160
rect 3830 55970 3870 56002
rect 3830 55850 3870 55890
rect 2972 55798 3148 55832
rect 3470 55798 3646 55832
rect 2888 55754 2922 55788
rect 3705 55754 3739 55788
rect 2972 55710 3148 55744
rect 3470 55710 3646 55744
rect 2760 55650 2800 55692
rect 3830 55692 3842 55850
rect 3842 55692 3870 55850
rect 3830 55650 3870 55692
rect 7750 56160 7790 56210
rect 7750 56002 7776 56160
rect 7776 56002 7790 56160
rect 8820 56160 8860 56210
rect 7962 56108 8138 56142
rect 8460 56108 8636 56142
rect 7878 56064 7912 56098
rect 8695 56064 8729 56098
rect 7962 56020 8138 56054
rect 8460 56020 8636 56054
rect 7750 55950 7790 56002
rect 7750 55850 7790 55890
rect 7750 55692 7776 55850
rect 7776 55692 7790 55850
rect 8820 56002 8832 56160
rect 8832 56002 8860 56160
rect 8820 55970 8860 56002
rect 8820 55850 8860 55890
rect 7962 55798 8138 55832
rect 8460 55798 8636 55832
rect 7878 55754 7912 55788
rect 8695 55754 8729 55788
rect 7962 55710 8138 55744
rect 8460 55710 8636 55744
rect 7750 55650 7790 55692
rect 8820 55692 8832 55850
rect 8832 55692 8860 55850
rect 8820 55650 8860 55692
rect 12740 56160 12780 56210
rect 12740 56002 12766 56160
rect 12766 56002 12780 56160
rect 13810 56160 13850 56210
rect 12952 56108 13128 56142
rect 13450 56108 13626 56142
rect 12868 56064 12902 56098
rect 13685 56064 13719 56098
rect 12952 56020 13128 56054
rect 13450 56020 13626 56054
rect 12740 55950 12780 56002
rect 12740 55850 12780 55890
rect 12740 55692 12766 55850
rect 12766 55692 12780 55850
rect 13810 56002 13822 56160
rect 13822 56002 13850 56160
rect 13810 55970 13850 56002
rect 13810 55850 13850 55890
rect 12952 55798 13128 55832
rect 13450 55798 13626 55832
rect 12868 55754 12902 55788
rect 13685 55754 13719 55788
rect 12952 55710 13128 55744
rect 13450 55710 13626 55744
rect 12740 55650 12780 55692
rect 13810 55692 13822 55850
rect 13822 55692 13850 55850
rect 13810 55650 13850 55692
rect 17730 56160 17770 56210
rect 17730 56002 17756 56160
rect 17756 56002 17770 56160
rect 18800 56160 18840 56210
rect 17942 56108 18118 56142
rect 18440 56108 18616 56142
rect 17858 56064 17892 56098
rect 18675 56064 18709 56098
rect 17942 56020 18118 56054
rect 18440 56020 18616 56054
rect 17730 55950 17770 56002
rect 17730 55850 17770 55890
rect 17730 55692 17756 55850
rect 17756 55692 17770 55850
rect 18800 56002 18812 56160
rect 18812 56002 18840 56160
rect 18800 55970 18840 56002
rect 18800 55850 18840 55890
rect 17942 55798 18118 55832
rect 18440 55798 18616 55832
rect 17858 55754 17892 55788
rect 18675 55754 18709 55788
rect 17942 55710 18118 55744
rect 18440 55710 18616 55744
rect 17730 55650 17770 55692
rect 18800 55692 18812 55850
rect 18812 55692 18840 55850
rect 18800 55650 18840 55692
rect 22720 56160 22760 56210
rect 22720 56002 22746 56160
rect 22746 56002 22760 56160
rect 23790 56160 23830 56210
rect 22932 56108 23108 56142
rect 23430 56108 23606 56142
rect 22848 56064 22882 56098
rect 23665 56064 23699 56098
rect 22932 56020 23108 56054
rect 23430 56020 23606 56054
rect 22720 55950 22760 56002
rect 22720 55850 22760 55890
rect 22720 55692 22746 55850
rect 22746 55692 22760 55850
rect 23790 56002 23802 56160
rect 23802 56002 23830 56160
rect 23790 55970 23830 56002
rect 23790 55850 23830 55890
rect 22932 55798 23108 55832
rect 23430 55798 23606 55832
rect 22848 55754 22882 55788
rect 23665 55754 23699 55788
rect 22932 55710 23108 55744
rect 23430 55710 23606 55744
rect 22720 55650 22760 55692
rect 23790 55692 23802 55850
rect 23802 55692 23830 55850
rect 23790 55650 23830 55692
rect 27710 56160 27750 56210
rect 27710 56002 27736 56160
rect 27736 56002 27750 56160
rect 28780 56160 28820 56210
rect 27922 56108 28098 56142
rect 28420 56108 28596 56142
rect 27838 56064 27872 56098
rect 28655 56064 28689 56098
rect 27922 56020 28098 56054
rect 28420 56020 28596 56054
rect 27710 55950 27750 56002
rect 27710 55850 27750 55890
rect 27710 55692 27736 55850
rect 27736 55692 27750 55850
rect 28780 56002 28792 56160
rect 28792 56002 28820 56160
rect 28780 55970 28820 56002
rect 28780 55850 28820 55890
rect 27922 55798 28098 55832
rect 28420 55798 28596 55832
rect 27838 55754 27872 55788
rect 28655 55754 28689 55788
rect 27922 55710 28098 55744
rect 28420 55710 28596 55744
rect 27710 55650 27750 55692
rect 28780 55692 28792 55850
rect 28792 55692 28820 55850
rect 28780 55650 28820 55692
rect 32700 56160 32740 56210
rect 32700 56002 32726 56160
rect 32726 56002 32740 56160
rect 33770 56160 33810 56210
rect 32912 56108 33088 56142
rect 33410 56108 33586 56142
rect 32828 56064 32862 56098
rect 33645 56064 33679 56098
rect 32912 56020 33088 56054
rect 33410 56020 33586 56054
rect 32700 55950 32740 56002
rect 32700 55850 32740 55890
rect 32700 55692 32726 55850
rect 32726 55692 32740 55850
rect 33770 56002 33782 56160
rect 33782 56002 33810 56160
rect 33770 55970 33810 56002
rect 33770 55850 33810 55890
rect 32912 55798 33088 55832
rect 33410 55798 33586 55832
rect 32828 55754 32862 55788
rect 33645 55754 33679 55788
rect 32912 55710 33088 55744
rect 33410 55710 33586 55744
rect 32700 55650 32740 55692
rect 33770 55692 33782 55850
rect 33782 55692 33810 55850
rect 33770 55650 33810 55692
rect 37690 56160 37730 56210
rect 37690 56002 37716 56160
rect 37716 56002 37730 56160
rect 38760 56160 38800 56210
rect 37902 56108 38078 56142
rect 38400 56108 38576 56142
rect 37818 56064 37852 56098
rect 38635 56064 38669 56098
rect 37902 56020 38078 56054
rect 38400 56020 38576 56054
rect 37690 55950 37730 56002
rect 37690 55850 37730 55890
rect 37690 55692 37716 55850
rect 37716 55692 37730 55850
rect 38760 56002 38772 56160
rect 38772 56002 38800 56160
rect 38760 55970 38800 56002
rect 38760 55850 38800 55890
rect 37902 55798 38078 55832
rect 38400 55798 38576 55832
rect 37818 55754 37852 55788
rect 38635 55754 38669 55788
rect 37902 55710 38078 55744
rect 38400 55710 38576 55744
rect 37690 55650 37730 55692
rect 38760 55692 38772 55850
rect 38772 55692 38800 55850
rect 38760 55650 38800 55692
rect 42680 56160 42720 56210
rect 42680 56002 42706 56160
rect 42706 56002 42720 56160
rect 43750 56160 43790 56210
rect 42892 56108 43068 56142
rect 43390 56108 43566 56142
rect 42808 56064 42842 56098
rect 43625 56064 43659 56098
rect 42892 56020 43068 56054
rect 43390 56020 43566 56054
rect 42680 55950 42720 56002
rect 42680 55850 42720 55890
rect 42680 55692 42706 55850
rect 42706 55692 42720 55850
rect 43750 56002 43762 56160
rect 43762 56002 43790 56160
rect 43750 55970 43790 56002
rect 43750 55850 43790 55890
rect 42892 55798 43068 55832
rect 43390 55798 43566 55832
rect 42808 55754 42842 55788
rect 43625 55754 43659 55788
rect 42892 55710 43068 55744
rect 43390 55710 43566 55744
rect 42680 55650 42720 55692
rect 43750 55692 43762 55850
rect 43762 55692 43790 55850
rect 43750 55650 43790 55692
rect 47670 56160 47710 56210
rect 47670 56002 47696 56160
rect 47696 56002 47710 56160
rect 48740 56160 48780 56210
rect 47882 56108 48058 56142
rect 48380 56108 48556 56142
rect 47798 56064 47832 56098
rect 48615 56064 48649 56098
rect 47882 56020 48058 56054
rect 48380 56020 48556 56054
rect 47670 55950 47710 56002
rect 47670 55850 47710 55890
rect 47670 55692 47696 55850
rect 47696 55692 47710 55850
rect 48740 56002 48752 56160
rect 48752 56002 48780 56160
rect 48740 55970 48780 56002
rect 48740 55850 48780 55890
rect 47882 55798 48058 55832
rect 48380 55798 48556 55832
rect 47798 55754 47832 55788
rect 48615 55754 48649 55788
rect 47882 55710 48058 55744
rect 48380 55710 48556 55744
rect 47670 55650 47710 55692
rect 48740 55692 48752 55850
rect 48752 55692 48780 55850
rect 48740 55650 48780 55692
rect 52660 56160 52700 56210
rect 52660 56002 52686 56160
rect 52686 56002 52700 56160
rect 53730 56160 53770 56210
rect 52872 56108 53048 56142
rect 53370 56108 53546 56142
rect 52788 56064 52822 56098
rect 53605 56064 53639 56098
rect 52872 56020 53048 56054
rect 53370 56020 53546 56054
rect 52660 55950 52700 56002
rect 52660 55850 52700 55890
rect 52660 55692 52686 55850
rect 52686 55692 52700 55850
rect 53730 56002 53742 56160
rect 53742 56002 53770 56160
rect 53730 55970 53770 56002
rect 53730 55850 53770 55890
rect 52872 55798 53048 55832
rect 53370 55798 53546 55832
rect 52788 55754 52822 55788
rect 53605 55754 53639 55788
rect 52872 55710 53048 55744
rect 53370 55710 53546 55744
rect 52660 55650 52700 55692
rect 53730 55692 53742 55850
rect 53742 55692 53770 55850
rect 53730 55650 53770 55692
rect 57650 56160 57690 56210
rect 57650 56002 57676 56160
rect 57676 56002 57690 56160
rect 58720 56160 58760 56210
rect 57862 56108 58038 56142
rect 58360 56108 58536 56142
rect 57778 56064 57812 56098
rect 58595 56064 58629 56098
rect 57862 56020 58038 56054
rect 58360 56020 58536 56054
rect 57650 55950 57690 56002
rect 57650 55850 57690 55890
rect 57650 55692 57676 55850
rect 57676 55692 57690 55850
rect 58720 56002 58732 56160
rect 58732 56002 58760 56160
rect 58720 55970 58760 56002
rect 58720 55850 58760 55890
rect 57862 55798 58038 55832
rect 58360 55798 58536 55832
rect 57778 55754 57812 55788
rect 58595 55754 58629 55788
rect 57862 55710 58038 55744
rect 58360 55710 58536 55744
rect 57650 55650 57690 55692
rect 58720 55692 58732 55850
rect 58732 55692 58760 55850
rect 58720 55650 58760 55692
rect 62640 56160 62680 56210
rect 62640 56002 62666 56160
rect 62666 56002 62680 56160
rect 63710 56160 63750 56210
rect 62852 56108 63028 56142
rect 63350 56108 63526 56142
rect 62768 56064 62802 56098
rect 63585 56064 63619 56098
rect 62852 56020 63028 56054
rect 63350 56020 63526 56054
rect 62640 55950 62680 56002
rect 62640 55850 62680 55890
rect 62640 55692 62666 55850
rect 62666 55692 62680 55850
rect 63710 56002 63722 56160
rect 63722 56002 63750 56160
rect 63710 55970 63750 56002
rect 63710 55850 63750 55890
rect 62852 55798 63028 55832
rect 63350 55798 63526 55832
rect 62768 55754 62802 55788
rect 63585 55754 63619 55788
rect 62852 55710 63028 55744
rect 63350 55710 63526 55744
rect 62640 55650 62680 55692
rect 63710 55692 63722 55850
rect 63722 55692 63750 55850
rect 63710 55650 63750 55692
rect 67630 56160 67670 56210
rect 67630 56002 67656 56160
rect 67656 56002 67670 56160
rect 68700 56160 68740 56210
rect 67842 56108 68018 56142
rect 68340 56108 68516 56142
rect 67758 56064 67792 56098
rect 68575 56064 68609 56098
rect 67842 56020 68018 56054
rect 68340 56020 68516 56054
rect 67630 55950 67670 56002
rect 67630 55850 67670 55890
rect 67630 55692 67656 55850
rect 67656 55692 67670 55850
rect 68700 56002 68712 56160
rect 68712 56002 68740 56160
rect 68700 55970 68740 56002
rect 68700 55850 68740 55890
rect 67842 55798 68018 55832
rect 68340 55798 68516 55832
rect 67758 55754 67792 55788
rect 68575 55754 68609 55788
rect 67842 55710 68018 55744
rect 68340 55710 68516 55744
rect 67630 55650 67670 55692
rect 68700 55692 68712 55850
rect 68712 55692 68740 55850
rect 68700 55650 68740 55692
rect 72620 56160 72660 56210
rect 72620 56002 72646 56160
rect 72646 56002 72660 56160
rect 73690 56160 73730 56210
rect 72832 56108 73008 56142
rect 73330 56108 73506 56142
rect 72748 56064 72782 56098
rect 73565 56064 73599 56098
rect 72832 56020 73008 56054
rect 73330 56020 73506 56054
rect 72620 55950 72660 56002
rect 72620 55850 72660 55890
rect 72620 55692 72646 55850
rect 72646 55692 72660 55850
rect 73690 56002 73702 56160
rect 73702 56002 73730 56160
rect 73690 55970 73730 56002
rect 73690 55850 73730 55890
rect 72832 55798 73008 55832
rect 73330 55798 73506 55832
rect 72748 55754 72782 55788
rect 73565 55754 73599 55788
rect 72832 55710 73008 55744
rect 73330 55710 73506 55744
rect 72620 55650 72660 55692
rect 73690 55692 73702 55850
rect 73702 55692 73730 55850
rect 73690 55650 73730 55692
rect 77610 56160 77650 56210
rect 77610 56002 77636 56160
rect 77636 56002 77650 56160
rect 78680 56160 78720 56210
rect 77822 56108 77998 56142
rect 78320 56108 78496 56142
rect 77738 56064 77772 56098
rect 78555 56064 78589 56098
rect 77822 56020 77998 56054
rect 78320 56020 78496 56054
rect 77610 55950 77650 56002
rect 77610 55850 77650 55890
rect 77610 55692 77636 55850
rect 77636 55692 77650 55850
rect 78680 56002 78692 56160
rect 78692 56002 78720 56160
rect 78680 55970 78720 56002
rect 78680 55850 78720 55890
rect 77822 55798 77998 55832
rect 78320 55798 78496 55832
rect 77738 55754 77772 55788
rect 78555 55754 78589 55788
rect 77822 55710 77998 55744
rect 78320 55710 78496 55744
rect 77610 55650 77650 55692
rect 78680 55692 78692 55850
rect 78692 55692 78720 55850
rect 78680 55650 78720 55692
rect 2760 54450 2800 54500
rect 2760 54292 2786 54450
rect 2786 54292 2800 54450
rect 3830 54450 3870 54500
rect 2972 54398 3148 54432
rect 3470 54398 3646 54432
rect 2888 54354 2922 54388
rect 3705 54354 3739 54388
rect 2972 54310 3148 54344
rect 3470 54310 3646 54344
rect 2760 54240 2800 54292
rect 2760 54140 2800 54180
rect 2760 53982 2786 54140
rect 2786 53982 2800 54140
rect 3830 54292 3842 54450
rect 3842 54292 3870 54450
rect 3830 54260 3870 54292
rect 3830 54140 3870 54180
rect 2972 54088 3148 54122
rect 3470 54088 3646 54122
rect 2888 54044 2922 54078
rect 3705 54044 3739 54078
rect 2972 54000 3148 54034
rect 3470 54000 3646 54034
rect 2760 53940 2800 53982
rect 3830 53982 3842 54140
rect 3842 53982 3870 54140
rect 3830 53940 3870 53982
rect 7750 54450 7790 54500
rect 7750 54292 7776 54450
rect 7776 54292 7790 54450
rect 8820 54450 8860 54500
rect 7962 54398 8138 54432
rect 8460 54398 8636 54432
rect 7878 54354 7912 54388
rect 8695 54354 8729 54388
rect 7962 54310 8138 54344
rect 8460 54310 8636 54344
rect 7750 54240 7790 54292
rect 7750 54140 7790 54180
rect 7750 53982 7776 54140
rect 7776 53982 7790 54140
rect 8820 54292 8832 54450
rect 8832 54292 8860 54450
rect 8820 54260 8860 54292
rect 8820 54140 8860 54180
rect 7962 54088 8138 54122
rect 8460 54088 8636 54122
rect 7878 54044 7912 54078
rect 8695 54044 8729 54078
rect 7962 54000 8138 54034
rect 8460 54000 8636 54034
rect 7750 53940 7790 53982
rect 8820 53982 8832 54140
rect 8832 53982 8860 54140
rect 8820 53940 8860 53982
rect 12740 54450 12780 54500
rect 12740 54292 12766 54450
rect 12766 54292 12780 54450
rect 13810 54450 13850 54500
rect 12952 54398 13128 54432
rect 13450 54398 13626 54432
rect 12868 54354 12902 54388
rect 13685 54354 13719 54388
rect 12952 54310 13128 54344
rect 13450 54310 13626 54344
rect 12740 54240 12780 54292
rect 12740 54140 12780 54180
rect 12740 53982 12766 54140
rect 12766 53982 12780 54140
rect 13810 54292 13822 54450
rect 13822 54292 13850 54450
rect 13810 54260 13850 54292
rect 13810 54140 13850 54180
rect 12952 54088 13128 54122
rect 13450 54088 13626 54122
rect 12868 54044 12902 54078
rect 13685 54044 13719 54078
rect 12952 54000 13128 54034
rect 13450 54000 13626 54034
rect 12740 53940 12780 53982
rect 13810 53982 13822 54140
rect 13822 53982 13850 54140
rect 13810 53940 13850 53982
rect 17730 54450 17770 54500
rect 17730 54292 17756 54450
rect 17756 54292 17770 54450
rect 18800 54450 18840 54500
rect 17942 54398 18118 54432
rect 18440 54398 18616 54432
rect 17858 54354 17892 54388
rect 18675 54354 18709 54388
rect 17942 54310 18118 54344
rect 18440 54310 18616 54344
rect 17730 54240 17770 54292
rect 17730 54140 17770 54180
rect 17730 53982 17756 54140
rect 17756 53982 17770 54140
rect 18800 54292 18812 54450
rect 18812 54292 18840 54450
rect 18800 54260 18840 54292
rect 18800 54140 18840 54180
rect 17942 54088 18118 54122
rect 18440 54088 18616 54122
rect 17858 54044 17892 54078
rect 18675 54044 18709 54078
rect 17942 54000 18118 54034
rect 18440 54000 18616 54034
rect 17730 53940 17770 53982
rect 18800 53982 18812 54140
rect 18812 53982 18840 54140
rect 18800 53940 18840 53982
rect 22720 54450 22760 54500
rect 22720 54292 22746 54450
rect 22746 54292 22760 54450
rect 23790 54450 23830 54500
rect 22932 54398 23108 54432
rect 23430 54398 23606 54432
rect 22848 54354 22882 54388
rect 23665 54354 23699 54388
rect 22932 54310 23108 54344
rect 23430 54310 23606 54344
rect 22720 54240 22760 54292
rect 22720 54140 22760 54180
rect 22720 53982 22746 54140
rect 22746 53982 22760 54140
rect 23790 54292 23802 54450
rect 23802 54292 23830 54450
rect 23790 54260 23830 54292
rect 23790 54140 23830 54180
rect 22932 54088 23108 54122
rect 23430 54088 23606 54122
rect 22848 54044 22882 54078
rect 23665 54044 23699 54078
rect 22932 54000 23108 54034
rect 23430 54000 23606 54034
rect 22720 53940 22760 53982
rect 23790 53982 23802 54140
rect 23802 53982 23830 54140
rect 23790 53940 23830 53982
rect 27710 54450 27750 54500
rect 27710 54292 27736 54450
rect 27736 54292 27750 54450
rect 28780 54450 28820 54500
rect 27922 54398 28098 54432
rect 28420 54398 28596 54432
rect 27838 54354 27872 54388
rect 28655 54354 28689 54388
rect 27922 54310 28098 54344
rect 28420 54310 28596 54344
rect 27710 54240 27750 54292
rect 27710 54140 27750 54180
rect 27710 53982 27736 54140
rect 27736 53982 27750 54140
rect 28780 54292 28792 54450
rect 28792 54292 28820 54450
rect 28780 54260 28820 54292
rect 28780 54140 28820 54180
rect 27922 54088 28098 54122
rect 28420 54088 28596 54122
rect 27838 54044 27872 54078
rect 28655 54044 28689 54078
rect 27922 54000 28098 54034
rect 28420 54000 28596 54034
rect 27710 53940 27750 53982
rect 28780 53982 28792 54140
rect 28792 53982 28820 54140
rect 28780 53940 28820 53982
rect 32700 54450 32740 54500
rect 32700 54292 32726 54450
rect 32726 54292 32740 54450
rect 33770 54450 33810 54500
rect 32912 54398 33088 54432
rect 33410 54398 33586 54432
rect 32828 54354 32862 54388
rect 33645 54354 33679 54388
rect 32912 54310 33088 54344
rect 33410 54310 33586 54344
rect 32700 54240 32740 54292
rect 32700 54140 32740 54180
rect 32700 53982 32726 54140
rect 32726 53982 32740 54140
rect 33770 54292 33782 54450
rect 33782 54292 33810 54450
rect 33770 54260 33810 54292
rect 33770 54140 33810 54180
rect 32912 54088 33088 54122
rect 33410 54088 33586 54122
rect 32828 54044 32862 54078
rect 33645 54044 33679 54078
rect 32912 54000 33088 54034
rect 33410 54000 33586 54034
rect 32700 53940 32740 53982
rect 33770 53982 33782 54140
rect 33782 53982 33810 54140
rect 33770 53940 33810 53982
rect 37690 54450 37730 54500
rect 37690 54292 37716 54450
rect 37716 54292 37730 54450
rect 38760 54450 38800 54500
rect 37902 54398 38078 54432
rect 38400 54398 38576 54432
rect 37818 54354 37852 54388
rect 38635 54354 38669 54388
rect 37902 54310 38078 54344
rect 38400 54310 38576 54344
rect 37690 54240 37730 54292
rect 37690 54140 37730 54180
rect 37690 53982 37716 54140
rect 37716 53982 37730 54140
rect 38760 54292 38772 54450
rect 38772 54292 38800 54450
rect 38760 54260 38800 54292
rect 38760 54140 38800 54180
rect 37902 54088 38078 54122
rect 38400 54088 38576 54122
rect 37818 54044 37852 54078
rect 38635 54044 38669 54078
rect 37902 54000 38078 54034
rect 38400 54000 38576 54034
rect 37690 53940 37730 53982
rect 38760 53982 38772 54140
rect 38772 53982 38800 54140
rect 38760 53940 38800 53982
rect 42680 54450 42720 54500
rect 42680 54292 42706 54450
rect 42706 54292 42720 54450
rect 43750 54450 43790 54500
rect 42892 54398 43068 54432
rect 43390 54398 43566 54432
rect 42808 54354 42842 54388
rect 43625 54354 43659 54388
rect 42892 54310 43068 54344
rect 43390 54310 43566 54344
rect 42680 54240 42720 54292
rect 42680 54140 42720 54180
rect 42680 53982 42706 54140
rect 42706 53982 42720 54140
rect 43750 54292 43762 54450
rect 43762 54292 43790 54450
rect 43750 54260 43790 54292
rect 43750 54140 43790 54180
rect 42892 54088 43068 54122
rect 43390 54088 43566 54122
rect 42808 54044 42842 54078
rect 43625 54044 43659 54078
rect 42892 54000 43068 54034
rect 43390 54000 43566 54034
rect 42680 53940 42720 53982
rect 43750 53982 43762 54140
rect 43762 53982 43790 54140
rect 43750 53940 43790 53982
rect 47670 54450 47710 54500
rect 47670 54292 47696 54450
rect 47696 54292 47710 54450
rect 48740 54450 48780 54500
rect 47882 54398 48058 54432
rect 48380 54398 48556 54432
rect 47798 54354 47832 54388
rect 48615 54354 48649 54388
rect 47882 54310 48058 54344
rect 48380 54310 48556 54344
rect 47670 54240 47710 54292
rect 47670 54140 47710 54180
rect 47670 53982 47696 54140
rect 47696 53982 47710 54140
rect 48740 54292 48752 54450
rect 48752 54292 48780 54450
rect 48740 54260 48780 54292
rect 48740 54140 48780 54180
rect 47882 54088 48058 54122
rect 48380 54088 48556 54122
rect 47798 54044 47832 54078
rect 48615 54044 48649 54078
rect 47882 54000 48058 54034
rect 48380 54000 48556 54034
rect 47670 53940 47710 53982
rect 48740 53982 48752 54140
rect 48752 53982 48780 54140
rect 48740 53940 48780 53982
rect 52660 54450 52700 54500
rect 52660 54292 52686 54450
rect 52686 54292 52700 54450
rect 53730 54450 53770 54500
rect 52872 54398 53048 54432
rect 53370 54398 53546 54432
rect 52788 54354 52822 54388
rect 53605 54354 53639 54388
rect 52872 54310 53048 54344
rect 53370 54310 53546 54344
rect 52660 54240 52700 54292
rect 52660 54140 52700 54180
rect 52660 53982 52686 54140
rect 52686 53982 52700 54140
rect 53730 54292 53742 54450
rect 53742 54292 53770 54450
rect 53730 54260 53770 54292
rect 53730 54140 53770 54180
rect 52872 54088 53048 54122
rect 53370 54088 53546 54122
rect 52788 54044 52822 54078
rect 53605 54044 53639 54078
rect 52872 54000 53048 54034
rect 53370 54000 53546 54034
rect 52660 53940 52700 53982
rect 53730 53982 53742 54140
rect 53742 53982 53770 54140
rect 53730 53940 53770 53982
rect 57650 54450 57690 54500
rect 57650 54292 57676 54450
rect 57676 54292 57690 54450
rect 58720 54450 58760 54500
rect 57862 54398 58038 54432
rect 58360 54398 58536 54432
rect 57778 54354 57812 54388
rect 58595 54354 58629 54388
rect 57862 54310 58038 54344
rect 58360 54310 58536 54344
rect 57650 54240 57690 54292
rect 57650 54140 57690 54180
rect 57650 53982 57676 54140
rect 57676 53982 57690 54140
rect 58720 54292 58732 54450
rect 58732 54292 58760 54450
rect 58720 54260 58760 54292
rect 58720 54140 58760 54180
rect 57862 54088 58038 54122
rect 58360 54088 58536 54122
rect 57778 54044 57812 54078
rect 58595 54044 58629 54078
rect 57862 54000 58038 54034
rect 58360 54000 58536 54034
rect 57650 53940 57690 53982
rect 58720 53982 58732 54140
rect 58732 53982 58760 54140
rect 58720 53940 58760 53982
rect 62640 54450 62680 54500
rect 62640 54292 62666 54450
rect 62666 54292 62680 54450
rect 63710 54450 63750 54500
rect 62852 54398 63028 54432
rect 63350 54398 63526 54432
rect 62768 54354 62802 54388
rect 63585 54354 63619 54388
rect 62852 54310 63028 54344
rect 63350 54310 63526 54344
rect 62640 54240 62680 54292
rect 62640 54140 62680 54180
rect 62640 53982 62666 54140
rect 62666 53982 62680 54140
rect 63710 54292 63722 54450
rect 63722 54292 63750 54450
rect 63710 54260 63750 54292
rect 63710 54140 63750 54180
rect 62852 54088 63028 54122
rect 63350 54088 63526 54122
rect 62768 54044 62802 54078
rect 63585 54044 63619 54078
rect 62852 54000 63028 54034
rect 63350 54000 63526 54034
rect 62640 53940 62680 53982
rect 63710 53982 63722 54140
rect 63722 53982 63750 54140
rect 63710 53940 63750 53982
rect 67630 54450 67670 54500
rect 67630 54292 67656 54450
rect 67656 54292 67670 54450
rect 68700 54450 68740 54500
rect 67842 54398 68018 54432
rect 68340 54398 68516 54432
rect 67758 54354 67792 54388
rect 68575 54354 68609 54388
rect 67842 54310 68018 54344
rect 68340 54310 68516 54344
rect 67630 54240 67670 54292
rect 67630 54140 67670 54180
rect 67630 53982 67656 54140
rect 67656 53982 67670 54140
rect 68700 54292 68712 54450
rect 68712 54292 68740 54450
rect 68700 54260 68740 54292
rect 68700 54140 68740 54180
rect 67842 54088 68018 54122
rect 68340 54088 68516 54122
rect 67758 54044 67792 54078
rect 68575 54044 68609 54078
rect 67842 54000 68018 54034
rect 68340 54000 68516 54034
rect 67630 53940 67670 53982
rect 68700 53982 68712 54140
rect 68712 53982 68740 54140
rect 68700 53940 68740 53982
rect 72620 54450 72660 54500
rect 72620 54292 72646 54450
rect 72646 54292 72660 54450
rect 73690 54450 73730 54500
rect 72832 54398 73008 54432
rect 73330 54398 73506 54432
rect 72748 54354 72782 54388
rect 73565 54354 73599 54388
rect 72832 54310 73008 54344
rect 73330 54310 73506 54344
rect 72620 54240 72660 54292
rect 72620 54140 72660 54180
rect 72620 53982 72646 54140
rect 72646 53982 72660 54140
rect 73690 54292 73702 54450
rect 73702 54292 73730 54450
rect 73690 54260 73730 54292
rect 73690 54140 73730 54180
rect 72832 54088 73008 54122
rect 73330 54088 73506 54122
rect 72748 54044 72782 54078
rect 73565 54044 73599 54078
rect 72832 54000 73008 54034
rect 73330 54000 73506 54034
rect 72620 53940 72660 53982
rect 73690 53982 73702 54140
rect 73702 53982 73730 54140
rect 73690 53940 73730 53982
rect 77610 54450 77650 54500
rect 77610 54292 77636 54450
rect 77636 54292 77650 54450
rect 78680 54450 78720 54500
rect 77822 54398 77998 54432
rect 78320 54398 78496 54432
rect 77738 54354 77772 54388
rect 78555 54354 78589 54388
rect 77822 54310 77998 54344
rect 78320 54310 78496 54344
rect 77610 54240 77650 54292
rect 77610 54140 77650 54180
rect 77610 53982 77636 54140
rect 77636 53982 77650 54140
rect 78680 54292 78692 54450
rect 78692 54292 78720 54450
rect 78680 54260 78720 54292
rect 78680 54140 78720 54180
rect 77822 54088 77998 54122
rect 78320 54088 78496 54122
rect 77738 54044 77772 54078
rect 78555 54044 78589 54078
rect 77822 54000 77998 54034
rect 78320 54000 78496 54034
rect 77610 53940 77650 53982
rect 78680 53982 78692 54140
rect 78692 53982 78720 54140
rect 78680 53940 78720 53982
rect 2760 52740 2800 52790
rect 2760 52582 2786 52740
rect 2786 52582 2800 52740
rect 3830 52740 3870 52790
rect 2972 52688 3148 52722
rect 3470 52688 3646 52722
rect 2888 52644 2922 52678
rect 3705 52644 3739 52678
rect 2972 52600 3148 52634
rect 3470 52600 3646 52634
rect 2760 52530 2800 52582
rect 2760 52430 2800 52470
rect 2760 52272 2786 52430
rect 2786 52272 2800 52430
rect 3830 52582 3842 52740
rect 3842 52582 3870 52740
rect 3830 52550 3870 52582
rect 3830 52430 3870 52470
rect 2972 52378 3148 52412
rect 3470 52378 3646 52412
rect 2888 52334 2922 52368
rect 3705 52334 3739 52368
rect 2972 52290 3148 52324
rect 3470 52290 3646 52324
rect 2760 52230 2800 52272
rect 3830 52272 3842 52430
rect 3842 52272 3870 52430
rect 3830 52230 3870 52272
rect 7750 52740 7790 52790
rect 7750 52582 7776 52740
rect 7776 52582 7790 52740
rect 8820 52740 8860 52790
rect 7962 52688 8138 52722
rect 8460 52688 8636 52722
rect 7878 52644 7912 52678
rect 8695 52644 8729 52678
rect 7962 52600 8138 52634
rect 8460 52600 8636 52634
rect 7750 52530 7790 52582
rect 7750 52430 7790 52470
rect 7750 52272 7776 52430
rect 7776 52272 7790 52430
rect 8820 52582 8832 52740
rect 8832 52582 8860 52740
rect 8820 52550 8860 52582
rect 8820 52430 8860 52470
rect 7962 52378 8138 52412
rect 8460 52378 8636 52412
rect 7878 52334 7912 52368
rect 8695 52334 8729 52368
rect 7962 52290 8138 52324
rect 8460 52290 8636 52324
rect 7750 52230 7790 52272
rect 8820 52272 8832 52430
rect 8832 52272 8860 52430
rect 8820 52230 8860 52272
rect 12740 52740 12780 52790
rect 12740 52582 12766 52740
rect 12766 52582 12780 52740
rect 13810 52740 13850 52790
rect 12952 52688 13128 52722
rect 13450 52688 13626 52722
rect 12868 52644 12902 52678
rect 13685 52644 13719 52678
rect 12952 52600 13128 52634
rect 13450 52600 13626 52634
rect 12740 52530 12780 52582
rect 12740 52430 12780 52470
rect 12740 52272 12766 52430
rect 12766 52272 12780 52430
rect 13810 52582 13822 52740
rect 13822 52582 13850 52740
rect 13810 52550 13850 52582
rect 13810 52430 13850 52470
rect 12952 52378 13128 52412
rect 13450 52378 13626 52412
rect 12868 52334 12902 52368
rect 13685 52334 13719 52368
rect 12952 52290 13128 52324
rect 13450 52290 13626 52324
rect 12740 52230 12780 52272
rect 13810 52272 13822 52430
rect 13822 52272 13850 52430
rect 13810 52230 13850 52272
rect 17730 52740 17770 52790
rect 17730 52582 17756 52740
rect 17756 52582 17770 52740
rect 18800 52740 18840 52790
rect 17942 52688 18118 52722
rect 18440 52688 18616 52722
rect 17858 52644 17892 52678
rect 18675 52644 18709 52678
rect 17942 52600 18118 52634
rect 18440 52600 18616 52634
rect 17730 52530 17770 52582
rect 17730 52430 17770 52470
rect 17730 52272 17756 52430
rect 17756 52272 17770 52430
rect 18800 52582 18812 52740
rect 18812 52582 18840 52740
rect 18800 52550 18840 52582
rect 18800 52430 18840 52470
rect 17942 52378 18118 52412
rect 18440 52378 18616 52412
rect 17858 52334 17892 52368
rect 18675 52334 18709 52368
rect 17942 52290 18118 52324
rect 18440 52290 18616 52324
rect 17730 52230 17770 52272
rect 18800 52272 18812 52430
rect 18812 52272 18840 52430
rect 18800 52230 18840 52272
rect 22720 52740 22760 52790
rect 22720 52582 22746 52740
rect 22746 52582 22760 52740
rect 23790 52740 23830 52790
rect 22932 52688 23108 52722
rect 23430 52688 23606 52722
rect 22848 52644 22882 52678
rect 23665 52644 23699 52678
rect 22932 52600 23108 52634
rect 23430 52600 23606 52634
rect 22720 52530 22760 52582
rect 22720 52430 22760 52470
rect 22720 52272 22746 52430
rect 22746 52272 22760 52430
rect 23790 52582 23802 52740
rect 23802 52582 23830 52740
rect 23790 52550 23830 52582
rect 23790 52430 23830 52470
rect 22932 52378 23108 52412
rect 23430 52378 23606 52412
rect 22848 52334 22882 52368
rect 23665 52334 23699 52368
rect 22932 52290 23108 52324
rect 23430 52290 23606 52324
rect 22720 52230 22760 52272
rect 23790 52272 23802 52430
rect 23802 52272 23830 52430
rect 23790 52230 23830 52272
rect 27710 52740 27750 52790
rect 27710 52582 27736 52740
rect 27736 52582 27750 52740
rect 28780 52740 28820 52790
rect 27922 52688 28098 52722
rect 28420 52688 28596 52722
rect 27838 52644 27872 52678
rect 28655 52644 28689 52678
rect 27922 52600 28098 52634
rect 28420 52600 28596 52634
rect 27710 52530 27750 52582
rect 27710 52430 27750 52470
rect 27710 52272 27736 52430
rect 27736 52272 27750 52430
rect 28780 52582 28792 52740
rect 28792 52582 28820 52740
rect 28780 52550 28820 52582
rect 28780 52430 28820 52470
rect 27922 52378 28098 52412
rect 28420 52378 28596 52412
rect 27838 52334 27872 52368
rect 28655 52334 28689 52368
rect 27922 52290 28098 52324
rect 28420 52290 28596 52324
rect 27710 52230 27750 52272
rect 28780 52272 28792 52430
rect 28792 52272 28820 52430
rect 28780 52230 28820 52272
rect 32700 52740 32740 52790
rect 32700 52582 32726 52740
rect 32726 52582 32740 52740
rect 33770 52740 33810 52790
rect 32912 52688 33088 52722
rect 33410 52688 33586 52722
rect 32828 52644 32862 52678
rect 33645 52644 33679 52678
rect 32912 52600 33088 52634
rect 33410 52600 33586 52634
rect 32700 52530 32740 52582
rect 32700 52430 32740 52470
rect 32700 52272 32726 52430
rect 32726 52272 32740 52430
rect 33770 52582 33782 52740
rect 33782 52582 33810 52740
rect 33770 52550 33810 52582
rect 33770 52430 33810 52470
rect 32912 52378 33088 52412
rect 33410 52378 33586 52412
rect 32828 52334 32862 52368
rect 33645 52334 33679 52368
rect 32912 52290 33088 52324
rect 33410 52290 33586 52324
rect 32700 52230 32740 52272
rect 33770 52272 33782 52430
rect 33782 52272 33810 52430
rect 33770 52230 33810 52272
rect 37690 52740 37730 52790
rect 37690 52582 37716 52740
rect 37716 52582 37730 52740
rect 38760 52740 38800 52790
rect 37902 52688 38078 52722
rect 38400 52688 38576 52722
rect 37818 52644 37852 52678
rect 38635 52644 38669 52678
rect 37902 52600 38078 52634
rect 38400 52600 38576 52634
rect 37690 52530 37730 52582
rect 37690 52430 37730 52470
rect 37690 52272 37716 52430
rect 37716 52272 37730 52430
rect 38760 52582 38772 52740
rect 38772 52582 38800 52740
rect 38760 52550 38800 52582
rect 38760 52430 38800 52470
rect 37902 52378 38078 52412
rect 38400 52378 38576 52412
rect 37818 52334 37852 52368
rect 38635 52334 38669 52368
rect 37902 52290 38078 52324
rect 38400 52290 38576 52324
rect 37690 52230 37730 52272
rect 38760 52272 38772 52430
rect 38772 52272 38800 52430
rect 38760 52230 38800 52272
rect 42680 52740 42720 52790
rect 42680 52582 42706 52740
rect 42706 52582 42720 52740
rect 43750 52740 43790 52790
rect 42892 52688 43068 52722
rect 43390 52688 43566 52722
rect 42808 52644 42842 52678
rect 43625 52644 43659 52678
rect 42892 52600 43068 52634
rect 43390 52600 43566 52634
rect 42680 52530 42720 52582
rect 42680 52430 42720 52470
rect 42680 52272 42706 52430
rect 42706 52272 42720 52430
rect 43750 52582 43762 52740
rect 43762 52582 43790 52740
rect 43750 52550 43790 52582
rect 43750 52430 43790 52470
rect 42892 52378 43068 52412
rect 43390 52378 43566 52412
rect 42808 52334 42842 52368
rect 43625 52334 43659 52368
rect 42892 52290 43068 52324
rect 43390 52290 43566 52324
rect 42680 52230 42720 52272
rect 43750 52272 43762 52430
rect 43762 52272 43790 52430
rect 43750 52230 43790 52272
rect 47670 52740 47710 52790
rect 47670 52582 47696 52740
rect 47696 52582 47710 52740
rect 48740 52740 48780 52790
rect 47882 52688 48058 52722
rect 48380 52688 48556 52722
rect 47798 52644 47832 52678
rect 48615 52644 48649 52678
rect 47882 52600 48058 52634
rect 48380 52600 48556 52634
rect 47670 52530 47710 52582
rect 47670 52430 47710 52470
rect 47670 52272 47696 52430
rect 47696 52272 47710 52430
rect 48740 52582 48752 52740
rect 48752 52582 48780 52740
rect 48740 52550 48780 52582
rect 48740 52430 48780 52470
rect 47882 52378 48058 52412
rect 48380 52378 48556 52412
rect 47798 52334 47832 52368
rect 48615 52334 48649 52368
rect 47882 52290 48058 52324
rect 48380 52290 48556 52324
rect 47670 52230 47710 52272
rect 48740 52272 48752 52430
rect 48752 52272 48780 52430
rect 48740 52230 48780 52272
rect 52660 52740 52700 52790
rect 52660 52582 52686 52740
rect 52686 52582 52700 52740
rect 53730 52740 53770 52790
rect 52872 52688 53048 52722
rect 53370 52688 53546 52722
rect 52788 52644 52822 52678
rect 53605 52644 53639 52678
rect 52872 52600 53048 52634
rect 53370 52600 53546 52634
rect 52660 52530 52700 52582
rect 52660 52430 52700 52470
rect 52660 52272 52686 52430
rect 52686 52272 52700 52430
rect 53730 52582 53742 52740
rect 53742 52582 53770 52740
rect 53730 52550 53770 52582
rect 53730 52430 53770 52470
rect 52872 52378 53048 52412
rect 53370 52378 53546 52412
rect 52788 52334 52822 52368
rect 53605 52334 53639 52368
rect 52872 52290 53048 52324
rect 53370 52290 53546 52324
rect 52660 52230 52700 52272
rect 53730 52272 53742 52430
rect 53742 52272 53770 52430
rect 53730 52230 53770 52272
rect 57650 52740 57690 52790
rect 57650 52582 57676 52740
rect 57676 52582 57690 52740
rect 58720 52740 58760 52790
rect 57862 52688 58038 52722
rect 58360 52688 58536 52722
rect 57778 52644 57812 52678
rect 58595 52644 58629 52678
rect 57862 52600 58038 52634
rect 58360 52600 58536 52634
rect 57650 52530 57690 52582
rect 57650 52430 57690 52470
rect 57650 52272 57676 52430
rect 57676 52272 57690 52430
rect 58720 52582 58732 52740
rect 58732 52582 58760 52740
rect 58720 52550 58760 52582
rect 58720 52430 58760 52470
rect 57862 52378 58038 52412
rect 58360 52378 58536 52412
rect 57778 52334 57812 52368
rect 58595 52334 58629 52368
rect 57862 52290 58038 52324
rect 58360 52290 58536 52324
rect 57650 52230 57690 52272
rect 58720 52272 58732 52430
rect 58732 52272 58760 52430
rect 58720 52230 58760 52272
rect 62640 52740 62680 52790
rect 62640 52582 62666 52740
rect 62666 52582 62680 52740
rect 63710 52740 63750 52790
rect 62852 52688 63028 52722
rect 63350 52688 63526 52722
rect 62768 52644 62802 52678
rect 63585 52644 63619 52678
rect 62852 52600 63028 52634
rect 63350 52600 63526 52634
rect 62640 52530 62680 52582
rect 62640 52430 62680 52470
rect 62640 52272 62666 52430
rect 62666 52272 62680 52430
rect 63710 52582 63722 52740
rect 63722 52582 63750 52740
rect 63710 52550 63750 52582
rect 63710 52430 63750 52470
rect 62852 52378 63028 52412
rect 63350 52378 63526 52412
rect 62768 52334 62802 52368
rect 63585 52334 63619 52368
rect 62852 52290 63028 52324
rect 63350 52290 63526 52324
rect 62640 52230 62680 52272
rect 63710 52272 63722 52430
rect 63722 52272 63750 52430
rect 63710 52230 63750 52272
rect 67630 52740 67670 52790
rect 67630 52582 67656 52740
rect 67656 52582 67670 52740
rect 68700 52740 68740 52790
rect 67842 52688 68018 52722
rect 68340 52688 68516 52722
rect 67758 52644 67792 52678
rect 68575 52644 68609 52678
rect 67842 52600 68018 52634
rect 68340 52600 68516 52634
rect 67630 52530 67670 52582
rect 67630 52430 67670 52470
rect 67630 52272 67656 52430
rect 67656 52272 67670 52430
rect 68700 52582 68712 52740
rect 68712 52582 68740 52740
rect 68700 52550 68740 52582
rect 68700 52430 68740 52470
rect 67842 52378 68018 52412
rect 68340 52378 68516 52412
rect 67758 52334 67792 52368
rect 68575 52334 68609 52368
rect 67842 52290 68018 52324
rect 68340 52290 68516 52324
rect 67630 52230 67670 52272
rect 68700 52272 68712 52430
rect 68712 52272 68740 52430
rect 68700 52230 68740 52272
rect 72620 52740 72660 52790
rect 72620 52582 72646 52740
rect 72646 52582 72660 52740
rect 73690 52740 73730 52790
rect 72832 52688 73008 52722
rect 73330 52688 73506 52722
rect 72748 52644 72782 52678
rect 73565 52644 73599 52678
rect 72832 52600 73008 52634
rect 73330 52600 73506 52634
rect 72620 52530 72660 52582
rect 72620 52430 72660 52470
rect 72620 52272 72646 52430
rect 72646 52272 72660 52430
rect 73690 52582 73702 52740
rect 73702 52582 73730 52740
rect 73690 52550 73730 52582
rect 73690 52430 73730 52470
rect 72832 52378 73008 52412
rect 73330 52378 73506 52412
rect 72748 52334 72782 52368
rect 73565 52334 73599 52368
rect 72832 52290 73008 52324
rect 73330 52290 73506 52324
rect 72620 52230 72660 52272
rect 73690 52272 73702 52430
rect 73702 52272 73730 52430
rect 73690 52230 73730 52272
rect 77610 52740 77650 52790
rect 77610 52582 77636 52740
rect 77636 52582 77650 52740
rect 78680 52740 78720 52790
rect 77822 52688 77998 52722
rect 78320 52688 78496 52722
rect 77738 52644 77772 52678
rect 78555 52644 78589 52678
rect 77822 52600 77998 52634
rect 78320 52600 78496 52634
rect 77610 52530 77650 52582
rect 77610 52430 77650 52470
rect 77610 52272 77636 52430
rect 77636 52272 77650 52430
rect 78680 52582 78692 52740
rect 78692 52582 78720 52740
rect 78680 52550 78720 52582
rect 78680 52430 78720 52470
rect 77822 52378 77998 52412
rect 78320 52378 78496 52412
rect 77738 52334 77772 52368
rect 78555 52334 78589 52368
rect 77822 52290 77998 52324
rect 78320 52290 78496 52324
rect 77610 52230 77650 52272
rect 78680 52272 78692 52430
rect 78692 52272 78720 52430
rect 78680 52230 78720 52272
rect 2760 51030 2800 51080
rect 2760 50872 2786 51030
rect 2786 50872 2800 51030
rect 3830 51030 3870 51080
rect 2972 50978 3148 51012
rect 3470 50978 3646 51012
rect 2888 50934 2922 50968
rect 3705 50934 3739 50968
rect 2972 50890 3148 50924
rect 3470 50890 3646 50924
rect 2760 50820 2800 50872
rect 2760 50720 2800 50760
rect 2760 50562 2786 50720
rect 2786 50562 2800 50720
rect 3830 50872 3842 51030
rect 3842 50872 3870 51030
rect 3830 50840 3870 50872
rect 3830 50720 3870 50760
rect 2972 50668 3148 50702
rect 3470 50668 3646 50702
rect 2888 50624 2922 50658
rect 3705 50624 3739 50658
rect 2972 50580 3148 50614
rect 3470 50580 3646 50614
rect 2760 50520 2800 50562
rect 3830 50562 3842 50720
rect 3842 50562 3870 50720
rect 3830 50520 3870 50562
rect 7750 51030 7790 51080
rect 7750 50872 7776 51030
rect 7776 50872 7790 51030
rect 8820 51030 8860 51080
rect 7962 50978 8138 51012
rect 8460 50978 8636 51012
rect 7878 50934 7912 50968
rect 8695 50934 8729 50968
rect 7962 50890 8138 50924
rect 8460 50890 8636 50924
rect 7750 50820 7790 50872
rect 7750 50720 7790 50760
rect 7750 50562 7776 50720
rect 7776 50562 7790 50720
rect 8820 50872 8832 51030
rect 8832 50872 8860 51030
rect 8820 50840 8860 50872
rect 8820 50720 8860 50760
rect 7962 50668 8138 50702
rect 8460 50668 8636 50702
rect 7878 50624 7912 50658
rect 8695 50624 8729 50658
rect 7962 50580 8138 50614
rect 8460 50580 8636 50614
rect 7750 50520 7790 50562
rect 8820 50562 8832 50720
rect 8832 50562 8860 50720
rect 8820 50520 8860 50562
rect 12740 51030 12780 51080
rect 12740 50872 12766 51030
rect 12766 50872 12780 51030
rect 13810 51030 13850 51080
rect 12952 50978 13128 51012
rect 13450 50978 13626 51012
rect 12868 50934 12902 50968
rect 13685 50934 13719 50968
rect 12952 50890 13128 50924
rect 13450 50890 13626 50924
rect 12740 50820 12780 50872
rect 12740 50720 12780 50760
rect 12740 50562 12766 50720
rect 12766 50562 12780 50720
rect 13810 50872 13822 51030
rect 13822 50872 13850 51030
rect 13810 50840 13850 50872
rect 13810 50720 13850 50760
rect 12952 50668 13128 50702
rect 13450 50668 13626 50702
rect 12868 50624 12902 50658
rect 13685 50624 13719 50658
rect 12952 50580 13128 50614
rect 13450 50580 13626 50614
rect 12740 50520 12780 50562
rect 13810 50562 13822 50720
rect 13822 50562 13850 50720
rect 13810 50520 13850 50562
rect 17730 51030 17770 51080
rect 17730 50872 17756 51030
rect 17756 50872 17770 51030
rect 18800 51030 18840 51080
rect 17942 50978 18118 51012
rect 18440 50978 18616 51012
rect 17858 50934 17892 50968
rect 18675 50934 18709 50968
rect 17942 50890 18118 50924
rect 18440 50890 18616 50924
rect 17730 50820 17770 50872
rect 17730 50720 17770 50760
rect 17730 50562 17756 50720
rect 17756 50562 17770 50720
rect 18800 50872 18812 51030
rect 18812 50872 18840 51030
rect 18800 50840 18840 50872
rect 18800 50720 18840 50760
rect 17942 50668 18118 50702
rect 18440 50668 18616 50702
rect 17858 50624 17892 50658
rect 18675 50624 18709 50658
rect 17942 50580 18118 50614
rect 18440 50580 18616 50614
rect 17730 50520 17770 50562
rect 18800 50562 18812 50720
rect 18812 50562 18840 50720
rect 18800 50520 18840 50562
rect 22720 51030 22760 51080
rect 22720 50872 22746 51030
rect 22746 50872 22760 51030
rect 23790 51030 23830 51080
rect 22932 50978 23108 51012
rect 23430 50978 23606 51012
rect 22848 50934 22882 50968
rect 23665 50934 23699 50968
rect 22932 50890 23108 50924
rect 23430 50890 23606 50924
rect 22720 50820 22760 50872
rect 22720 50720 22760 50760
rect 22720 50562 22746 50720
rect 22746 50562 22760 50720
rect 23790 50872 23802 51030
rect 23802 50872 23830 51030
rect 23790 50840 23830 50872
rect 23790 50720 23830 50760
rect 22932 50668 23108 50702
rect 23430 50668 23606 50702
rect 22848 50624 22882 50658
rect 23665 50624 23699 50658
rect 22932 50580 23108 50614
rect 23430 50580 23606 50614
rect 22720 50520 22760 50562
rect 23790 50562 23802 50720
rect 23802 50562 23830 50720
rect 23790 50520 23830 50562
rect 27710 51030 27750 51080
rect 27710 50872 27736 51030
rect 27736 50872 27750 51030
rect 28780 51030 28820 51080
rect 27922 50978 28098 51012
rect 28420 50978 28596 51012
rect 27838 50934 27872 50968
rect 28655 50934 28689 50968
rect 27922 50890 28098 50924
rect 28420 50890 28596 50924
rect 27710 50820 27750 50872
rect 27710 50720 27750 50760
rect 27710 50562 27736 50720
rect 27736 50562 27750 50720
rect 28780 50872 28792 51030
rect 28792 50872 28820 51030
rect 28780 50840 28820 50872
rect 28780 50720 28820 50760
rect 27922 50668 28098 50702
rect 28420 50668 28596 50702
rect 27838 50624 27872 50658
rect 28655 50624 28689 50658
rect 27922 50580 28098 50614
rect 28420 50580 28596 50614
rect 27710 50520 27750 50562
rect 28780 50562 28792 50720
rect 28792 50562 28820 50720
rect 28780 50520 28820 50562
rect 32700 51030 32740 51080
rect 32700 50872 32726 51030
rect 32726 50872 32740 51030
rect 33770 51030 33810 51080
rect 32912 50978 33088 51012
rect 33410 50978 33586 51012
rect 32828 50934 32862 50968
rect 33645 50934 33679 50968
rect 32912 50890 33088 50924
rect 33410 50890 33586 50924
rect 32700 50820 32740 50872
rect 32700 50720 32740 50760
rect 32700 50562 32726 50720
rect 32726 50562 32740 50720
rect 33770 50872 33782 51030
rect 33782 50872 33810 51030
rect 33770 50840 33810 50872
rect 33770 50720 33810 50760
rect 32912 50668 33088 50702
rect 33410 50668 33586 50702
rect 32828 50624 32862 50658
rect 33645 50624 33679 50658
rect 32912 50580 33088 50614
rect 33410 50580 33586 50614
rect 32700 50520 32740 50562
rect 33770 50562 33782 50720
rect 33782 50562 33810 50720
rect 33770 50520 33810 50562
rect 37690 51030 37730 51080
rect 37690 50872 37716 51030
rect 37716 50872 37730 51030
rect 38760 51030 38800 51080
rect 37902 50978 38078 51012
rect 38400 50978 38576 51012
rect 37818 50934 37852 50968
rect 38635 50934 38669 50968
rect 37902 50890 38078 50924
rect 38400 50890 38576 50924
rect 37690 50820 37730 50872
rect 37690 50720 37730 50760
rect 37690 50562 37716 50720
rect 37716 50562 37730 50720
rect 38760 50872 38772 51030
rect 38772 50872 38800 51030
rect 38760 50840 38800 50872
rect 38760 50720 38800 50760
rect 37902 50668 38078 50702
rect 38400 50668 38576 50702
rect 37818 50624 37852 50658
rect 38635 50624 38669 50658
rect 37902 50580 38078 50614
rect 38400 50580 38576 50614
rect 37690 50520 37730 50562
rect 38760 50562 38772 50720
rect 38772 50562 38800 50720
rect 38760 50520 38800 50562
rect 42680 51030 42720 51080
rect 42680 50872 42706 51030
rect 42706 50872 42720 51030
rect 43750 51030 43790 51080
rect 42892 50978 43068 51012
rect 43390 50978 43566 51012
rect 42808 50934 42842 50968
rect 43625 50934 43659 50968
rect 42892 50890 43068 50924
rect 43390 50890 43566 50924
rect 42680 50820 42720 50872
rect 42680 50720 42720 50760
rect 42680 50562 42706 50720
rect 42706 50562 42720 50720
rect 43750 50872 43762 51030
rect 43762 50872 43790 51030
rect 43750 50840 43790 50872
rect 43750 50720 43790 50760
rect 42892 50668 43068 50702
rect 43390 50668 43566 50702
rect 42808 50624 42842 50658
rect 43625 50624 43659 50658
rect 42892 50580 43068 50614
rect 43390 50580 43566 50614
rect 42680 50520 42720 50562
rect 43750 50562 43762 50720
rect 43762 50562 43790 50720
rect 43750 50520 43790 50562
rect 47670 51030 47710 51080
rect 47670 50872 47696 51030
rect 47696 50872 47710 51030
rect 48740 51030 48780 51080
rect 47882 50978 48058 51012
rect 48380 50978 48556 51012
rect 47798 50934 47832 50968
rect 48615 50934 48649 50968
rect 47882 50890 48058 50924
rect 48380 50890 48556 50924
rect 47670 50820 47710 50872
rect 47670 50720 47710 50760
rect 47670 50562 47696 50720
rect 47696 50562 47710 50720
rect 48740 50872 48752 51030
rect 48752 50872 48780 51030
rect 48740 50840 48780 50872
rect 48740 50720 48780 50760
rect 47882 50668 48058 50702
rect 48380 50668 48556 50702
rect 47798 50624 47832 50658
rect 48615 50624 48649 50658
rect 47882 50580 48058 50614
rect 48380 50580 48556 50614
rect 47670 50520 47710 50562
rect 48740 50562 48752 50720
rect 48752 50562 48780 50720
rect 48740 50520 48780 50562
rect 52660 51030 52700 51080
rect 52660 50872 52686 51030
rect 52686 50872 52700 51030
rect 53730 51030 53770 51080
rect 52872 50978 53048 51012
rect 53370 50978 53546 51012
rect 52788 50934 52822 50968
rect 53605 50934 53639 50968
rect 52872 50890 53048 50924
rect 53370 50890 53546 50924
rect 52660 50820 52700 50872
rect 52660 50720 52700 50760
rect 52660 50562 52686 50720
rect 52686 50562 52700 50720
rect 53730 50872 53742 51030
rect 53742 50872 53770 51030
rect 53730 50840 53770 50872
rect 53730 50720 53770 50760
rect 52872 50668 53048 50702
rect 53370 50668 53546 50702
rect 52788 50624 52822 50658
rect 53605 50624 53639 50658
rect 52872 50580 53048 50614
rect 53370 50580 53546 50614
rect 52660 50520 52700 50562
rect 53730 50562 53742 50720
rect 53742 50562 53770 50720
rect 53730 50520 53770 50562
rect 57650 51030 57690 51080
rect 57650 50872 57676 51030
rect 57676 50872 57690 51030
rect 58720 51030 58760 51080
rect 57862 50978 58038 51012
rect 58360 50978 58536 51012
rect 57778 50934 57812 50968
rect 58595 50934 58629 50968
rect 57862 50890 58038 50924
rect 58360 50890 58536 50924
rect 57650 50820 57690 50872
rect 57650 50720 57690 50760
rect 57650 50562 57676 50720
rect 57676 50562 57690 50720
rect 58720 50872 58732 51030
rect 58732 50872 58760 51030
rect 58720 50840 58760 50872
rect 58720 50720 58760 50760
rect 57862 50668 58038 50702
rect 58360 50668 58536 50702
rect 57778 50624 57812 50658
rect 58595 50624 58629 50658
rect 57862 50580 58038 50614
rect 58360 50580 58536 50614
rect 57650 50520 57690 50562
rect 58720 50562 58732 50720
rect 58732 50562 58760 50720
rect 58720 50520 58760 50562
rect 62640 51030 62680 51080
rect 62640 50872 62666 51030
rect 62666 50872 62680 51030
rect 63710 51030 63750 51080
rect 62852 50978 63028 51012
rect 63350 50978 63526 51012
rect 62768 50934 62802 50968
rect 63585 50934 63619 50968
rect 62852 50890 63028 50924
rect 63350 50890 63526 50924
rect 62640 50820 62680 50872
rect 62640 50720 62680 50760
rect 62640 50562 62666 50720
rect 62666 50562 62680 50720
rect 63710 50872 63722 51030
rect 63722 50872 63750 51030
rect 63710 50840 63750 50872
rect 63710 50720 63750 50760
rect 62852 50668 63028 50702
rect 63350 50668 63526 50702
rect 62768 50624 62802 50658
rect 63585 50624 63619 50658
rect 62852 50580 63028 50614
rect 63350 50580 63526 50614
rect 62640 50520 62680 50562
rect 63710 50562 63722 50720
rect 63722 50562 63750 50720
rect 63710 50520 63750 50562
rect 67630 51030 67670 51080
rect 67630 50872 67656 51030
rect 67656 50872 67670 51030
rect 68700 51030 68740 51080
rect 67842 50978 68018 51012
rect 68340 50978 68516 51012
rect 67758 50934 67792 50968
rect 68575 50934 68609 50968
rect 67842 50890 68018 50924
rect 68340 50890 68516 50924
rect 67630 50820 67670 50872
rect 67630 50720 67670 50760
rect 67630 50562 67656 50720
rect 67656 50562 67670 50720
rect 68700 50872 68712 51030
rect 68712 50872 68740 51030
rect 68700 50840 68740 50872
rect 68700 50720 68740 50760
rect 67842 50668 68018 50702
rect 68340 50668 68516 50702
rect 67758 50624 67792 50658
rect 68575 50624 68609 50658
rect 67842 50580 68018 50614
rect 68340 50580 68516 50614
rect 67630 50520 67670 50562
rect 68700 50562 68712 50720
rect 68712 50562 68740 50720
rect 68700 50520 68740 50562
rect 72620 51030 72660 51080
rect 72620 50872 72646 51030
rect 72646 50872 72660 51030
rect 73690 51030 73730 51080
rect 72832 50978 73008 51012
rect 73330 50978 73506 51012
rect 72748 50934 72782 50968
rect 73565 50934 73599 50968
rect 72832 50890 73008 50924
rect 73330 50890 73506 50924
rect 72620 50820 72660 50872
rect 72620 50720 72660 50760
rect 72620 50562 72646 50720
rect 72646 50562 72660 50720
rect 73690 50872 73702 51030
rect 73702 50872 73730 51030
rect 73690 50840 73730 50872
rect 73690 50720 73730 50760
rect 72832 50668 73008 50702
rect 73330 50668 73506 50702
rect 72748 50624 72782 50658
rect 73565 50624 73599 50658
rect 72832 50580 73008 50614
rect 73330 50580 73506 50614
rect 72620 50520 72660 50562
rect 73690 50562 73702 50720
rect 73702 50562 73730 50720
rect 73690 50520 73730 50562
rect 77610 51030 77650 51080
rect 77610 50872 77636 51030
rect 77636 50872 77650 51030
rect 78680 51030 78720 51080
rect 77822 50978 77998 51012
rect 78320 50978 78496 51012
rect 77738 50934 77772 50968
rect 78555 50934 78589 50968
rect 77822 50890 77998 50924
rect 78320 50890 78496 50924
rect 77610 50820 77650 50872
rect 77610 50720 77650 50760
rect 77610 50562 77636 50720
rect 77636 50562 77650 50720
rect 78680 50872 78692 51030
rect 78692 50872 78720 51030
rect 78680 50840 78720 50872
rect 78680 50720 78720 50760
rect 77822 50668 77998 50702
rect 78320 50668 78496 50702
rect 77738 50624 77772 50658
rect 78555 50624 78589 50658
rect 77822 50580 77998 50614
rect 78320 50580 78496 50614
rect 77610 50520 77650 50562
rect 78680 50562 78692 50720
rect 78692 50562 78720 50720
rect 78680 50520 78720 50562
rect 2760 49320 2800 49370
rect 2760 49162 2786 49320
rect 2786 49162 2800 49320
rect 3830 49320 3870 49370
rect 2972 49268 3148 49302
rect 3470 49268 3646 49302
rect 2888 49224 2922 49258
rect 3705 49224 3739 49258
rect 2972 49180 3148 49214
rect 3470 49180 3646 49214
rect 2760 49110 2800 49162
rect 2760 49010 2800 49050
rect 2760 48852 2786 49010
rect 2786 48852 2800 49010
rect 3830 49162 3842 49320
rect 3842 49162 3870 49320
rect 3830 49130 3870 49162
rect 3830 49010 3870 49050
rect 2972 48958 3148 48992
rect 3470 48958 3646 48992
rect 2888 48914 2922 48948
rect 3705 48914 3739 48948
rect 2972 48870 3148 48904
rect 3470 48870 3646 48904
rect 2760 48810 2800 48852
rect 3830 48852 3842 49010
rect 3842 48852 3870 49010
rect 3830 48810 3870 48852
rect 7750 49320 7790 49370
rect 7750 49162 7776 49320
rect 7776 49162 7790 49320
rect 8820 49320 8860 49370
rect 7962 49268 8138 49302
rect 8460 49268 8636 49302
rect 7878 49224 7912 49258
rect 8695 49224 8729 49258
rect 7962 49180 8138 49214
rect 8460 49180 8636 49214
rect 7750 49110 7790 49162
rect 7750 49010 7790 49050
rect 7750 48852 7776 49010
rect 7776 48852 7790 49010
rect 8820 49162 8832 49320
rect 8832 49162 8860 49320
rect 8820 49130 8860 49162
rect 8820 49010 8860 49050
rect 7962 48958 8138 48992
rect 8460 48958 8636 48992
rect 7878 48914 7912 48948
rect 8695 48914 8729 48948
rect 7962 48870 8138 48904
rect 8460 48870 8636 48904
rect 7750 48810 7790 48852
rect 8820 48852 8832 49010
rect 8832 48852 8860 49010
rect 8820 48810 8860 48852
rect 12740 49320 12780 49370
rect 12740 49162 12766 49320
rect 12766 49162 12780 49320
rect 13810 49320 13850 49370
rect 12952 49268 13128 49302
rect 13450 49268 13626 49302
rect 12868 49224 12902 49258
rect 13685 49224 13719 49258
rect 12952 49180 13128 49214
rect 13450 49180 13626 49214
rect 12740 49110 12780 49162
rect 12740 49010 12780 49050
rect 12740 48852 12766 49010
rect 12766 48852 12780 49010
rect 13810 49162 13822 49320
rect 13822 49162 13850 49320
rect 13810 49130 13850 49162
rect 13810 49010 13850 49050
rect 12952 48958 13128 48992
rect 13450 48958 13626 48992
rect 12868 48914 12902 48948
rect 13685 48914 13719 48948
rect 12952 48870 13128 48904
rect 13450 48870 13626 48904
rect 12740 48810 12780 48852
rect 13810 48852 13822 49010
rect 13822 48852 13850 49010
rect 13810 48810 13850 48852
rect 17730 49320 17770 49370
rect 17730 49162 17756 49320
rect 17756 49162 17770 49320
rect 18800 49320 18840 49370
rect 17942 49268 18118 49302
rect 18440 49268 18616 49302
rect 17858 49224 17892 49258
rect 18675 49224 18709 49258
rect 17942 49180 18118 49214
rect 18440 49180 18616 49214
rect 17730 49110 17770 49162
rect 17730 49010 17770 49050
rect 17730 48852 17756 49010
rect 17756 48852 17770 49010
rect 18800 49162 18812 49320
rect 18812 49162 18840 49320
rect 18800 49130 18840 49162
rect 18800 49010 18840 49050
rect 17942 48958 18118 48992
rect 18440 48958 18616 48992
rect 17858 48914 17892 48948
rect 18675 48914 18709 48948
rect 17942 48870 18118 48904
rect 18440 48870 18616 48904
rect 17730 48810 17770 48852
rect 18800 48852 18812 49010
rect 18812 48852 18840 49010
rect 18800 48810 18840 48852
rect 22720 49320 22760 49370
rect 22720 49162 22746 49320
rect 22746 49162 22760 49320
rect 23790 49320 23830 49370
rect 22932 49268 23108 49302
rect 23430 49268 23606 49302
rect 22848 49224 22882 49258
rect 23665 49224 23699 49258
rect 22932 49180 23108 49214
rect 23430 49180 23606 49214
rect 22720 49110 22760 49162
rect 22720 49010 22760 49050
rect 22720 48852 22746 49010
rect 22746 48852 22760 49010
rect 23790 49162 23802 49320
rect 23802 49162 23830 49320
rect 23790 49130 23830 49162
rect 23790 49010 23830 49050
rect 22932 48958 23108 48992
rect 23430 48958 23606 48992
rect 22848 48914 22882 48948
rect 23665 48914 23699 48948
rect 22932 48870 23108 48904
rect 23430 48870 23606 48904
rect 22720 48810 22760 48852
rect 23790 48852 23802 49010
rect 23802 48852 23830 49010
rect 23790 48810 23830 48852
rect 27710 49320 27750 49370
rect 27710 49162 27736 49320
rect 27736 49162 27750 49320
rect 28780 49320 28820 49370
rect 27922 49268 28098 49302
rect 28420 49268 28596 49302
rect 27838 49224 27872 49258
rect 28655 49224 28689 49258
rect 27922 49180 28098 49214
rect 28420 49180 28596 49214
rect 27710 49110 27750 49162
rect 27710 49010 27750 49050
rect 27710 48852 27736 49010
rect 27736 48852 27750 49010
rect 28780 49162 28792 49320
rect 28792 49162 28820 49320
rect 28780 49130 28820 49162
rect 28780 49010 28820 49050
rect 27922 48958 28098 48992
rect 28420 48958 28596 48992
rect 27838 48914 27872 48948
rect 28655 48914 28689 48948
rect 27922 48870 28098 48904
rect 28420 48870 28596 48904
rect 27710 48810 27750 48852
rect 28780 48852 28792 49010
rect 28792 48852 28820 49010
rect 28780 48810 28820 48852
rect 32700 49320 32740 49370
rect 32700 49162 32726 49320
rect 32726 49162 32740 49320
rect 33770 49320 33810 49370
rect 32912 49268 33088 49302
rect 33410 49268 33586 49302
rect 32828 49224 32862 49258
rect 33645 49224 33679 49258
rect 32912 49180 33088 49214
rect 33410 49180 33586 49214
rect 32700 49110 32740 49162
rect 32700 49010 32740 49050
rect 32700 48852 32726 49010
rect 32726 48852 32740 49010
rect 33770 49162 33782 49320
rect 33782 49162 33810 49320
rect 33770 49130 33810 49162
rect 33770 49010 33810 49050
rect 32912 48958 33088 48992
rect 33410 48958 33586 48992
rect 32828 48914 32862 48948
rect 33645 48914 33679 48948
rect 32912 48870 33088 48904
rect 33410 48870 33586 48904
rect 32700 48810 32740 48852
rect 33770 48852 33782 49010
rect 33782 48852 33810 49010
rect 33770 48810 33810 48852
rect 37690 49320 37730 49370
rect 37690 49162 37716 49320
rect 37716 49162 37730 49320
rect 38760 49320 38800 49370
rect 37902 49268 38078 49302
rect 38400 49268 38576 49302
rect 37818 49224 37852 49258
rect 38635 49224 38669 49258
rect 37902 49180 38078 49214
rect 38400 49180 38576 49214
rect 37690 49110 37730 49162
rect 37690 49010 37730 49050
rect 37690 48852 37716 49010
rect 37716 48852 37730 49010
rect 38760 49162 38772 49320
rect 38772 49162 38800 49320
rect 38760 49130 38800 49162
rect 38760 49010 38800 49050
rect 37902 48958 38078 48992
rect 38400 48958 38576 48992
rect 37818 48914 37852 48948
rect 38635 48914 38669 48948
rect 37902 48870 38078 48904
rect 38400 48870 38576 48904
rect 37690 48810 37730 48852
rect 38760 48852 38772 49010
rect 38772 48852 38800 49010
rect 38760 48810 38800 48852
rect 42680 49320 42720 49370
rect 42680 49162 42706 49320
rect 42706 49162 42720 49320
rect 43750 49320 43790 49370
rect 42892 49268 43068 49302
rect 43390 49268 43566 49302
rect 42808 49224 42842 49258
rect 43625 49224 43659 49258
rect 42892 49180 43068 49214
rect 43390 49180 43566 49214
rect 42680 49110 42720 49162
rect 42680 49010 42720 49050
rect 42680 48852 42706 49010
rect 42706 48852 42720 49010
rect 43750 49162 43762 49320
rect 43762 49162 43790 49320
rect 43750 49130 43790 49162
rect 43750 49010 43790 49050
rect 42892 48958 43068 48992
rect 43390 48958 43566 48992
rect 42808 48914 42842 48948
rect 43625 48914 43659 48948
rect 42892 48870 43068 48904
rect 43390 48870 43566 48904
rect 42680 48810 42720 48852
rect 43750 48852 43762 49010
rect 43762 48852 43790 49010
rect 43750 48810 43790 48852
rect 47670 49320 47710 49370
rect 47670 49162 47696 49320
rect 47696 49162 47710 49320
rect 48740 49320 48780 49370
rect 47882 49268 48058 49302
rect 48380 49268 48556 49302
rect 47798 49224 47832 49258
rect 48615 49224 48649 49258
rect 47882 49180 48058 49214
rect 48380 49180 48556 49214
rect 47670 49110 47710 49162
rect 47670 49010 47710 49050
rect 47670 48852 47696 49010
rect 47696 48852 47710 49010
rect 48740 49162 48752 49320
rect 48752 49162 48780 49320
rect 48740 49130 48780 49162
rect 48740 49010 48780 49050
rect 47882 48958 48058 48992
rect 48380 48958 48556 48992
rect 47798 48914 47832 48948
rect 48615 48914 48649 48948
rect 47882 48870 48058 48904
rect 48380 48870 48556 48904
rect 47670 48810 47710 48852
rect 48740 48852 48752 49010
rect 48752 48852 48780 49010
rect 48740 48810 48780 48852
rect 52660 49320 52700 49370
rect 52660 49162 52686 49320
rect 52686 49162 52700 49320
rect 53730 49320 53770 49370
rect 52872 49268 53048 49302
rect 53370 49268 53546 49302
rect 52788 49224 52822 49258
rect 53605 49224 53639 49258
rect 52872 49180 53048 49214
rect 53370 49180 53546 49214
rect 52660 49110 52700 49162
rect 52660 49010 52700 49050
rect 52660 48852 52686 49010
rect 52686 48852 52700 49010
rect 53730 49162 53742 49320
rect 53742 49162 53770 49320
rect 53730 49130 53770 49162
rect 53730 49010 53770 49050
rect 52872 48958 53048 48992
rect 53370 48958 53546 48992
rect 52788 48914 52822 48948
rect 53605 48914 53639 48948
rect 52872 48870 53048 48904
rect 53370 48870 53546 48904
rect 52660 48810 52700 48852
rect 53730 48852 53742 49010
rect 53742 48852 53770 49010
rect 53730 48810 53770 48852
rect 57650 49320 57690 49370
rect 57650 49162 57676 49320
rect 57676 49162 57690 49320
rect 58720 49320 58760 49370
rect 57862 49268 58038 49302
rect 58360 49268 58536 49302
rect 57778 49224 57812 49258
rect 58595 49224 58629 49258
rect 57862 49180 58038 49214
rect 58360 49180 58536 49214
rect 57650 49110 57690 49162
rect 57650 49010 57690 49050
rect 57650 48852 57676 49010
rect 57676 48852 57690 49010
rect 58720 49162 58732 49320
rect 58732 49162 58760 49320
rect 58720 49130 58760 49162
rect 58720 49010 58760 49050
rect 57862 48958 58038 48992
rect 58360 48958 58536 48992
rect 57778 48914 57812 48948
rect 58595 48914 58629 48948
rect 57862 48870 58038 48904
rect 58360 48870 58536 48904
rect 57650 48810 57690 48852
rect 58720 48852 58732 49010
rect 58732 48852 58760 49010
rect 58720 48810 58760 48852
rect 62640 49320 62680 49370
rect 62640 49162 62666 49320
rect 62666 49162 62680 49320
rect 63710 49320 63750 49370
rect 62852 49268 63028 49302
rect 63350 49268 63526 49302
rect 62768 49224 62802 49258
rect 63585 49224 63619 49258
rect 62852 49180 63028 49214
rect 63350 49180 63526 49214
rect 62640 49110 62680 49162
rect 62640 49010 62680 49050
rect 62640 48852 62666 49010
rect 62666 48852 62680 49010
rect 63710 49162 63722 49320
rect 63722 49162 63750 49320
rect 63710 49130 63750 49162
rect 63710 49010 63750 49050
rect 62852 48958 63028 48992
rect 63350 48958 63526 48992
rect 62768 48914 62802 48948
rect 63585 48914 63619 48948
rect 62852 48870 63028 48904
rect 63350 48870 63526 48904
rect 62640 48810 62680 48852
rect 63710 48852 63722 49010
rect 63722 48852 63750 49010
rect 63710 48810 63750 48852
rect 67630 49320 67670 49370
rect 67630 49162 67656 49320
rect 67656 49162 67670 49320
rect 68700 49320 68740 49370
rect 67842 49268 68018 49302
rect 68340 49268 68516 49302
rect 67758 49224 67792 49258
rect 68575 49224 68609 49258
rect 67842 49180 68018 49214
rect 68340 49180 68516 49214
rect 67630 49110 67670 49162
rect 67630 49010 67670 49050
rect 67630 48852 67656 49010
rect 67656 48852 67670 49010
rect 68700 49162 68712 49320
rect 68712 49162 68740 49320
rect 68700 49130 68740 49162
rect 68700 49010 68740 49050
rect 67842 48958 68018 48992
rect 68340 48958 68516 48992
rect 67758 48914 67792 48948
rect 68575 48914 68609 48948
rect 67842 48870 68018 48904
rect 68340 48870 68516 48904
rect 67630 48810 67670 48852
rect 68700 48852 68712 49010
rect 68712 48852 68740 49010
rect 68700 48810 68740 48852
rect 72620 49320 72660 49370
rect 72620 49162 72646 49320
rect 72646 49162 72660 49320
rect 73690 49320 73730 49370
rect 72832 49268 73008 49302
rect 73330 49268 73506 49302
rect 72748 49224 72782 49258
rect 73565 49224 73599 49258
rect 72832 49180 73008 49214
rect 73330 49180 73506 49214
rect 72620 49110 72660 49162
rect 72620 49010 72660 49050
rect 72620 48852 72646 49010
rect 72646 48852 72660 49010
rect 73690 49162 73702 49320
rect 73702 49162 73730 49320
rect 73690 49130 73730 49162
rect 73690 49010 73730 49050
rect 72832 48958 73008 48992
rect 73330 48958 73506 48992
rect 72748 48914 72782 48948
rect 73565 48914 73599 48948
rect 72832 48870 73008 48904
rect 73330 48870 73506 48904
rect 72620 48810 72660 48852
rect 73690 48852 73702 49010
rect 73702 48852 73730 49010
rect 73690 48810 73730 48852
rect 77610 49320 77650 49370
rect 77610 49162 77636 49320
rect 77636 49162 77650 49320
rect 78680 49320 78720 49370
rect 77822 49268 77998 49302
rect 78320 49268 78496 49302
rect 77738 49224 77772 49258
rect 78555 49224 78589 49258
rect 77822 49180 77998 49214
rect 78320 49180 78496 49214
rect 77610 49110 77650 49162
rect 77610 49010 77650 49050
rect 77610 48852 77636 49010
rect 77636 48852 77650 49010
rect 78680 49162 78692 49320
rect 78692 49162 78720 49320
rect 78680 49130 78720 49162
rect 78680 49010 78720 49050
rect 77822 48958 77998 48992
rect 78320 48958 78496 48992
rect 77738 48914 77772 48948
rect 78555 48914 78589 48948
rect 77822 48870 77998 48904
rect 78320 48870 78496 48904
rect 77610 48810 77650 48852
rect 78680 48852 78692 49010
rect 78692 48852 78720 49010
rect 78680 48810 78720 48852
rect 2760 47610 2800 47660
rect 2760 47452 2786 47610
rect 2786 47452 2800 47610
rect 3830 47610 3870 47660
rect 2972 47558 3148 47592
rect 3470 47558 3646 47592
rect 2888 47514 2922 47548
rect 3705 47514 3739 47548
rect 2972 47470 3148 47504
rect 3470 47470 3646 47504
rect 2760 47400 2800 47452
rect 2760 47300 2800 47340
rect 2760 47142 2786 47300
rect 2786 47142 2800 47300
rect 3830 47452 3842 47610
rect 3842 47452 3870 47610
rect 3830 47420 3870 47452
rect 3830 47300 3870 47340
rect 2972 47248 3148 47282
rect 3470 47248 3646 47282
rect 2888 47204 2922 47238
rect 3705 47204 3739 47238
rect 2972 47160 3148 47194
rect 3470 47160 3646 47194
rect 2760 47100 2800 47142
rect 3830 47142 3842 47300
rect 3842 47142 3870 47300
rect 3830 47100 3870 47142
rect 7750 47610 7790 47660
rect 7750 47452 7776 47610
rect 7776 47452 7790 47610
rect 8820 47610 8860 47660
rect 7962 47558 8138 47592
rect 8460 47558 8636 47592
rect 7878 47514 7912 47548
rect 8695 47514 8729 47548
rect 7962 47470 8138 47504
rect 8460 47470 8636 47504
rect 7750 47400 7790 47452
rect 7750 47300 7790 47340
rect 7750 47142 7776 47300
rect 7776 47142 7790 47300
rect 8820 47452 8832 47610
rect 8832 47452 8860 47610
rect 8820 47420 8860 47452
rect 8820 47300 8860 47340
rect 7962 47248 8138 47282
rect 8460 47248 8636 47282
rect 7878 47204 7912 47238
rect 8695 47204 8729 47238
rect 7962 47160 8138 47194
rect 8460 47160 8636 47194
rect 7750 47100 7790 47142
rect 8820 47142 8832 47300
rect 8832 47142 8860 47300
rect 8820 47100 8860 47142
rect 12740 47610 12780 47660
rect 12740 47452 12766 47610
rect 12766 47452 12780 47610
rect 13810 47610 13850 47660
rect 12952 47558 13128 47592
rect 13450 47558 13626 47592
rect 12868 47514 12902 47548
rect 13685 47514 13719 47548
rect 12952 47470 13128 47504
rect 13450 47470 13626 47504
rect 12740 47400 12780 47452
rect 12740 47300 12780 47340
rect 12740 47142 12766 47300
rect 12766 47142 12780 47300
rect 13810 47452 13822 47610
rect 13822 47452 13850 47610
rect 13810 47420 13850 47452
rect 13810 47300 13850 47340
rect 12952 47248 13128 47282
rect 13450 47248 13626 47282
rect 12868 47204 12902 47238
rect 13685 47204 13719 47238
rect 12952 47160 13128 47194
rect 13450 47160 13626 47194
rect 12740 47100 12780 47142
rect 13810 47142 13822 47300
rect 13822 47142 13850 47300
rect 13810 47100 13850 47142
rect 17730 47610 17770 47660
rect 17730 47452 17756 47610
rect 17756 47452 17770 47610
rect 18800 47610 18840 47660
rect 17942 47558 18118 47592
rect 18440 47558 18616 47592
rect 17858 47514 17892 47548
rect 18675 47514 18709 47548
rect 17942 47470 18118 47504
rect 18440 47470 18616 47504
rect 17730 47400 17770 47452
rect 17730 47300 17770 47340
rect 17730 47142 17756 47300
rect 17756 47142 17770 47300
rect 18800 47452 18812 47610
rect 18812 47452 18840 47610
rect 18800 47420 18840 47452
rect 18800 47300 18840 47340
rect 17942 47248 18118 47282
rect 18440 47248 18616 47282
rect 17858 47204 17892 47238
rect 18675 47204 18709 47238
rect 17942 47160 18118 47194
rect 18440 47160 18616 47194
rect 17730 47100 17770 47142
rect 18800 47142 18812 47300
rect 18812 47142 18840 47300
rect 18800 47100 18840 47142
rect 22720 47610 22760 47660
rect 22720 47452 22746 47610
rect 22746 47452 22760 47610
rect 23790 47610 23830 47660
rect 22932 47558 23108 47592
rect 23430 47558 23606 47592
rect 22848 47514 22882 47548
rect 23665 47514 23699 47548
rect 22932 47470 23108 47504
rect 23430 47470 23606 47504
rect 22720 47400 22760 47452
rect 22720 47300 22760 47340
rect 22720 47142 22746 47300
rect 22746 47142 22760 47300
rect 23790 47452 23802 47610
rect 23802 47452 23830 47610
rect 23790 47420 23830 47452
rect 23790 47300 23830 47340
rect 22932 47248 23108 47282
rect 23430 47248 23606 47282
rect 22848 47204 22882 47238
rect 23665 47204 23699 47238
rect 22932 47160 23108 47194
rect 23430 47160 23606 47194
rect 22720 47100 22760 47142
rect 23790 47142 23802 47300
rect 23802 47142 23830 47300
rect 23790 47100 23830 47142
rect 27710 47610 27750 47660
rect 27710 47452 27736 47610
rect 27736 47452 27750 47610
rect 28780 47610 28820 47660
rect 27922 47558 28098 47592
rect 28420 47558 28596 47592
rect 27838 47514 27872 47548
rect 28655 47514 28689 47548
rect 27922 47470 28098 47504
rect 28420 47470 28596 47504
rect 27710 47400 27750 47452
rect 27710 47300 27750 47340
rect 27710 47142 27736 47300
rect 27736 47142 27750 47300
rect 28780 47452 28792 47610
rect 28792 47452 28820 47610
rect 28780 47420 28820 47452
rect 28780 47300 28820 47340
rect 27922 47248 28098 47282
rect 28420 47248 28596 47282
rect 27838 47204 27872 47238
rect 28655 47204 28689 47238
rect 27922 47160 28098 47194
rect 28420 47160 28596 47194
rect 27710 47100 27750 47142
rect 28780 47142 28792 47300
rect 28792 47142 28820 47300
rect 28780 47100 28820 47142
rect 32700 47610 32740 47660
rect 32700 47452 32726 47610
rect 32726 47452 32740 47610
rect 33770 47610 33810 47660
rect 32912 47558 33088 47592
rect 33410 47558 33586 47592
rect 32828 47514 32862 47548
rect 33645 47514 33679 47548
rect 32912 47470 33088 47504
rect 33410 47470 33586 47504
rect 32700 47400 32740 47452
rect 32700 47300 32740 47340
rect 32700 47142 32726 47300
rect 32726 47142 32740 47300
rect 33770 47452 33782 47610
rect 33782 47452 33810 47610
rect 33770 47420 33810 47452
rect 33770 47300 33810 47340
rect 32912 47248 33088 47282
rect 33410 47248 33586 47282
rect 32828 47204 32862 47238
rect 33645 47204 33679 47238
rect 32912 47160 33088 47194
rect 33410 47160 33586 47194
rect 32700 47100 32740 47142
rect 33770 47142 33782 47300
rect 33782 47142 33810 47300
rect 33770 47100 33810 47142
rect 37690 47610 37730 47660
rect 37690 47452 37716 47610
rect 37716 47452 37730 47610
rect 38760 47610 38800 47660
rect 37902 47558 38078 47592
rect 38400 47558 38576 47592
rect 37818 47514 37852 47548
rect 38635 47514 38669 47548
rect 37902 47470 38078 47504
rect 38400 47470 38576 47504
rect 37690 47400 37730 47452
rect 37690 47300 37730 47340
rect 37690 47142 37716 47300
rect 37716 47142 37730 47300
rect 38760 47452 38772 47610
rect 38772 47452 38800 47610
rect 38760 47420 38800 47452
rect 38760 47300 38800 47340
rect 37902 47248 38078 47282
rect 38400 47248 38576 47282
rect 37818 47204 37852 47238
rect 38635 47204 38669 47238
rect 37902 47160 38078 47194
rect 38400 47160 38576 47194
rect 37690 47100 37730 47142
rect 38760 47142 38772 47300
rect 38772 47142 38800 47300
rect 38760 47100 38800 47142
rect 42680 47610 42720 47660
rect 42680 47452 42706 47610
rect 42706 47452 42720 47610
rect 43750 47610 43790 47660
rect 42892 47558 43068 47592
rect 43390 47558 43566 47592
rect 42808 47514 42842 47548
rect 43625 47514 43659 47548
rect 42892 47470 43068 47504
rect 43390 47470 43566 47504
rect 42680 47400 42720 47452
rect 42680 47300 42720 47340
rect 42680 47142 42706 47300
rect 42706 47142 42720 47300
rect 43750 47452 43762 47610
rect 43762 47452 43790 47610
rect 43750 47420 43790 47452
rect 43750 47300 43790 47340
rect 42892 47248 43068 47282
rect 43390 47248 43566 47282
rect 42808 47204 42842 47238
rect 43625 47204 43659 47238
rect 42892 47160 43068 47194
rect 43390 47160 43566 47194
rect 42680 47100 42720 47142
rect 43750 47142 43762 47300
rect 43762 47142 43790 47300
rect 43750 47100 43790 47142
rect 47670 47610 47710 47660
rect 47670 47452 47696 47610
rect 47696 47452 47710 47610
rect 48740 47610 48780 47660
rect 47882 47558 48058 47592
rect 48380 47558 48556 47592
rect 47798 47514 47832 47548
rect 48615 47514 48649 47548
rect 47882 47470 48058 47504
rect 48380 47470 48556 47504
rect 47670 47400 47710 47452
rect 47670 47300 47710 47340
rect 47670 47142 47696 47300
rect 47696 47142 47710 47300
rect 48740 47452 48752 47610
rect 48752 47452 48780 47610
rect 48740 47420 48780 47452
rect 48740 47300 48780 47340
rect 47882 47248 48058 47282
rect 48380 47248 48556 47282
rect 47798 47204 47832 47238
rect 48615 47204 48649 47238
rect 47882 47160 48058 47194
rect 48380 47160 48556 47194
rect 47670 47100 47710 47142
rect 48740 47142 48752 47300
rect 48752 47142 48780 47300
rect 48740 47100 48780 47142
rect 52660 47610 52700 47660
rect 52660 47452 52686 47610
rect 52686 47452 52700 47610
rect 53730 47610 53770 47660
rect 52872 47558 53048 47592
rect 53370 47558 53546 47592
rect 52788 47514 52822 47548
rect 53605 47514 53639 47548
rect 52872 47470 53048 47504
rect 53370 47470 53546 47504
rect 52660 47400 52700 47452
rect 52660 47300 52700 47340
rect 52660 47142 52686 47300
rect 52686 47142 52700 47300
rect 53730 47452 53742 47610
rect 53742 47452 53770 47610
rect 53730 47420 53770 47452
rect 53730 47300 53770 47340
rect 52872 47248 53048 47282
rect 53370 47248 53546 47282
rect 52788 47204 52822 47238
rect 53605 47204 53639 47238
rect 52872 47160 53048 47194
rect 53370 47160 53546 47194
rect 52660 47100 52700 47142
rect 53730 47142 53742 47300
rect 53742 47142 53770 47300
rect 53730 47100 53770 47142
rect 57650 47610 57690 47660
rect 57650 47452 57676 47610
rect 57676 47452 57690 47610
rect 58720 47610 58760 47660
rect 57862 47558 58038 47592
rect 58360 47558 58536 47592
rect 57778 47514 57812 47548
rect 58595 47514 58629 47548
rect 57862 47470 58038 47504
rect 58360 47470 58536 47504
rect 57650 47400 57690 47452
rect 57650 47300 57690 47340
rect 57650 47142 57676 47300
rect 57676 47142 57690 47300
rect 58720 47452 58732 47610
rect 58732 47452 58760 47610
rect 58720 47420 58760 47452
rect 58720 47300 58760 47340
rect 57862 47248 58038 47282
rect 58360 47248 58536 47282
rect 57778 47204 57812 47238
rect 58595 47204 58629 47238
rect 57862 47160 58038 47194
rect 58360 47160 58536 47194
rect 57650 47100 57690 47142
rect 58720 47142 58732 47300
rect 58732 47142 58760 47300
rect 58720 47100 58760 47142
rect 62640 47610 62680 47660
rect 62640 47452 62666 47610
rect 62666 47452 62680 47610
rect 63710 47610 63750 47660
rect 62852 47558 63028 47592
rect 63350 47558 63526 47592
rect 62768 47514 62802 47548
rect 63585 47514 63619 47548
rect 62852 47470 63028 47504
rect 63350 47470 63526 47504
rect 62640 47400 62680 47452
rect 62640 47300 62680 47340
rect 62640 47142 62666 47300
rect 62666 47142 62680 47300
rect 63710 47452 63722 47610
rect 63722 47452 63750 47610
rect 63710 47420 63750 47452
rect 63710 47300 63750 47340
rect 62852 47248 63028 47282
rect 63350 47248 63526 47282
rect 62768 47204 62802 47238
rect 63585 47204 63619 47238
rect 62852 47160 63028 47194
rect 63350 47160 63526 47194
rect 62640 47100 62680 47142
rect 63710 47142 63722 47300
rect 63722 47142 63750 47300
rect 63710 47100 63750 47142
rect 67630 47610 67670 47660
rect 67630 47452 67656 47610
rect 67656 47452 67670 47610
rect 68700 47610 68740 47660
rect 67842 47558 68018 47592
rect 68340 47558 68516 47592
rect 67758 47514 67792 47548
rect 68575 47514 68609 47548
rect 67842 47470 68018 47504
rect 68340 47470 68516 47504
rect 67630 47400 67670 47452
rect 67630 47300 67670 47340
rect 67630 47142 67656 47300
rect 67656 47142 67670 47300
rect 68700 47452 68712 47610
rect 68712 47452 68740 47610
rect 68700 47420 68740 47452
rect 68700 47300 68740 47340
rect 67842 47248 68018 47282
rect 68340 47248 68516 47282
rect 67758 47204 67792 47238
rect 68575 47204 68609 47238
rect 67842 47160 68018 47194
rect 68340 47160 68516 47194
rect 67630 47100 67670 47142
rect 68700 47142 68712 47300
rect 68712 47142 68740 47300
rect 68700 47100 68740 47142
rect 72620 47610 72660 47660
rect 72620 47452 72646 47610
rect 72646 47452 72660 47610
rect 73690 47610 73730 47660
rect 72832 47558 73008 47592
rect 73330 47558 73506 47592
rect 72748 47514 72782 47548
rect 73565 47514 73599 47548
rect 72832 47470 73008 47504
rect 73330 47470 73506 47504
rect 72620 47400 72660 47452
rect 72620 47300 72660 47340
rect 72620 47142 72646 47300
rect 72646 47142 72660 47300
rect 73690 47452 73702 47610
rect 73702 47452 73730 47610
rect 73690 47420 73730 47452
rect 73690 47300 73730 47340
rect 72832 47248 73008 47282
rect 73330 47248 73506 47282
rect 72748 47204 72782 47238
rect 73565 47204 73599 47238
rect 72832 47160 73008 47194
rect 73330 47160 73506 47194
rect 72620 47100 72660 47142
rect 73690 47142 73702 47300
rect 73702 47142 73730 47300
rect 73690 47100 73730 47142
rect 77610 47610 77650 47660
rect 77610 47452 77636 47610
rect 77636 47452 77650 47610
rect 78680 47610 78720 47660
rect 77822 47558 77998 47592
rect 78320 47558 78496 47592
rect 77738 47514 77772 47548
rect 78555 47514 78589 47548
rect 77822 47470 77998 47504
rect 78320 47470 78496 47504
rect 77610 47400 77650 47452
rect 77610 47300 77650 47340
rect 77610 47142 77636 47300
rect 77636 47142 77650 47300
rect 78680 47452 78692 47610
rect 78692 47452 78720 47610
rect 78680 47420 78720 47452
rect 78680 47300 78720 47340
rect 77822 47248 77998 47282
rect 78320 47248 78496 47282
rect 77738 47204 77772 47238
rect 78555 47204 78589 47238
rect 77822 47160 77998 47194
rect 78320 47160 78496 47194
rect 77610 47100 77650 47142
rect 78680 47142 78692 47300
rect 78692 47142 78720 47300
rect 78680 47100 78720 47142
rect 2760 45900 2800 45950
rect 2760 45742 2786 45900
rect 2786 45742 2800 45900
rect 3830 45900 3870 45950
rect 2972 45848 3148 45882
rect 3470 45848 3646 45882
rect 2888 45804 2922 45838
rect 3705 45804 3739 45838
rect 2972 45760 3148 45794
rect 3470 45760 3646 45794
rect 2760 45690 2800 45742
rect 2760 45590 2800 45630
rect 2760 45432 2786 45590
rect 2786 45432 2800 45590
rect 3830 45742 3842 45900
rect 3842 45742 3870 45900
rect 3830 45710 3870 45742
rect 3830 45590 3870 45630
rect 2972 45538 3148 45572
rect 3470 45538 3646 45572
rect 2888 45494 2922 45528
rect 3705 45494 3739 45528
rect 2972 45450 3148 45484
rect 3470 45450 3646 45484
rect 2760 45390 2800 45432
rect 3830 45432 3842 45590
rect 3842 45432 3870 45590
rect 3830 45390 3870 45432
rect 7750 45900 7790 45950
rect 7750 45742 7776 45900
rect 7776 45742 7790 45900
rect 8820 45900 8860 45950
rect 7962 45848 8138 45882
rect 8460 45848 8636 45882
rect 7878 45804 7912 45838
rect 8695 45804 8729 45838
rect 7962 45760 8138 45794
rect 8460 45760 8636 45794
rect 7750 45690 7790 45742
rect 7750 45590 7790 45630
rect 7750 45432 7776 45590
rect 7776 45432 7790 45590
rect 8820 45742 8832 45900
rect 8832 45742 8860 45900
rect 8820 45710 8860 45742
rect 8820 45590 8860 45630
rect 7962 45538 8138 45572
rect 8460 45538 8636 45572
rect 7878 45494 7912 45528
rect 8695 45494 8729 45528
rect 7962 45450 8138 45484
rect 8460 45450 8636 45484
rect 7750 45390 7790 45432
rect 8820 45432 8832 45590
rect 8832 45432 8860 45590
rect 8820 45390 8860 45432
rect 12740 45900 12780 45950
rect 12740 45742 12766 45900
rect 12766 45742 12780 45900
rect 13810 45900 13850 45950
rect 12952 45848 13128 45882
rect 13450 45848 13626 45882
rect 12868 45804 12902 45838
rect 13685 45804 13719 45838
rect 12952 45760 13128 45794
rect 13450 45760 13626 45794
rect 12740 45690 12780 45742
rect 12740 45590 12780 45630
rect 12740 45432 12766 45590
rect 12766 45432 12780 45590
rect 13810 45742 13822 45900
rect 13822 45742 13850 45900
rect 13810 45710 13850 45742
rect 13810 45590 13850 45630
rect 12952 45538 13128 45572
rect 13450 45538 13626 45572
rect 12868 45494 12902 45528
rect 13685 45494 13719 45528
rect 12952 45450 13128 45484
rect 13450 45450 13626 45484
rect 12740 45390 12780 45432
rect 13810 45432 13822 45590
rect 13822 45432 13850 45590
rect 13810 45390 13850 45432
rect 17730 45900 17770 45950
rect 17730 45742 17756 45900
rect 17756 45742 17770 45900
rect 18800 45900 18840 45950
rect 17942 45848 18118 45882
rect 18440 45848 18616 45882
rect 17858 45804 17892 45838
rect 18675 45804 18709 45838
rect 17942 45760 18118 45794
rect 18440 45760 18616 45794
rect 17730 45690 17770 45742
rect 17730 45590 17770 45630
rect 17730 45432 17756 45590
rect 17756 45432 17770 45590
rect 18800 45742 18812 45900
rect 18812 45742 18840 45900
rect 18800 45710 18840 45742
rect 18800 45590 18840 45630
rect 17942 45538 18118 45572
rect 18440 45538 18616 45572
rect 17858 45494 17892 45528
rect 18675 45494 18709 45528
rect 17942 45450 18118 45484
rect 18440 45450 18616 45484
rect 17730 45390 17770 45432
rect 18800 45432 18812 45590
rect 18812 45432 18840 45590
rect 18800 45390 18840 45432
rect 22720 45900 22760 45950
rect 22720 45742 22746 45900
rect 22746 45742 22760 45900
rect 23790 45900 23830 45950
rect 22932 45848 23108 45882
rect 23430 45848 23606 45882
rect 22848 45804 22882 45838
rect 23665 45804 23699 45838
rect 22932 45760 23108 45794
rect 23430 45760 23606 45794
rect 22720 45690 22760 45742
rect 22720 45590 22760 45630
rect 22720 45432 22746 45590
rect 22746 45432 22760 45590
rect 23790 45742 23802 45900
rect 23802 45742 23830 45900
rect 23790 45710 23830 45742
rect 23790 45590 23830 45630
rect 22932 45538 23108 45572
rect 23430 45538 23606 45572
rect 22848 45494 22882 45528
rect 23665 45494 23699 45528
rect 22932 45450 23108 45484
rect 23430 45450 23606 45484
rect 22720 45390 22760 45432
rect 23790 45432 23802 45590
rect 23802 45432 23830 45590
rect 23790 45390 23830 45432
rect 27710 45900 27750 45950
rect 27710 45742 27736 45900
rect 27736 45742 27750 45900
rect 28780 45900 28820 45950
rect 27922 45848 28098 45882
rect 28420 45848 28596 45882
rect 27838 45804 27872 45838
rect 28655 45804 28689 45838
rect 27922 45760 28098 45794
rect 28420 45760 28596 45794
rect 27710 45690 27750 45742
rect 27710 45590 27750 45630
rect 27710 45432 27736 45590
rect 27736 45432 27750 45590
rect 28780 45742 28792 45900
rect 28792 45742 28820 45900
rect 28780 45710 28820 45742
rect 28780 45590 28820 45630
rect 27922 45538 28098 45572
rect 28420 45538 28596 45572
rect 27838 45494 27872 45528
rect 28655 45494 28689 45528
rect 27922 45450 28098 45484
rect 28420 45450 28596 45484
rect 27710 45390 27750 45432
rect 28780 45432 28792 45590
rect 28792 45432 28820 45590
rect 28780 45390 28820 45432
rect 32700 45900 32740 45950
rect 32700 45742 32726 45900
rect 32726 45742 32740 45900
rect 33770 45900 33810 45950
rect 32912 45848 33088 45882
rect 33410 45848 33586 45882
rect 32828 45804 32862 45838
rect 33645 45804 33679 45838
rect 32912 45760 33088 45794
rect 33410 45760 33586 45794
rect 32700 45690 32740 45742
rect 32700 45590 32740 45630
rect 32700 45432 32726 45590
rect 32726 45432 32740 45590
rect 33770 45742 33782 45900
rect 33782 45742 33810 45900
rect 33770 45710 33810 45742
rect 33770 45590 33810 45630
rect 32912 45538 33088 45572
rect 33410 45538 33586 45572
rect 32828 45494 32862 45528
rect 33645 45494 33679 45528
rect 32912 45450 33088 45484
rect 33410 45450 33586 45484
rect 32700 45390 32740 45432
rect 33770 45432 33782 45590
rect 33782 45432 33810 45590
rect 33770 45390 33810 45432
rect 37690 45900 37730 45950
rect 37690 45742 37716 45900
rect 37716 45742 37730 45900
rect 38760 45900 38800 45950
rect 37902 45848 38078 45882
rect 38400 45848 38576 45882
rect 37818 45804 37852 45838
rect 38635 45804 38669 45838
rect 37902 45760 38078 45794
rect 38400 45760 38576 45794
rect 37690 45690 37730 45742
rect 37690 45590 37730 45630
rect 37690 45432 37716 45590
rect 37716 45432 37730 45590
rect 38760 45742 38772 45900
rect 38772 45742 38800 45900
rect 38760 45710 38800 45742
rect 38760 45590 38800 45630
rect 37902 45538 38078 45572
rect 38400 45538 38576 45572
rect 37818 45494 37852 45528
rect 38635 45494 38669 45528
rect 37902 45450 38078 45484
rect 38400 45450 38576 45484
rect 37690 45390 37730 45432
rect 38760 45432 38772 45590
rect 38772 45432 38800 45590
rect 38760 45390 38800 45432
rect 42680 45900 42720 45950
rect 42680 45742 42706 45900
rect 42706 45742 42720 45900
rect 43750 45900 43790 45950
rect 42892 45848 43068 45882
rect 43390 45848 43566 45882
rect 42808 45804 42842 45838
rect 43625 45804 43659 45838
rect 42892 45760 43068 45794
rect 43390 45760 43566 45794
rect 42680 45690 42720 45742
rect 42680 45590 42720 45630
rect 42680 45432 42706 45590
rect 42706 45432 42720 45590
rect 43750 45742 43762 45900
rect 43762 45742 43790 45900
rect 43750 45710 43790 45742
rect 43750 45590 43790 45630
rect 42892 45538 43068 45572
rect 43390 45538 43566 45572
rect 42808 45494 42842 45528
rect 43625 45494 43659 45528
rect 42892 45450 43068 45484
rect 43390 45450 43566 45484
rect 42680 45390 42720 45432
rect 43750 45432 43762 45590
rect 43762 45432 43790 45590
rect 43750 45390 43790 45432
rect 47670 45900 47710 45950
rect 47670 45742 47696 45900
rect 47696 45742 47710 45900
rect 48740 45900 48780 45950
rect 47882 45848 48058 45882
rect 48380 45848 48556 45882
rect 47798 45804 47832 45838
rect 48615 45804 48649 45838
rect 47882 45760 48058 45794
rect 48380 45760 48556 45794
rect 47670 45690 47710 45742
rect 47670 45590 47710 45630
rect 47670 45432 47696 45590
rect 47696 45432 47710 45590
rect 48740 45742 48752 45900
rect 48752 45742 48780 45900
rect 48740 45710 48780 45742
rect 48740 45590 48780 45630
rect 47882 45538 48058 45572
rect 48380 45538 48556 45572
rect 47798 45494 47832 45528
rect 48615 45494 48649 45528
rect 47882 45450 48058 45484
rect 48380 45450 48556 45484
rect 47670 45390 47710 45432
rect 48740 45432 48752 45590
rect 48752 45432 48780 45590
rect 48740 45390 48780 45432
rect 52660 45900 52700 45950
rect 52660 45742 52686 45900
rect 52686 45742 52700 45900
rect 53730 45900 53770 45950
rect 52872 45848 53048 45882
rect 53370 45848 53546 45882
rect 52788 45804 52822 45838
rect 53605 45804 53639 45838
rect 52872 45760 53048 45794
rect 53370 45760 53546 45794
rect 52660 45690 52700 45742
rect 52660 45590 52700 45630
rect 52660 45432 52686 45590
rect 52686 45432 52700 45590
rect 53730 45742 53742 45900
rect 53742 45742 53770 45900
rect 53730 45710 53770 45742
rect 53730 45590 53770 45630
rect 52872 45538 53048 45572
rect 53370 45538 53546 45572
rect 52788 45494 52822 45528
rect 53605 45494 53639 45528
rect 52872 45450 53048 45484
rect 53370 45450 53546 45484
rect 52660 45390 52700 45432
rect 53730 45432 53742 45590
rect 53742 45432 53770 45590
rect 53730 45390 53770 45432
rect 57650 45900 57690 45950
rect 57650 45742 57676 45900
rect 57676 45742 57690 45900
rect 58720 45900 58760 45950
rect 57862 45848 58038 45882
rect 58360 45848 58536 45882
rect 57778 45804 57812 45838
rect 58595 45804 58629 45838
rect 57862 45760 58038 45794
rect 58360 45760 58536 45794
rect 57650 45690 57690 45742
rect 57650 45590 57690 45630
rect 57650 45432 57676 45590
rect 57676 45432 57690 45590
rect 58720 45742 58732 45900
rect 58732 45742 58760 45900
rect 58720 45710 58760 45742
rect 58720 45590 58760 45630
rect 57862 45538 58038 45572
rect 58360 45538 58536 45572
rect 57778 45494 57812 45528
rect 58595 45494 58629 45528
rect 57862 45450 58038 45484
rect 58360 45450 58536 45484
rect 57650 45390 57690 45432
rect 58720 45432 58732 45590
rect 58732 45432 58760 45590
rect 58720 45390 58760 45432
rect 62640 45900 62680 45950
rect 62640 45742 62666 45900
rect 62666 45742 62680 45900
rect 63710 45900 63750 45950
rect 62852 45848 63028 45882
rect 63350 45848 63526 45882
rect 62768 45804 62802 45838
rect 63585 45804 63619 45838
rect 62852 45760 63028 45794
rect 63350 45760 63526 45794
rect 62640 45690 62680 45742
rect 62640 45590 62680 45630
rect 62640 45432 62666 45590
rect 62666 45432 62680 45590
rect 63710 45742 63722 45900
rect 63722 45742 63750 45900
rect 63710 45710 63750 45742
rect 63710 45590 63750 45630
rect 62852 45538 63028 45572
rect 63350 45538 63526 45572
rect 62768 45494 62802 45528
rect 63585 45494 63619 45528
rect 62852 45450 63028 45484
rect 63350 45450 63526 45484
rect 62640 45390 62680 45432
rect 63710 45432 63722 45590
rect 63722 45432 63750 45590
rect 63710 45390 63750 45432
rect 67630 45900 67670 45950
rect 67630 45742 67656 45900
rect 67656 45742 67670 45900
rect 68700 45900 68740 45950
rect 67842 45848 68018 45882
rect 68340 45848 68516 45882
rect 67758 45804 67792 45838
rect 68575 45804 68609 45838
rect 67842 45760 68018 45794
rect 68340 45760 68516 45794
rect 67630 45690 67670 45742
rect 67630 45590 67670 45630
rect 67630 45432 67656 45590
rect 67656 45432 67670 45590
rect 68700 45742 68712 45900
rect 68712 45742 68740 45900
rect 68700 45710 68740 45742
rect 68700 45590 68740 45630
rect 67842 45538 68018 45572
rect 68340 45538 68516 45572
rect 67758 45494 67792 45528
rect 68575 45494 68609 45528
rect 67842 45450 68018 45484
rect 68340 45450 68516 45484
rect 67630 45390 67670 45432
rect 68700 45432 68712 45590
rect 68712 45432 68740 45590
rect 68700 45390 68740 45432
rect 72620 45900 72660 45950
rect 72620 45742 72646 45900
rect 72646 45742 72660 45900
rect 73690 45900 73730 45950
rect 72832 45848 73008 45882
rect 73330 45848 73506 45882
rect 72748 45804 72782 45838
rect 73565 45804 73599 45838
rect 72832 45760 73008 45794
rect 73330 45760 73506 45794
rect 72620 45690 72660 45742
rect 72620 45590 72660 45630
rect 72620 45432 72646 45590
rect 72646 45432 72660 45590
rect 73690 45742 73702 45900
rect 73702 45742 73730 45900
rect 73690 45710 73730 45742
rect 73690 45590 73730 45630
rect 72832 45538 73008 45572
rect 73330 45538 73506 45572
rect 72748 45494 72782 45528
rect 73565 45494 73599 45528
rect 72832 45450 73008 45484
rect 73330 45450 73506 45484
rect 72620 45390 72660 45432
rect 73690 45432 73702 45590
rect 73702 45432 73730 45590
rect 73690 45390 73730 45432
rect 77610 45900 77650 45950
rect 77610 45742 77636 45900
rect 77636 45742 77650 45900
rect 78680 45900 78720 45950
rect 77822 45848 77998 45882
rect 78320 45848 78496 45882
rect 77738 45804 77772 45838
rect 78555 45804 78589 45838
rect 77822 45760 77998 45794
rect 78320 45760 78496 45794
rect 77610 45690 77650 45742
rect 77610 45590 77650 45630
rect 77610 45432 77636 45590
rect 77636 45432 77650 45590
rect 78680 45742 78692 45900
rect 78692 45742 78720 45900
rect 78680 45710 78720 45742
rect 78680 45590 78720 45630
rect 77822 45538 77998 45572
rect 78320 45538 78496 45572
rect 77738 45494 77772 45528
rect 78555 45494 78589 45528
rect 77822 45450 77998 45484
rect 78320 45450 78496 45484
rect 77610 45390 77650 45432
rect 78680 45432 78692 45590
rect 78692 45432 78720 45590
rect 78680 45390 78720 45432
rect 2760 44190 2800 44240
rect 2760 44032 2786 44190
rect 2786 44032 2800 44190
rect 3830 44190 3870 44240
rect 2972 44138 3148 44172
rect 3470 44138 3646 44172
rect 2888 44094 2922 44128
rect 3705 44094 3739 44128
rect 2972 44050 3148 44084
rect 3470 44050 3646 44084
rect 2760 43980 2800 44032
rect 2760 43880 2800 43920
rect 2760 43722 2786 43880
rect 2786 43722 2800 43880
rect 3830 44032 3842 44190
rect 3842 44032 3870 44190
rect 3830 44000 3870 44032
rect 3830 43880 3870 43920
rect 2972 43828 3148 43862
rect 3470 43828 3646 43862
rect 2888 43784 2922 43818
rect 3705 43784 3739 43818
rect 2972 43740 3148 43774
rect 3470 43740 3646 43774
rect 2760 43680 2800 43722
rect 3830 43722 3842 43880
rect 3842 43722 3870 43880
rect 3830 43680 3870 43722
rect 7750 44190 7790 44240
rect 7750 44032 7776 44190
rect 7776 44032 7790 44190
rect 8820 44190 8860 44240
rect 7962 44138 8138 44172
rect 8460 44138 8636 44172
rect 7878 44094 7912 44128
rect 8695 44094 8729 44128
rect 7962 44050 8138 44084
rect 8460 44050 8636 44084
rect 7750 43980 7790 44032
rect 7750 43880 7790 43920
rect 7750 43722 7776 43880
rect 7776 43722 7790 43880
rect 8820 44032 8832 44190
rect 8832 44032 8860 44190
rect 8820 44000 8860 44032
rect 8820 43880 8860 43920
rect 7962 43828 8138 43862
rect 8460 43828 8636 43862
rect 7878 43784 7912 43818
rect 8695 43784 8729 43818
rect 7962 43740 8138 43774
rect 8460 43740 8636 43774
rect 7750 43680 7790 43722
rect 8820 43722 8832 43880
rect 8832 43722 8860 43880
rect 8820 43680 8860 43722
rect 12740 44190 12780 44240
rect 12740 44032 12766 44190
rect 12766 44032 12780 44190
rect 13810 44190 13850 44240
rect 12952 44138 13128 44172
rect 13450 44138 13626 44172
rect 12868 44094 12902 44128
rect 13685 44094 13719 44128
rect 12952 44050 13128 44084
rect 13450 44050 13626 44084
rect 12740 43980 12780 44032
rect 12740 43880 12780 43920
rect 12740 43722 12766 43880
rect 12766 43722 12780 43880
rect 13810 44032 13822 44190
rect 13822 44032 13850 44190
rect 13810 44000 13850 44032
rect 13810 43880 13850 43920
rect 12952 43828 13128 43862
rect 13450 43828 13626 43862
rect 12868 43784 12902 43818
rect 13685 43784 13719 43818
rect 12952 43740 13128 43774
rect 13450 43740 13626 43774
rect 12740 43680 12780 43722
rect 13810 43722 13822 43880
rect 13822 43722 13850 43880
rect 13810 43680 13850 43722
rect 17730 44190 17770 44240
rect 17730 44032 17756 44190
rect 17756 44032 17770 44190
rect 18800 44190 18840 44240
rect 17942 44138 18118 44172
rect 18440 44138 18616 44172
rect 17858 44094 17892 44128
rect 18675 44094 18709 44128
rect 17942 44050 18118 44084
rect 18440 44050 18616 44084
rect 17730 43980 17770 44032
rect 17730 43880 17770 43920
rect 17730 43722 17756 43880
rect 17756 43722 17770 43880
rect 18800 44032 18812 44190
rect 18812 44032 18840 44190
rect 18800 44000 18840 44032
rect 18800 43880 18840 43920
rect 17942 43828 18118 43862
rect 18440 43828 18616 43862
rect 17858 43784 17892 43818
rect 18675 43784 18709 43818
rect 17942 43740 18118 43774
rect 18440 43740 18616 43774
rect 17730 43680 17770 43722
rect 18800 43722 18812 43880
rect 18812 43722 18840 43880
rect 18800 43680 18840 43722
rect 22720 44190 22760 44240
rect 22720 44032 22746 44190
rect 22746 44032 22760 44190
rect 23790 44190 23830 44240
rect 22932 44138 23108 44172
rect 23430 44138 23606 44172
rect 22848 44094 22882 44128
rect 23665 44094 23699 44128
rect 22932 44050 23108 44084
rect 23430 44050 23606 44084
rect 22720 43980 22760 44032
rect 22720 43880 22760 43920
rect 22720 43722 22746 43880
rect 22746 43722 22760 43880
rect 23790 44032 23802 44190
rect 23802 44032 23830 44190
rect 23790 44000 23830 44032
rect 23790 43880 23830 43920
rect 22932 43828 23108 43862
rect 23430 43828 23606 43862
rect 22848 43784 22882 43818
rect 23665 43784 23699 43818
rect 22932 43740 23108 43774
rect 23430 43740 23606 43774
rect 22720 43680 22760 43722
rect 23790 43722 23802 43880
rect 23802 43722 23830 43880
rect 23790 43680 23830 43722
rect 27710 44190 27750 44240
rect 27710 44032 27736 44190
rect 27736 44032 27750 44190
rect 28780 44190 28820 44240
rect 27922 44138 28098 44172
rect 28420 44138 28596 44172
rect 27838 44094 27872 44128
rect 28655 44094 28689 44128
rect 27922 44050 28098 44084
rect 28420 44050 28596 44084
rect 27710 43980 27750 44032
rect 27710 43880 27750 43920
rect 27710 43722 27736 43880
rect 27736 43722 27750 43880
rect 28780 44032 28792 44190
rect 28792 44032 28820 44190
rect 28780 44000 28820 44032
rect 28780 43880 28820 43920
rect 27922 43828 28098 43862
rect 28420 43828 28596 43862
rect 27838 43784 27872 43818
rect 28655 43784 28689 43818
rect 27922 43740 28098 43774
rect 28420 43740 28596 43774
rect 27710 43680 27750 43722
rect 28780 43722 28792 43880
rect 28792 43722 28820 43880
rect 28780 43680 28820 43722
rect 32700 44190 32740 44240
rect 32700 44032 32726 44190
rect 32726 44032 32740 44190
rect 33770 44190 33810 44240
rect 32912 44138 33088 44172
rect 33410 44138 33586 44172
rect 32828 44094 32862 44128
rect 33645 44094 33679 44128
rect 32912 44050 33088 44084
rect 33410 44050 33586 44084
rect 32700 43980 32740 44032
rect 32700 43880 32740 43920
rect 32700 43722 32726 43880
rect 32726 43722 32740 43880
rect 33770 44032 33782 44190
rect 33782 44032 33810 44190
rect 33770 44000 33810 44032
rect 33770 43880 33810 43920
rect 32912 43828 33088 43862
rect 33410 43828 33586 43862
rect 32828 43784 32862 43818
rect 33645 43784 33679 43818
rect 32912 43740 33088 43774
rect 33410 43740 33586 43774
rect 32700 43680 32740 43722
rect 33770 43722 33782 43880
rect 33782 43722 33810 43880
rect 33770 43680 33810 43722
rect 37690 44190 37730 44240
rect 37690 44032 37716 44190
rect 37716 44032 37730 44190
rect 38760 44190 38800 44240
rect 37902 44138 38078 44172
rect 38400 44138 38576 44172
rect 37818 44094 37852 44128
rect 38635 44094 38669 44128
rect 37902 44050 38078 44084
rect 38400 44050 38576 44084
rect 37690 43980 37730 44032
rect 37690 43880 37730 43920
rect 37690 43722 37716 43880
rect 37716 43722 37730 43880
rect 38760 44032 38772 44190
rect 38772 44032 38800 44190
rect 38760 44000 38800 44032
rect 38760 43880 38800 43920
rect 37902 43828 38078 43862
rect 38400 43828 38576 43862
rect 37818 43784 37852 43818
rect 38635 43784 38669 43818
rect 37902 43740 38078 43774
rect 38400 43740 38576 43774
rect 37690 43680 37730 43722
rect 38760 43722 38772 43880
rect 38772 43722 38800 43880
rect 38760 43680 38800 43722
rect 42680 44190 42720 44240
rect 42680 44032 42706 44190
rect 42706 44032 42720 44190
rect 43750 44190 43790 44240
rect 42892 44138 43068 44172
rect 43390 44138 43566 44172
rect 42808 44094 42842 44128
rect 43625 44094 43659 44128
rect 42892 44050 43068 44084
rect 43390 44050 43566 44084
rect 42680 43980 42720 44032
rect 42680 43880 42720 43920
rect 42680 43722 42706 43880
rect 42706 43722 42720 43880
rect 43750 44032 43762 44190
rect 43762 44032 43790 44190
rect 43750 44000 43790 44032
rect 43750 43880 43790 43920
rect 42892 43828 43068 43862
rect 43390 43828 43566 43862
rect 42808 43784 42842 43818
rect 43625 43784 43659 43818
rect 42892 43740 43068 43774
rect 43390 43740 43566 43774
rect 42680 43680 42720 43722
rect 43750 43722 43762 43880
rect 43762 43722 43790 43880
rect 43750 43680 43790 43722
rect 47670 44190 47710 44240
rect 47670 44032 47696 44190
rect 47696 44032 47710 44190
rect 48740 44190 48780 44240
rect 47882 44138 48058 44172
rect 48380 44138 48556 44172
rect 47798 44094 47832 44128
rect 48615 44094 48649 44128
rect 47882 44050 48058 44084
rect 48380 44050 48556 44084
rect 47670 43980 47710 44032
rect 47670 43880 47710 43920
rect 47670 43722 47696 43880
rect 47696 43722 47710 43880
rect 48740 44032 48752 44190
rect 48752 44032 48780 44190
rect 48740 44000 48780 44032
rect 48740 43880 48780 43920
rect 47882 43828 48058 43862
rect 48380 43828 48556 43862
rect 47798 43784 47832 43818
rect 48615 43784 48649 43818
rect 47882 43740 48058 43774
rect 48380 43740 48556 43774
rect 47670 43680 47710 43722
rect 48740 43722 48752 43880
rect 48752 43722 48780 43880
rect 48740 43680 48780 43722
rect 52660 44190 52700 44240
rect 52660 44032 52686 44190
rect 52686 44032 52700 44190
rect 53730 44190 53770 44240
rect 52872 44138 53048 44172
rect 53370 44138 53546 44172
rect 52788 44094 52822 44128
rect 53605 44094 53639 44128
rect 52872 44050 53048 44084
rect 53370 44050 53546 44084
rect 52660 43980 52700 44032
rect 52660 43880 52700 43920
rect 52660 43722 52686 43880
rect 52686 43722 52700 43880
rect 53730 44032 53742 44190
rect 53742 44032 53770 44190
rect 53730 44000 53770 44032
rect 53730 43880 53770 43920
rect 52872 43828 53048 43862
rect 53370 43828 53546 43862
rect 52788 43784 52822 43818
rect 53605 43784 53639 43818
rect 52872 43740 53048 43774
rect 53370 43740 53546 43774
rect 52660 43680 52700 43722
rect 53730 43722 53742 43880
rect 53742 43722 53770 43880
rect 53730 43680 53770 43722
rect 57650 44190 57690 44240
rect 57650 44032 57676 44190
rect 57676 44032 57690 44190
rect 58720 44190 58760 44240
rect 57862 44138 58038 44172
rect 58360 44138 58536 44172
rect 57778 44094 57812 44128
rect 58595 44094 58629 44128
rect 57862 44050 58038 44084
rect 58360 44050 58536 44084
rect 57650 43980 57690 44032
rect 57650 43880 57690 43920
rect 57650 43722 57676 43880
rect 57676 43722 57690 43880
rect 58720 44032 58732 44190
rect 58732 44032 58760 44190
rect 58720 44000 58760 44032
rect 58720 43880 58760 43920
rect 57862 43828 58038 43862
rect 58360 43828 58536 43862
rect 57778 43784 57812 43818
rect 58595 43784 58629 43818
rect 57862 43740 58038 43774
rect 58360 43740 58536 43774
rect 57650 43680 57690 43722
rect 58720 43722 58732 43880
rect 58732 43722 58760 43880
rect 58720 43680 58760 43722
rect 62640 44190 62680 44240
rect 62640 44032 62666 44190
rect 62666 44032 62680 44190
rect 63710 44190 63750 44240
rect 62852 44138 63028 44172
rect 63350 44138 63526 44172
rect 62768 44094 62802 44128
rect 63585 44094 63619 44128
rect 62852 44050 63028 44084
rect 63350 44050 63526 44084
rect 62640 43980 62680 44032
rect 62640 43880 62680 43920
rect 62640 43722 62666 43880
rect 62666 43722 62680 43880
rect 63710 44032 63722 44190
rect 63722 44032 63750 44190
rect 63710 44000 63750 44032
rect 63710 43880 63750 43920
rect 62852 43828 63028 43862
rect 63350 43828 63526 43862
rect 62768 43784 62802 43818
rect 63585 43784 63619 43818
rect 62852 43740 63028 43774
rect 63350 43740 63526 43774
rect 62640 43680 62680 43722
rect 63710 43722 63722 43880
rect 63722 43722 63750 43880
rect 63710 43680 63750 43722
rect 67630 44190 67670 44240
rect 67630 44032 67656 44190
rect 67656 44032 67670 44190
rect 68700 44190 68740 44240
rect 67842 44138 68018 44172
rect 68340 44138 68516 44172
rect 67758 44094 67792 44128
rect 68575 44094 68609 44128
rect 67842 44050 68018 44084
rect 68340 44050 68516 44084
rect 67630 43980 67670 44032
rect 67630 43880 67670 43920
rect 67630 43722 67656 43880
rect 67656 43722 67670 43880
rect 68700 44032 68712 44190
rect 68712 44032 68740 44190
rect 68700 44000 68740 44032
rect 68700 43880 68740 43920
rect 67842 43828 68018 43862
rect 68340 43828 68516 43862
rect 67758 43784 67792 43818
rect 68575 43784 68609 43818
rect 67842 43740 68018 43774
rect 68340 43740 68516 43774
rect 67630 43680 67670 43722
rect 68700 43722 68712 43880
rect 68712 43722 68740 43880
rect 68700 43680 68740 43722
rect 72620 44190 72660 44240
rect 72620 44032 72646 44190
rect 72646 44032 72660 44190
rect 73690 44190 73730 44240
rect 72832 44138 73008 44172
rect 73330 44138 73506 44172
rect 72748 44094 72782 44128
rect 73565 44094 73599 44128
rect 72832 44050 73008 44084
rect 73330 44050 73506 44084
rect 72620 43980 72660 44032
rect 72620 43880 72660 43920
rect 72620 43722 72646 43880
rect 72646 43722 72660 43880
rect 73690 44032 73702 44190
rect 73702 44032 73730 44190
rect 73690 44000 73730 44032
rect 73690 43880 73730 43920
rect 72832 43828 73008 43862
rect 73330 43828 73506 43862
rect 72748 43784 72782 43818
rect 73565 43784 73599 43818
rect 72832 43740 73008 43774
rect 73330 43740 73506 43774
rect 72620 43680 72660 43722
rect 73690 43722 73702 43880
rect 73702 43722 73730 43880
rect 73690 43680 73730 43722
rect 77610 44190 77650 44240
rect 77610 44032 77636 44190
rect 77636 44032 77650 44190
rect 78680 44190 78720 44240
rect 77822 44138 77998 44172
rect 78320 44138 78496 44172
rect 77738 44094 77772 44128
rect 78555 44094 78589 44128
rect 77822 44050 77998 44084
rect 78320 44050 78496 44084
rect 77610 43980 77650 44032
rect 77610 43880 77650 43920
rect 77610 43722 77636 43880
rect 77636 43722 77650 43880
rect 78680 44032 78692 44190
rect 78692 44032 78720 44190
rect 78680 44000 78720 44032
rect 78680 43880 78720 43920
rect 77822 43828 77998 43862
rect 78320 43828 78496 43862
rect 77738 43784 77772 43818
rect 78555 43784 78589 43818
rect 77822 43740 77998 43774
rect 78320 43740 78496 43774
rect 77610 43680 77650 43722
rect 78680 43722 78692 43880
rect 78692 43722 78720 43880
rect 78680 43680 78720 43722
rect 2760 42480 2800 42530
rect 2760 42322 2786 42480
rect 2786 42322 2800 42480
rect 3830 42480 3870 42530
rect 2972 42428 3148 42462
rect 3470 42428 3646 42462
rect 2888 42384 2922 42418
rect 3705 42384 3739 42418
rect 2972 42340 3148 42374
rect 3470 42340 3646 42374
rect 2760 42270 2800 42322
rect 2760 42170 2800 42210
rect 2760 42012 2786 42170
rect 2786 42012 2800 42170
rect 3830 42322 3842 42480
rect 3842 42322 3870 42480
rect 3830 42290 3870 42322
rect 3830 42170 3870 42210
rect 2972 42118 3148 42152
rect 3470 42118 3646 42152
rect 2888 42074 2922 42108
rect 3705 42074 3739 42108
rect 2972 42030 3148 42064
rect 3470 42030 3646 42064
rect 2760 41970 2800 42012
rect 3830 42012 3842 42170
rect 3842 42012 3870 42170
rect 3830 41970 3870 42012
rect 7750 42480 7790 42530
rect 7750 42322 7776 42480
rect 7776 42322 7790 42480
rect 8820 42480 8860 42530
rect 7962 42428 8138 42462
rect 8460 42428 8636 42462
rect 7878 42384 7912 42418
rect 8695 42384 8729 42418
rect 7962 42340 8138 42374
rect 8460 42340 8636 42374
rect 7750 42270 7790 42322
rect 7750 42170 7790 42210
rect 7750 42012 7776 42170
rect 7776 42012 7790 42170
rect 8820 42322 8832 42480
rect 8832 42322 8860 42480
rect 8820 42290 8860 42322
rect 8820 42170 8860 42210
rect 7962 42118 8138 42152
rect 8460 42118 8636 42152
rect 7878 42074 7912 42108
rect 8695 42074 8729 42108
rect 7962 42030 8138 42064
rect 8460 42030 8636 42064
rect 7750 41970 7790 42012
rect 8820 42012 8832 42170
rect 8832 42012 8860 42170
rect 8820 41970 8860 42012
rect 12740 42480 12780 42530
rect 12740 42322 12766 42480
rect 12766 42322 12780 42480
rect 13810 42480 13850 42530
rect 12952 42428 13128 42462
rect 13450 42428 13626 42462
rect 12868 42384 12902 42418
rect 13685 42384 13719 42418
rect 12952 42340 13128 42374
rect 13450 42340 13626 42374
rect 12740 42270 12780 42322
rect 12740 42170 12780 42210
rect 12740 42012 12766 42170
rect 12766 42012 12780 42170
rect 13810 42322 13822 42480
rect 13822 42322 13850 42480
rect 13810 42290 13850 42322
rect 13810 42170 13850 42210
rect 12952 42118 13128 42152
rect 13450 42118 13626 42152
rect 12868 42074 12902 42108
rect 13685 42074 13719 42108
rect 12952 42030 13128 42064
rect 13450 42030 13626 42064
rect 12740 41970 12780 42012
rect 13810 42012 13822 42170
rect 13822 42012 13850 42170
rect 13810 41970 13850 42012
rect 17730 42480 17770 42530
rect 17730 42322 17756 42480
rect 17756 42322 17770 42480
rect 18800 42480 18840 42530
rect 17942 42428 18118 42462
rect 18440 42428 18616 42462
rect 17858 42384 17892 42418
rect 18675 42384 18709 42418
rect 17942 42340 18118 42374
rect 18440 42340 18616 42374
rect 17730 42270 17770 42322
rect 17730 42170 17770 42210
rect 17730 42012 17756 42170
rect 17756 42012 17770 42170
rect 18800 42322 18812 42480
rect 18812 42322 18840 42480
rect 18800 42290 18840 42322
rect 18800 42170 18840 42210
rect 17942 42118 18118 42152
rect 18440 42118 18616 42152
rect 17858 42074 17892 42108
rect 18675 42074 18709 42108
rect 17942 42030 18118 42064
rect 18440 42030 18616 42064
rect 17730 41970 17770 42012
rect 18800 42012 18812 42170
rect 18812 42012 18840 42170
rect 18800 41970 18840 42012
rect 22720 42480 22760 42530
rect 22720 42322 22746 42480
rect 22746 42322 22760 42480
rect 23790 42480 23830 42530
rect 22932 42428 23108 42462
rect 23430 42428 23606 42462
rect 22848 42384 22882 42418
rect 23665 42384 23699 42418
rect 22932 42340 23108 42374
rect 23430 42340 23606 42374
rect 22720 42270 22760 42322
rect 22720 42170 22760 42210
rect 22720 42012 22746 42170
rect 22746 42012 22760 42170
rect 23790 42322 23802 42480
rect 23802 42322 23830 42480
rect 23790 42290 23830 42322
rect 23790 42170 23830 42210
rect 22932 42118 23108 42152
rect 23430 42118 23606 42152
rect 22848 42074 22882 42108
rect 23665 42074 23699 42108
rect 22932 42030 23108 42064
rect 23430 42030 23606 42064
rect 22720 41970 22760 42012
rect 23790 42012 23802 42170
rect 23802 42012 23830 42170
rect 23790 41970 23830 42012
rect 27710 42480 27750 42530
rect 27710 42322 27736 42480
rect 27736 42322 27750 42480
rect 28780 42480 28820 42530
rect 27922 42428 28098 42462
rect 28420 42428 28596 42462
rect 27838 42384 27872 42418
rect 28655 42384 28689 42418
rect 27922 42340 28098 42374
rect 28420 42340 28596 42374
rect 27710 42270 27750 42322
rect 27710 42170 27750 42210
rect 27710 42012 27736 42170
rect 27736 42012 27750 42170
rect 28780 42322 28792 42480
rect 28792 42322 28820 42480
rect 28780 42290 28820 42322
rect 28780 42170 28820 42210
rect 27922 42118 28098 42152
rect 28420 42118 28596 42152
rect 27838 42074 27872 42108
rect 28655 42074 28689 42108
rect 27922 42030 28098 42064
rect 28420 42030 28596 42064
rect 27710 41970 27750 42012
rect 28780 42012 28792 42170
rect 28792 42012 28820 42170
rect 28780 41970 28820 42012
rect 32700 42480 32740 42530
rect 32700 42322 32726 42480
rect 32726 42322 32740 42480
rect 33770 42480 33810 42530
rect 32912 42428 33088 42462
rect 33410 42428 33586 42462
rect 32828 42384 32862 42418
rect 33645 42384 33679 42418
rect 32912 42340 33088 42374
rect 33410 42340 33586 42374
rect 32700 42270 32740 42322
rect 32700 42170 32740 42210
rect 32700 42012 32726 42170
rect 32726 42012 32740 42170
rect 33770 42322 33782 42480
rect 33782 42322 33810 42480
rect 33770 42290 33810 42322
rect 33770 42170 33810 42210
rect 32912 42118 33088 42152
rect 33410 42118 33586 42152
rect 32828 42074 32862 42108
rect 33645 42074 33679 42108
rect 32912 42030 33088 42064
rect 33410 42030 33586 42064
rect 32700 41970 32740 42012
rect 33770 42012 33782 42170
rect 33782 42012 33810 42170
rect 33770 41970 33810 42012
rect 37690 42480 37730 42530
rect 37690 42322 37716 42480
rect 37716 42322 37730 42480
rect 38760 42480 38800 42530
rect 37902 42428 38078 42462
rect 38400 42428 38576 42462
rect 37818 42384 37852 42418
rect 38635 42384 38669 42418
rect 37902 42340 38078 42374
rect 38400 42340 38576 42374
rect 37690 42270 37730 42322
rect 37690 42170 37730 42210
rect 37690 42012 37716 42170
rect 37716 42012 37730 42170
rect 38760 42322 38772 42480
rect 38772 42322 38800 42480
rect 38760 42290 38800 42322
rect 38760 42170 38800 42210
rect 37902 42118 38078 42152
rect 38400 42118 38576 42152
rect 37818 42074 37852 42108
rect 38635 42074 38669 42108
rect 37902 42030 38078 42064
rect 38400 42030 38576 42064
rect 37690 41970 37730 42012
rect 38760 42012 38772 42170
rect 38772 42012 38800 42170
rect 38760 41970 38800 42012
rect 42680 42480 42720 42530
rect 42680 42322 42706 42480
rect 42706 42322 42720 42480
rect 43750 42480 43790 42530
rect 42892 42428 43068 42462
rect 43390 42428 43566 42462
rect 42808 42384 42842 42418
rect 43625 42384 43659 42418
rect 42892 42340 43068 42374
rect 43390 42340 43566 42374
rect 42680 42270 42720 42322
rect 42680 42170 42720 42210
rect 42680 42012 42706 42170
rect 42706 42012 42720 42170
rect 43750 42322 43762 42480
rect 43762 42322 43790 42480
rect 43750 42290 43790 42322
rect 43750 42170 43790 42210
rect 42892 42118 43068 42152
rect 43390 42118 43566 42152
rect 42808 42074 42842 42108
rect 43625 42074 43659 42108
rect 42892 42030 43068 42064
rect 43390 42030 43566 42064
rect 42680 41970 42720 42012
rect 43750 42012 43762 42170
rect 43762 42012 43790 42170
rect 43750 41970 43790 42012
rect 47670 42480 47710 42530
rect 47670 42322 47696 42480
rect 47696 42322 47710 42480
rect 48740 42480 48780 42530
rect 47882 42428 48058 42462
rect 48380 42428 48556 42462
rect 47798 42384 47832 42418
rect 48615 42384 48649 42418
rect 47882 42340 48058 42374
rect 48380 42340 48556 42374
rect 47670 42270 47710 42322
rect 47670 42170 47710 42210
rect 47670 42012 47696 42170
rect 47696 42012 47710 42170
rect 48740 42322 48752 42480
rect 48752 42322 48780 42480
rect 48740 42290 48780 42322
rect 48740 42170 48780 42210
rect 47882 42118 48058 42152
rect 48380 42118 48556 42152
rect 47798 42074 47832 42108
rect 48615 42074 48649 42108
rect 47882 42030 48058 42064
rect 48380 42030 48556 42064
rect 47670 41970 47710 42012
rect 48740 42012 48752 42170
rect 48752 42012 48780 42170
rect 48740 41970 48780 42012
rect 52660 42480 52700 42530
rect 52660 42322 52686 42480
rect 52686 42322 52700 42480
rect 53730 42480 53770 42530
rect 52872 42428 53048 42462
rect 53370 42428 53546 42462
rect 52788 42384 52822 42418
rect 53605 42384 53639 42418
rect 52872 42340 53048 42374
rect 53370 42340 53546 42374
rect 52660 42270 52700 42322
rect 52660 42170 52700 42210
rect 52660 42012 52686 42170
rect 52686 42012 52700 42170
rect 53730 42322 53742 42480
rect 53742 42322 53770 42480
rect 53730 42290 53770 42322
rect 53730 42170 53770 42210
rect 52872 42118 53048 42152
rect 53370 42118 53546 42152
rect 52788 42074 52822 42108
rect 53605 42074 53639 42108
rect 52872 42030 53048 42064
rect 53370 42030 53546 42064
rect 52660 41970 52700 42012
rect 53730 42012 53742 42170
rect 53742 42012 53770 42170
rect 53730 41970 53770 42012
rect 57650 42480 57690 42530
rect 57650 42322 57676 42480
rect 57676 42322 57690 42480
rect 58720 42480 58760 42530
rect 57862 42428 58038 42462
rect 58360 42428 58536 42462
rect 57778 42384 57812 42418
rect 58595 42384 58629 42418
rect 57862 42340 58038 42374
rect 58360 42340 58536 42374
rect 57650 42270 57690 42322
rect 57650 42170 57690 42210
rect 57650 42012 57676 42170
rect 57676 42012 57690 42170
rect 58720 42322 58732 42480
rect 58732 42322 58760 42480
rect 58720 42290 58760 42322
rect 58720 42170 58760 42210
rect 57862 42118 58038 42152
rect 58360 42118 58536 42152
rect 57778 42074 57812 42108
rect 58595 42074 58629 42108
rect 57862 42030 58038 42064
rect 58360 42030 58536 42064
rect 57650 41970 57690 42012
rect 58720 42012 58732 42170
rect 58732 42012 58760 42170
rect 58720 41970 58760 42012
rect 62640 42480 62680 42530
rect 62640 42322 62666 42480
rect 62666 42322 62680 42480
rect 63710 42480 63750 42530
rect 62852 42428 63028 42462
rect 63350 42428 63526 42462
rect 62768 42384 62802 42418
rect 63585 42384 63619 42418
rect 62852 42340 63028 42374
rect 63350 42340 63526 42374
rect 62640 42270 62680 42322
rect 62640 42170 62680 42210
rect 62640 42012 62666 42170
rect 62666 42012 62680 42170
rect 63710 42322 63722 42480
rect 63722 42322 63750 42480
rect 63710 42290 63750 42322
rect 63710 42170 63750 42210
rect 62852 42118 63028 42152
rect 63350 42118 63526 42152
rect 62768 42074 62802 42108
rect 63585 42074 63619 42108
rect 62852 42030 63028 42064
rect 63350 42030 63526 42064
rect 62640 41970 62680 42012
rect 63710 42012 63722 42170
rect 63722 42012 63750 42170
rect 63710 41970 63750 42012
rect 67630 42480 67670 42530
rect 67630 42322 67656 42480
rect 67656 42322 67670 42480
rect 68700 42480 68740 42530
rect 67842 42428 68018 42462
rect 68340 42428 68516 42462
rect 67758 42384 67792 42418
rect 68575 42384 68609 42418
rect 67842 42340 68018 42374
rect 68340 42340 68516 42374
rect 67630 42270 67670 42322
rect 67630 42170 67670 42210
rect 67630 42012 67656 42170
rect 67656 42012 67670 42170
rect 68700 42322 68712 42480
rect 68712 42322 68740 42480
rect 68700 42290 68740 42322
rect 68700 42170 68740 42210
rect 67842 42118 68018 42152
rect 68340 42118 68516 42152
rect 67758 42074 67792 42108
rect 68575 42074 68609 42108
rect 67842 42030 68018 42064
rect 68340 42030 68516 42064
rect 67630 41970 67670 42012
rect 68700 42012 68712 42170
rect 68712 42012 68740 42170
rect 68700 41970 68740 42012
rect 72620 42480 72660 42530
rect 72620 42322 72646 42480
rect 72646 42322 72660 42480
rect 73690 42480 73730 42530
rect 72832 42428 73008 42462
rect 73330 42428 73506 42462
rect 72748 42384 72782 42418
rect 73565 42384 73599 42418
rect 72832 42340 73008 42374
rect 73330 42340 73506 42374
rect 72620 42270 72660 42322
rect 72620 42170 72660 42210
rect 72620 42012 72646 42170
rect 72646 42012 72660 42170
rect 73690 42322 73702 42480
rect 73702 42322 73730 42480
rect 73690 42290 73730 42322
rect 73690 42170 73730 42210
rect 72832 42118 73008 42152
rect 73330 42118 73506 42152
rect 72748 42074 72782 42108
rect 73565 42074 73599 42108
rect 72832 42030 73008 42064
rect 73330 42030 73506 42064
rect 72620 41970 72660 42012
rect 73690 42012 73702 42170
rect 73702 42012 73730 42170
rect 73690 41970 73730 42012
rect 77610 42480 77650 42530
rect 77610 42322 77636 42480
rect 77636 42322 77650 42480
rect 78680 42480 78720 42530
rect 77822 42428 77998 42462
rect 78320 42428 78496 42462
rect 77738 42384 77772 42418
rect 78555 42384 78589 42418
rect 77822 42340 77998 42374
rect 78320 42340 78496 42374
rect 77610 42270 77650 42322
rect 77610 42170 77650 42210
rect 77610 42012 77636 42170
rect 77636 42012 77650 42170
rect 78680 42322 78692 42480
rect 78692 42322 78720 42480
rect 78680 42290 78720 42322
rect 78680 42170 78720 42210
rect 77822 42118 77998 42152
rect 78320 42118 78496 42152
rect 77738 42074 77772 42108
rect 78555 42074 78589 42108
rect 77822 42030 77998 42064
rect 78320 42030 78496 42064
rect 77610 41970 77650 42012
rect 78680 42012 78692 42170
rect 78692 42012 78720 42170
rect 78680 41970 78720 42012
rect 2760 40770 2800 40820
rect 2760 40612 2786 40770
rect 2786 40612 2800 40770
rect 3830 40770 3870 40820
rect 2972 40718 3148 40752
rect 3470 40718 3646 40752
rect 2888 40674 2922 40708
rect 3705 40674 3739 40708
rect 2972 40630 3148 40664
rect 3470 40630 3646 40664
rect 2760 40560 2800 40612
rect 2760 40460 2800 40500
rect 2760 40302 2786 40460
rect 2786 40302 2800 40460
rect 3830 40612 3842 40770
rect 3842 40612 3870 40770
rect 3830 40580 3870 40612
rect 3830 40460 3870 40500
rect 2972 40408 3148 40442
rect 3470 40408 3646 40442
rect 2888 40364 2922 40398
rect 3705 40364 3739 40398
rect 2972 40320 3148 40354
rect 3470 40320 3646 40354
rect 2760 40260 2800 40302
rect 3830 40302 3842 40460
rect 3842 40302 3870 40460
rect 3830 40260 3870 40302
rect 7750 40770 7790 40820
rect 7750 40612 7776 40770
rect 7776 40612 7790 40770
rect 8820 40770 8860 40820
rect 7962 40718 8138 40752
rect 8460 40718 8636 40752
rect 7878 40674 7912 40708
rect 8695 40674 8729 40708
rect 7962 40630 8138 40664
rect 8460 40630 8636 40664
rect 7750 40560 7790 40612
rect 7750 40460 7790 40500
rect 7750 40302 7776 40460
rect 7776 40302 7790 40460
rect 8820 40612 8832 40770
rect 8832 40612 8860 40770
rect 8820 40580 8860 40612
rect 8820 40460 8860 40500
rect 7962 40408 8138 40442
rect 8460 40408 8636 40442
rect 7878 40364 7912 40398
rect 8695 40364 8729 40398
rect 7962 40320 8138 40354
rect 8460 40320 8636 40354
rect 7750 40260 7790 40302
rect 8820 40302 8832 40460
rect 8832 40302 8860 40460
rect 8820 40260 8860 40302
rect 12740 40770 12780 40820
rect 12740 40612 12766 40770
rect 12766 40612 12780 40770
rect 13810 40770 13850 40820
rect 12952 40718 13128 40752
rect 13450 40718 13626 40752
rect 12868 40674 12902 40708
rect 13685 40674 13719 40708
rect 12952 40630 13128 40664
rect 13450 40630 13626 40664
rect 12740 40560 12780 40612
rect 12740 40460 12780 40500
rect 12740 40302 12766 40460
rect 12766 40302 12780 40460
rect 13810 40612 13822 40770
rect 13822 40612 13850 40770
rect 13810 40580 13850 40612
rect 13810 40460 13850 40500
rect 12952 40408 13128 40442
rect 13450 40408 13626 40442
rect 12868 40364 12902 40398
rect 13685 40364 13719 40398
rect 12952 40320 13128 40354
rect 13450 40320 13626 40354
rect 12740 40260 12780 40302
rect 13810 40302 13822 40460
rect 13822 40302 13850 40460
rect 13810 40260 13850 40302
rect 17730 40770 17770 40820
rect 17730 40612 17756 40770
rect 17756 40612 17770 40770
rect 18800 40770 18840 40820
rect 17942 40718 18118 40752
rect 18440 40718 18616 40752
rect 17858 40674 17892 40708
rect 18675 40674 18709 40708
rect 17942 40630 18118 40664
rect 18440 40630 18616 40664
rect 17730 40560 17770 40612
rect 17730 40460 17770 40500
rect 17730 40302 17756 40460
rect 17756 40302 17770 40460
rect 18800 40612 18812 40770
rect 18812 40612 18840 40770
rect 18800 40580 18840 40612
rect 18800 40460 18840 40500
rect 17942 40408 18118 40442
rect 18440 40408 18616 40442
rect 17858 40364 17892 40398
rect 18675 40364 18709 40398
rect 17942 40320 18118 40354
rect 18440 40320 18616 40354
rect 17730 40260 17770 40302
rect 18800 40302 18812 40460
rect 18812 40302 18840 40460
rect 18800 40260 18840 40302
rect 22720 40770 22760 40820
rect 22720 40612 22746 40770
rect 22746 40612 22760 40770
rect 23790 40770 23830 40820
rect 22932 40718 23108 40752
rect 23430 40718 23606 40752
rect 22848 40674 22882 40708
rect 23665 40674 23699 40708
rect 22932 40630 23108 40664
rect 23430 40630 23606 40664
rect 22720 40560 22760 40612
rect 22720 40460 22760 40500
rect 22720 40302 22746 40460
rect 22746 40302 22760 40460
rect 23790 40612 23802 40770
rect 23802 40612 23830 40770
rect 23790 40580 23830 40612
rect 23790 40460 23830 40500
rect 22932 40408 23108 40442
rect 23430 40408 23606 40442
rect 22848 40364 22882 40398
rect 23665 40364 23699 40398
rect 22932 40320 23108 40354
rect 23430 40320 23606 40354
rect 22720 40260 22760 40302
rect 23790 40302 23802 40460
rect 23802 40302 23830 40460
rect 23790 40260 23830 40302
rect 27710 40770 27750 40820
rect 27710 40612 27736 40770
rect 27736 40612 27750 40770
rect 28780 40770 28820 40820
rect 27922 40718 28098 40752
rect 28420 40718 28596 40752
rect 27838 40674 27872 40708
rect 28655 40674 28689 40708
rect 27922 40630 28098 40664
rect 28420 40630 28596 40664
rect 27710 40560 27750 40612
rect 27710 40460 27750 40500
rect 27710 40302 27736 40460
rect 27736 40302 27750 40460
rect 28780 40612 28792 40770
rect 28792 40612 28820 40770
rect 28780 40580 28820 40612
rect 28780 40460 28820 40500
rect 27922 40408 28098 40442
rect 28420 40408 28596 40442
rect 27838 40364 27872 40398
rect 28655 40364 28689 40398
rect 27922 40320 28098 40354
rect 28420 40320 28596 40354
rect 27710 40260 27750 40302
rect 28780 40302 28792 40460
rect 28792 40302 28820 40460
rect 28780 40260 28820 40302
rect 32700 40770 32740 40820
rect 32700 40612 32726 40770
rect 32726 40612 32740 40770
rect 33770 40770 33810 40820
rect 32912 40718 33088 40752
rect 33410 40718 33586 40752
rect 32828 40674 32862 40708
rect 33645 40674 33679 40708
rect 32912 40630 33088 40664
rect 33410 40630 33586 40664
rect 32700 40560 32740 40612
rect 32700 40460 32740 40500
rect 32700 40302 32726 40460
rect 32726 40302 32740 40460
rect 33770 40612 33782 40770
rect 33782 40612 33810 40770
rect 33770 40580 33810 40612
rect 33770 40460 33810 40500
rect 32912 40408 33088 40442
rect 33410 40408 33586 40442
rect 32828 40364 32862 40398
rect 33645 40364 33679 40398
rect 32912 40320 33088 40354
rect 33410 40320 33586 40354
rect 32700 40260 32740 40302
rect 33770 40302 33782 40460
rect 33782 40302 33810 40460
rect 33770 40260 33810 40302
rect 37690 40770 37730 40820
rect 37690 40612 37716 40770
rect 37716 40612 37730 40770
rect 38760 40770 38800 40820
rect 37902 40718 38078 40752
rect 38400 40718 38576 40752
rect 37818 40674 37852 40708
rect 38635 40674 38669 40708
rect 37902 40630 38078 40664
rect 38400 40630 38576 40664
rect 37690 40560 37730 40612
rect 37690 40460 37730 40500
rect 37690 40302 37716 40460
rect 37716 40302 37730 40460
rect 38760 40612 38772 40770
rect 38772 40612 38800 40770
rect 38760 40580 38800 40612
rect 38760 40460 38800 40500
rect 37902 40408 38078 40442
rect 38400 40408 38576 40442
rect 37818 40364 37852 40398
rect 38635 40364 38669 40398
rect 37902 40320 38078 40354
rect 38400 40320 38576 40354
rect 37690 40260 37730 40302
rect 38760 40302 38772 40460
rect 38772 40302 38800 40460
rect 38760 40260 38800 40302
rect 42680 40770 42720 40820
rect 42680 40612 42706 40770
rect 42706 40612 42720 40770
rect 43750 40770 43790 40820
rect 42892 40718 43068 40752
rect 43390 40718 43566 40752
rect 42808 40674 42842 40708
rect 43625 40674 43659 40708
rect 42892 40630 43068 40664
rect 43390 40630 43566 40664
rect 42680 40560 42720 40612
rect 42680 40460 42720 40500
rect 42680 40302 42706 40460
rect 42706 40302 42720 40460
rect 43750 40612 43762 40770
rect 43762 40612 43790 40770
rect 43750 40580 43790 40612
rect 43750 40460 43790 40500
rect 42892 40408 43068 40442
rect 43390 40408 43566 40442
rect 42808 40364 42842 40398
rect 43625 40364 43659 40398
rect 42892 40320 43068 40354
rect 43390 40320 43566 40354
rect 42680 40260 42720 40302
rect 43750 40302 43762 40460
rect 43762 40302 43790 40460
rect 43750 40260 43790 40302
rect 47670 40770 47710 40820
rect 47670 40612 47696 40770
rect 47696 40612 47710 40770
rect 48740 40770 48780 40820
rect 47882 40718 48058 40752
rect 48380 40718 48556 40752
rect 47798 40674 47832 40708
rect 48615 40674 48649 40708
rect 47882 40630 48058 40664
rect 48380 40630 48556 40664
rect 47670 40560 47710 40612
rect 47670 40460 47710 40500
rect 47670 40302 47696 40460
rect 47696 40302 47710 40460
rect 48740 40612 48752 40770
rect 48752 40612 48780 40770
rect 48740 40580 48780 40612
rect 48740 40460 48780 40500
rect 47882 40408 48058 40442
rect 48380 40408 48556 40442
rect 47798 40364 47832 40398
rect 48615 40364 48649 40398
rect 47882 40320 48058 40354
rect 48380 40320 48556 40354
rect 47670 40260 47710 40302
rect 48740 40302 48752 40460
rect 48752 40302 48780 40460
rect 48740 40260 48780 40302
rect 52660 40770 52700 40820
rect 52660 40612 52686 40770
rect 52686 40612 52700 40770
rect 53730 40770 53770 40820
rect 52872 40718 53048 40752
rect 53370 40718 53546 40752
rect 52788 40674 52822 40708
rect 53605 40674 53639 40708
rect 52872 40630 53048 40664
rect 53370 40630 53546 40664
rect 52660 40560 52700 40612
rect 52660 40460 52700 40500
rect 52660 40302 52686 40460
rect 52686 40302 52700 40460
rect 53730 40612 53742 40770
rect 53742 40612 53770 40770
rect 53730 40580 53770 40612
rect 53730 40460 53770 40500
rect 52872 40408 53048 40442
rect 53370 40408 53546 40442
rect 52788 40364 52822 40398
rect 53605 40364 53639 40398
rect 52872 40320 53048 40354
rect 53370 40320 53546 40354
rect 52660 40260 52700 40302
rect 53730 40302 53742 40460
rect 53742 40302 53770 40460
rect 53730 40260 53770 40302
rect 57650 40770 57690 40820
rect 57650 40612 57676 40770
rect 57676 40612 57690 40770
rect 58720 40770 58760 40820
rect 57862 40718 58038 40752
rect 58360 40718 58536 40752
rect 57778 40674 57812 40708
rect 58595 40674 58629 40708
rect 57862 40630 58038 40664
rect 58360 40630 58536 40664
rect 57650 40560 57690 40612
rect 57650 40460 57690 40500
rect 57650 40302 57676 40460
rect 57676 40302 57690 40460
rect 58720 40612 58732 40770
rect 58732 40612 58760 40770
rect 58720 40580 58760 40612
rect 58720 40460 58760 40500
rect 57862 40408 58038 40442
rect 58360 40408 58536 40442
rect 57778 40364 57812 40398
rect 58595 40364 58629 40398
rect 57862 40320 58038 40354
rect 58360 40320 58536 40354
rect 57650 40260 57690 40302
rect 58720 40302 58732 40460
rect 58732 40302 58760 40460
rect 58720 40260 58760 40302
rect 62640 40770 62680 40820
rect 62640 40612 62666 40770
rect 62666 40612 62680 40770
rect 63710 40770 63750 40820
rect 62852 40718 63028 40752
rect 63350 40718 63526 40752
rect 62768 40674 62802 40708
rect 63585 40674 63619 40708
rect 62852 40630 63028 40664
rect 63350 40630 63526 40664
rect 62640 40560 62680 40612
rect 62640 40460 62680 40500
rect 62640 40302 62666 40460
rect 62666 40302 62680 40460
rect 63710 40612 63722 40770
rect 63722 40612 63750 40770
rect 63710 40580 63750 40612
rect 63710 40460 63750 40500
rect 62852 40408 63028 40442
rect 63350 40408 63526 40442
rect 62768 40364 62802 40398
rect 63585 40364 63619 40398
rect 62852 40320 63028 40354
rect 63350 40320 63526 40354
rect 62640 40260 62680 40302
rect 63710 40302 63722 40460
rect 63722 40302 63750 40460
rect 63710 40260 63750 40302
rect 67630 40770 67670 40820
rect 67630 40612 67656 40770
rect 67656 40612 67670 40770
rect 68700 40770 68740 40820
rect 67842 40718 68018 40752
rect 68340 40718 68516 40752
rect 67758 40674 67792 40708
rect 68575 40674 68609 40708
rect 67842 40630 68018 40664
rect 68340 40630 68516 40664
rect 67630 40560 67670 40612
rect 67630 40460 67670 40500
rect 67630 40302 67656 40460
rect 67656 40302 67670 40460
rect 68700 40612 68712 40770
rect 68712 40612 68740 40770
rect 68700 40580 68740 40612
rect 68700 40460 68740 40500
rect 67842 40408 68018 40442
rect 68340 40408 68516 40442
rect 67758 40364 67792 40398
rect 68575 40364 68609 40398
rect 67842 40320 68018 40354
rect 68340 40320 68516 40354
rect 67630 40260 67670 40302
rect 68700 40302 68712 40460
rect 68712 40302 68740 40460
rect 68700 40260 68740 40302
rect 72620 40770 72660 40820
rect 72620 40612 72646 40770
rect 72646 40612 72660 40770
rect 73690 40770 73730 40820
rect 72832 40718 73008 40752
rect 73330 40718 73506 40752
rect 72748 40674 72782 40708
rect 73565 40674 73599 40708
rect 72832 40630 73008 40664
rect 73330 40630 73506 40664
rect 72620 40560 72660 40612
rect 72620 40460 72660 40500
rect 72620 40302 72646 40460
rect 72646 40302 72660 40460
rect 73690 40612 73702 40770
rect 73702 40612 73730 40770
rect 73690 40580 73730 40612
rect 73690 40460 73730 40500
rect 72832 40408 73008 40442
rect 73330 40408 73506 40442
rect 72748 40364 72782 40398
rect 73565 40364 73599 40398
rect 72832 40320 73008 40354
rect 73330 40320 73506 40354
rect 72620 40260 72660 40302
rect 73690 40302 73702 40460
rect 73702 40302 73730 40460
rect 73690 40260 73730 40302
rect 77610 40770 77650 40820
rect 77610 40612 77636 40770
rect 77636 40612 77650 40770
rect 78680 40770 78720 40820
rect 77822 40718 77998 40752
rect 78320 40718 78496 40752
rect 77738 40674 77772 40708
rect 78555 40674 78589 40708
rect 77822 40630 77998 40664
rect 78320 40630 78496 40664
rect 77610 40560 77650 40612
rect 77610 40460 77650 40500
rect 77610 40302 77636 40460
rect 77636 40302 77650 40460
rect 78680 40612 78692 40770
rect 78692 40612 78720 40770
rect 78680 40580 78720 40612
rect 78680 40460 78720 40500
rect 77822 40408 77998 40442
rect 78320 40408 78496 40442
rect 77738 40364 77772 40398
rect 78555 40364 78589 40398
rect 77822 40320 77998 40354
rect 78320 40320 78496 40354
rect 77610 40260 77650 40302
rect 78680 40302 78692 40460
rect 78692 40302 78720 40460
rect 78680 40260 78720 40302
<< metal1 >>
rect -9740 35752 -1824 53786
rect 1960 39690 1990 67050
rect 2080 39690 2110 67050
rect 2200 39690 2230 67050
rect 2320 39690 2350 67050
rect 2440 39690 2470 67050
rect 2560 39690 2590 67050
rect 2680 66390 2710 67050
rect 2650 66380 2710 66390
rect 2650 66310 2710 66320
rect 2680 64680 2710 66310
rect 2650 64670 2710 64680
rect 2650 64600 2710 64610
rect 2680 62970 2710 64600
rect 2650 62960 2710 62970
rect 2650 62890 2710 62900
rect 2680 61260 2710 62890
rect 2650 61250 2710 61260
rect 2650 61180 2710 61190
rect 2680 59550 2710 61180
rect 2650 59540 2710 59550
rect 2650 59470 2710 59480
rect 2680 57840 2710 59470
rect 2650 57830 2710 57840
rect 2650 57760 2710 57770
rect 2680 56130 2710 57760
rect 2650 56120 2710 56130
rect 2650 56050 2710 56060
rect 2680 54420 2710 56050
rect 2650 54410 2710 54420
rect 2650 54340 2710 54350
rect 2680 52710 2710 54340
rect 2650 52700 2710 52710
rect 2650 52630 2710 52640
rect 2680 51000 2710 52630
rect 2650 50990 2710 51000
rect 2650 50920 2710 50930
rect 2680 49290 2710 50920
rect 2650 49280 2710 49290
rect 2650 49210 2710 49220
rect 2680 47580 2710 49210
rect 2650 47570 2710 47580
rect 2650 47500 2710 47510
rect 2680 45870 2710 47500
rect 2650 45860 2710 45870
rect 2650 45790 2710 45800
rect 2680 44160 2710 45790
rect 2650 44150 2710 44160
rect 2650 44080 2710 44090
rect 2680 42450 2710 44080
rect 2650 42440 2710 42450
rect 2650 42370 2710 42380
rect 2680 40740 2710 42370
rect 2650 40730 2710 40740
rect 2650 40660 2710 40670
rect 2680 39240 2710 40660
rect 2740 66470 2810 67050
rect 2740 66210 2760 66470
rect 2800 66210 2810 66470
rect 3820 66470 3890 67050
rect 3270 66440 3350 66450
rect 2960 66402 3160 66408
rect 2850 66370 2930 66390
rect 2850 66310 2860 66370
rect 2920 66358 2930 66370
rect 2960 66368 2972 66402
rect 3148 66400 3160 66402
rect 3270 66400 3280 66440
rect 3148 66380 3280 66400
rect 3340 66400 3350 66440
rect 3458 66402 3658 66408
rect 3458 66400 3470 66402
rect 3340 66380 3470 66400
rect 3148 66370 3470 66380
rect 3148 66368 3160 66370
rect 2960 66362 3160 66368
rect 3458 66368 3470 66370
rect 3646 66368 3658 66402
rect 3458 66362 3658 66368
rect 3690 66370 3770 66390
rect 2922 66324 2930 66358
rect 2920 66310 2930 66324
rect 2850 66290 2930 66310
rect 2960 66314 3160 66320
rect 2960 66280 2972 66314
rect 3148 66310 3160 66314
rect 3458 66314 3658 66320
rect 3458 66310 3470 66314
rect 3148 66280 3470 66310
rect 3646 66280 3658 66314
rect 3690 66310 3700 66370
rect 3760 66310 3770 66370
rect 3690 66290 3770 66310
rect 2960 66274 3160 66280
rect 2740 66150 2810 66210
rect 2740 65910 2760 66150
rect 2800 65910 2810 66150
rect 3270 66270 3350 66280
rect 3458 66274 3658 66280
rect 3270 66210 3280 66270
rect 3340 66210 3350 66270
rect 3270 66160 3350 66210
rect 3270 66100 3280 66160
rect 3340 66100 3350 66160
rect 2960 66092 3160 66098
rect 2850 66060 2930 66080
rect 2850 66000 2860 66060
rect 2920 66048 2930 66060
rect 2960 66058 2972 66092
rect 3148 66090 3160 66092
rect 3270 66090 3350 66100
rect 3820 66230 3830 66470
rect 3870 66230 3890 66470
rect 3820 66150 3890 66230
rect 3458 66092 3658 66098
rect 3458 66090 3470 66092
rect 3148 66060 3470 66090
rect 3148 66058 3160 66060
rect 2960 66052 3160 66058
rect 3458 66058 3470 66060
rect 3646 66058 3658 66092
rect 3458 66052 3658 66058
rect 3690 66060 3770 66080
rect 2922 66014 2930 66048
rect 2920 66000 2930 66014
rect 2850 65980 2930 66000
rect 2960 66004 3160 66010
rect 2960 65970 2972 66004
rect 3148 66000 3160 66004
rect 3458 66004 3658 66010
rect 3458 66000 3470 66004
rect 3148 65990 3470 66000
rect 3148 65970 3280 65990
rect 2960 65964 3160 65970
rect 3270 65930 3280 65970
rect 3340 65970 3470 65990
rect 3646 65970 3658 66004
rect 3690 66000 3700 66060
rect 3760 66000 3770 66060
rect 3690 65980 3770 66000
rect 3340 65930 3350 65970
rect 3458 65964 3658 65970
rect 3270 65920 3350 65930
rect 2740 64760 2810 65910
rect 2740 64500 2760 64760
rect 2800 64500 2810 64760
rect 3820 65910 3830 66150
rect 3870 65910 3890 66150
rect 3820 64760 3890 65910
rect 3270 64730 3350 64740
rect 2960 64692 3160 64698
rect 2850 64660 2930 64680
rect 2850 64600 2860 64660
rect 2920 64648 2930 64660
rect 2960 64658 2972 64692
rect 3148 64690 3160 64692
rect 3270 64690 3280 64730
rect 3148 64670 3280 64690
rect 3340 64690 3350 64730
rect 3458 64692 3658 64698
rect 3458 64690 3470 64692
rect 3340 64670 3470 64690
rect 3148 64660 3470 64670
rect 3148 64658 3160 64660
rect 2960 64652 3160 64658
rect 3458 64658 3470 64660
rect 3646 64658 3658 64692
rect 3458 64652 3658 64658
rect 3690 64660 3770 64680
rect 2922 64614 2930 64648
rect 2920 64600 2930 64614
rect 2850 64580 2930 64600
rect 2960 64604 3160 64610
rect 2960 64570 2972 64604
rect 3148 64600 3160 64604
rect 3458 64604 3658 64610
rect 3458 64600 3470 64604
rect 3148 64570 3470 64600
rect 3646 64570 3658 64604
rect 3690 64600 3700 64660
rect 3760 64600 3770 64660
rect 3690 64580 3770 64600
rect 2960 64564 3160 64570
rect 2740 64440 2810 64500
rect 2740 64200 2760 64440
rect 2800 64200 2810 64440
rect 3270 64560 3350 64570
rect 3458 64564 3658 64570
rect 3270 64500 3280 64560
rect 3340 64500 3350 64560
rect 3270 64450 3350 64500
rect 3270 64390 3280 64450
rect 3340 64390 3350 64450
rect 2960 64382 3160 64388
rect 2850 64350 2930 64370
rect 2850 64290 2860 64350
rect 2920 64338 2930 64350
rect 2960 64348 2972 64382
rect 3148 64380 3160 64382
rect 3270 64380 3350 64390
rect 3820 64520 3830 64760
rect 3870 64520 3890 64760
rect 3820 64440 3890 64520
rect 3458 64382 3658 64388
rect 3458 64380 3470 64382
rect 3148 64350 3470 64380
rect 3148 64348 3160 64350
rect 2960 64342 3160 64348
rect 3458 64348 3470 64350
rect 3646 64348 3658 64382
rect 3458 64342 3658 64348
rect 3690 64350 3770 64370
rect 2922 64304 2930 64338
rect 2920 64290 2930 64304
rect 2850 64270 2930 64290
rect 2960 64294 3160 64300
rect 2960 64260 2972 64294
rect 3148 64290 3160 64294
rect 3458 64294 3658 64300
rect 3458 64290 3470 64294
rect 3148 64280 3470 64290
rect 3148 64260 3280 64280
rect 2960 64254 3160 64260
rect 3270 64220 3280 64260
rect 3340 64260 3470 64280
rect 3646 64260 3658 64294
rect 3690 64290 3700 64350
rect 3760 64290 3770 64350
rect 3690 64270 3770 64290
rect 3340 64220 3350 64260
rect 3458 64254 3658 64260
rect 3270 64210 3350 64220
rect 2740 63050 2810 64200
rect 2740 62790 2760 63050
rect 2800 62790 2810 63050
rect 3820 64200 3830 64440
rect 3870 64200 3890 64440
rect 3820 63050 3890 64200
rect 3270 63020 3350 63030
rect 2960 62982 3160 62988
rect 2850 62950 2930 62970
rect 2850 62890 2860 62950
rect 2920 62938 2930 62950
rect 2960 62948 2972 62982
rect 3148 62980 3160 62982
rect 3270 62980 3280 63020
rect 3148 62960 3280 62980
rect 3340 62980 3350 63020
rect 3458 62982 3658 62988
rect 3458 62980 3470 62982
rect 3340 62960 3470 62980
rect 3148 62950 3470 62960
rect 3148 62948 3160 62950
rect 2960 62942 3160 62948
rect 3458 62948 3470 62950
rect 3646 62948 3658 62982
rect 3458 62942 3658 62948
rect 3690 62950 3770 62970
rect 2922 62904 2930 62938
rect 2920 62890 2930 62904
rect 2850 62870 2930 62890
rect 2960 62894 3160 62900
rect 2960 62860 2972 62894
rect 3148 62890 3160 62894
rect 3458 62894 3658 62900
rect 3458 62890 3470 62894
rect 3148 62860 3470 62890
rect 3646 62860 3658 62894
rect 3690 62890 3700 62950
rect 3760 62890 3770 62950
rect 3690 62870 3770 62890
rect 2960 62854 3160 62860
rect 2740 62730 2810 62790
rect 2740 62490 2760 62730
rect 2800 62490 2810 62730
rect 3270 62850 3350 62860
rect 3458 62854 3658 62860
rect 3270 62790 3280 62850
rect 3340 62790 3350 62850
rect 3270 62740 3350 62790
rect 3270 62680 3280 62740
rect 3340 62680 3350 62740
rect 2960 62672 3160 62678
rect 2850 62640 2930 62660
rect 2850 62580 2860 62640
rect 2920 62628 2930 62640
rect 2960 62638 2972 62672
rect 3148 62670 3160 62672
rect 3270 62670 3350 62680
rect 3820 62810 3830 63050
rect 3870 62810 3890 63050
rect 3820 62730 3890 62810
rect 3458 62672 3658 62678
rect 3458 62670 3470 62672
rect 3148 62640 3470 62670
rect 3148 62638 3160 62640
rect 2960 62632 3160 62638
rect 3458 62638 3470 62640
rect 3646 62638 3658 62672
rect 3458 62632 3658 62638
rect 3690 62640 3770 62660
rect 2922 62594 2930 62628
rect 2920 62580 2930 62594
rect 2850 62560 2930 62580
rect 2960 62584 3160 62590
rect 2960 62550 2972 62584
rect 3148 62580 3160 62584
rect 3458 62584 3658 62590
rect 3458 62580 3470 62584
rect 3148 62570 3470 62580
rect 3148 62550 3280 62570
rect 2960 62544 3160 62550
rect 3270 62510 3280 62550
rect 3340 62550 3470 62570
rect 3646 62550 3658 62584
rect 3690 62580 3700 62640
rect 3760 62580 3770 62640
rect 3690 62560 3770 62580
rect 3340 62510 3350 62550
rect 3458 62544 3658 62550
rect 3270 62500 3350 62510
rect 2740 61340 2810 62490
rect 2740 61080 2760 61340
rect 2800 61080 2810 61340
rect 3820 62490 3830 62730
rect 3870 62490 3890 62730
rect 3820 61340 3890 62490
rect 3270 61310 3350 61320
rect 2960 61272 3160 61278
rect 2850 61240 2930 61260
rect 2850 61180 2860 61240
rect 2920 61228 2930 61240
rect 2960 61238 2972 61272
rect 3148 61270 3160 61272
rect 3270 61270 3280 61310
rect 3148 61250 3280 61270
rect 3340 61270 3350 61310
rect 3458 61272 3658 61278
rect 3458 61270 3470 61272
rect 3340 61250 3470 61270
rect 3148 61240 3470 61250
rect 3148 61238 3160 61240
rect 2960 61232 3160 61238
rect 3458 61238 3470 61240
rect 3646 61238 3658 61272
rect 3458 61232 3658 61238
rect 3690 61240 3770 61260
rect 2922 61194 2930 61228
rect 2920 61180 2930 61194
rect 2850 61160 2930 61180
rect 2960 61184 3160 61190
rect 2960 61150 2972 61184
rect 3148 61180 3160 61184
rect 3458 61184 3658 61190
rect 3458 61180 3470 61184
rect 3148 61150 3470 61180
rect 3646 61150 3658 61184
rect 3690 61180 3700 61240
rect 3760 61180 3770 61240
rect 3690 61160 3770 61180
rect 2960 61144 3160 61150
rect 2740 61020 2810 61080
rect 2740 60780 2760 61020
rect 2800 60780 2810 61020
rect 3270 61140 3350 61150
rect 3458 61144 3658 61150
rect 3270 61080 3280 61140
rect 3340 61080 3350 61140
rect 3270 61030 3350 61080
rect 3270 60970 3280 61030
rect 3340 60970 3350 61030
rect 2960 60962 3160 60968
rect 2850 60930 2930 60950
rect 2850 60870 2860 60930
rect 2920 60918 2930 60930
rect 2960 60928 2972 60962
rect 3148 60960 3160 60962
rect 3270 60960 3350 60970
rect 3820 61100 3830 61340
rect 3870 61100 3890 61340
rect 3820 61020 3890 61100
rect 3458 60962 3658 60968
rect 3458 60960 3470 60962
rect 3148 60930 3470 60960
rect 3148 60928 3160 60930
rect 2960 60922 3160 60928
rect 3458 60928 3470 60930
rect 3646 60928 3658 60962
rect 3458 60922 3658 60928
rect 3690 60930 3770 60950
rect 2922 60884 2930 60918
rect 2920 60870 2930 60884
rect 2850 60850 2930 60870
rect 2960 60874 3160 60880
rect 2960 60840 2972 60874
rect 3148 60870 3160 60874
rect 3458 60874 3658 60880
rect 3458 60870 3470 60874
rect 3148 60860 3470 60870
rect 3148 60840 3280 60860
rect 2960 60834 3160 60840
rect 3270 60800 3280 60840
rect 3340 60840 3470 60860
rect 3646 60840 3658 60874
rect 3690 60870 3700 60930
rect 3760 60870 3770 60930
rect 3690 60850 3770 60870
rect 3340 60800 3350 60840
rect 3458 60834 3658 60840
rect 3270 60790 3350 60800
rect 2740 59630 2810 60780
rect 2740 59370 2760 59630
rect 2800 59370 2810 59630
rect 3820 60780 3830 61020
rect 3870 60780 3890 61020
rect 3820 59630 3890 60780
rect 3270 59600 3350 59610
rect 2960 59562 3160 59568
rect 2850 59530 2930 59550
rect 2850 59470 2860 59530
rect 2920 59518 2930 59530
rect 2960 59528 2972 59562
rect 3148 59560 3160 59562
rect 3270 59560 3280 59600
rect 3148 59540 3280 59560
rect 3340 59560 3350 59600
rect 3458 59562 3658 59568
rect 3458 59560 3470 59562
rect 3340 59540 3470 59560
rect 3148 59530 3470 59540
rect 3148 59528 3160 59530
rect 2960 59522 3160 59528
rect 3458 59528 3470 59530
rect 3646 59528 3658 59562
rect 3458 59522 3658 59528
rect 3690 59530 3770 59550
rect 2922 59484 2930 59518
rect 2920 59470 2930 59484
rect 2850 59450 2930 59470
rect 2960 59474 3160 59480
rect 2960 59440 2972 59474
rect 3148 59470 3160 59474
rect 3458 59474 3658 59480
rect 3458 59470 3470 59474
rect 3148 59440 3470 59470
rect 3646 59440 3658 59474
rect 3690 59470 3700 59530
rect 3760 59470 3770 59530
rect 3690 59450 3770 59470
rect 2960 59434 3160 59440
rect 2740 59310 2810 59370
rect 2740 59070 2760 59310
rect 2800 59070 2810 59310
rect 3270 59430 3350 59440
rect 3458 59434 3658 59440
rect 3270 59370 3280 59430
rect 3340 59370 3350 59430
rect 3270 59320 3350 59370
rect 3270 59260 3280 59320
rect 3340 59260 3350 59320
rect 2960 59252 3160 59258
rect 2850 59220 2930 59240
rect 2850 59160 2860 59220
rect 2920 59208 2930 59220
rect 2960 59218 2972 59252
rect 3148 59250 3160 59252
rect 3270 59250 3350 59260
rect 3820 59390 3830 59630
rect 3870 59390 3890 59630
rect 3820 59310 3890 59390
rect 3458 59252 3658 59258
rect 3458 59250 3470 59252
rect 3148 59220 3470 59250
rect 3148 59218 3160 59220
rect 2960 59212 3160 59218
rect 3458 59218 3470 59220
rect 3646 59218 3658 59252
rect 3458 59212 3658 59218
rect 3690 59220 3770 59240
rect 2922 59174 2930 59208
rect 2920 59160 2930 59174
rect 2850 59140 2930 59160
rect 2960 59164 3160 59170
rect 2960 59130 2972 59164
rect 3148 59160 3160 59164
rect 3458 59164 3658 59170
rect 3458 59160 3470 59164
rect 3148 59150 3470 59160
rect 3148 59130 3280 59150
rect 2960 59124 3160 59130
rect 3270 59090 3280 59130
rect 3340 59130 3470 59150
rect 3646 59130 3658 59164
rect 3690 59160 3700 59220
rect 3760 59160 3770 59220
rect 3690 59140 3770 59160
rect 3340 59090 3350 59130
rect 3458 59124 3658 59130
rect 3270 59080 3350 59090
rect 2740 57920 2810 59070
rect 2740 57660 2760 57920
rect 2800 57660 2810 57920
rect 3820 59070 3830 59310
rect 3870 59070 3890 59310
rect 3820 57920 3890 59070
rect 3270 57890 3350 57900
rect 2960 57852 3160 57858
rect 2850 57820 2930 57840
rect 2850 57760 2860 57820
rect 2920 57808 2930 57820
rect 2960 57818 2972 57852
rect 3148 57850 3160 57852
rect 3270 57850 3280 57890
rect 3148 57830 3280 57850
rect 3340 57850 3350 57890
rect 3458 57852 3658 57858
rect 3458 57850 3470 57852
rect 3340 57830 3470 57850
rect 3148 57820 3470 57830
rect 3148 57818 3160 57820
rect 2960 57812 3160 57818
rect 3458 57818 3470 57820
rect 3646 57818 3658 57852
rect 3458 57812 3658 57818
rect 3690 57820 3770 57840
rect 2922 57774 2930 57808
rect 2920 57760 2930 57774
rect 2850 57740 2930 57760
rect 2960 57764 3160 57770
rect 2960 57730 2972 57764
rect 3148 57760 3160 57764
rect 3458 57764 3658 57770
rect 3458 57760 3470 57764
rect 3148 57730 3470 57760
rect 3646 57730 3658 57764
rect 3690 57760 3700 57820
rect 3760 57760 3770 57820
rect 3690 57740 3770 57760
rect 2960 57724 3160 57730
rect 2740 57600 2810 57660
rect 2740 57360 2760 57600
rect 2800 57360 2810 57600
rect 3270 57720 3350 57730
rect 3458 57724 3658 57730
rect 3270 57660 3280 57720
rect 3340 57660 3350 57720
rect 3270 57610 3350 57660
rect 3270 57550 3280 57610
rect 3340 57550 3350 57610
rect 2960 57542 3160 57548
rect 2850 57510 2930 57530
rect 2850 57450 2860 57510
rect 2920 57498 2930 57510
rect 2960 57508 2972 57542
rect 3148 57540 3160 57542
rect 3270 57540 3350 57550
rect 3820 57680 3830 57920
rect 3870 57680 3890 57920
rect 3820 57600 3890 57680
rect 3458 57542 3658 57548
rect 3458 57540 3470 57542
rect 3148 57510 3470 57540
rect 3148 57508 3160 57510
rect 2960 57502 3160 57508
rect 3458 57508 3470 57510
rect 3646 57508 3658 57542
rect 3458 57502 3658 57508
rect 3690 57510 3770 57530
rect 2922 57464 2930 57498
rect 2920 57450 2930 57464
rect 2850 57430 2930 57450
rect 2960 57454 3160 57460
rect 2960 57420 2972 57454
rect 3148 57450 3160 57454
rect 3458 57454 3658 57460
rect 3458 57450 3470 57454
rect 3148 57440 3470 57450
rect 3148 57420 3280 57440
rect 2960 57414 3160 57420
rect 3270 57380 3280 57420
rect 3340 57420 3470 57440
rect 3646 57420 3658 57454
rect 3690 57450 3700 57510
rect 3760 57450 3770 57510
rect 3690 57430 3770 57450
rect 3340 57380 3350 57420
rect 3458 57414 3658 57420
rect 3270 57370 3350 57380
rect 2740 56210 2810 57360
rect 2740 55950 2760 56210
rect 2800 55950 2810 56210
rect 3820 57360 3830 57600
rect 3870 57360 3890 57600
rect 3820 56210 3890 57360
rect 3270 56180 3350 56190
rect 2960 56142 3160 56148
rect 2850 56110 2930 56130
rect 2850 56050 2860 56110
rect 2920 56098 2930 56110
rect 2960 56108 2972 56142
rect 3148 56140 3160 56142
rect 3270 56140 3280 56180
rect 3148 56120 3280 56140
rect 3340 56140 3350 56180
rect 3458 56142 3658 56148
rect 3458 56140 3470 56142
rect 3340 56120 3470 56140
rect 3148 56110 3470 56120
rect 3148 56108 3160 56110
rect 2960 56102 3160 56108
rect 3458 56108 3470 56110
rect 3646 56108 3658 56142
rect 3458 56102 3658 56108
rect 3690 56110 3770 56130
rect 2922 56064 2930 56098
rect 2920 56050 2930 56064
rect 2850 56030 2930 56050
rect 2960 56054 3160 56060
rect 2960 56020 2972 56054
rect 3148 56050 3160 56054
rect 3458 56054 3658 56060
rect 3458 56050 3470 56054
rect 3148 56020 3470 56050
rect 3646 56020 3658 56054
rect 3690 56050 3700 56110
rect 3760 56050 3770 56110
rect 3690 56030 3770 56050
rect 2960 56014 3160 56020
rect 2740 55890 2810 55950
rect 2740 55650 2760 55890
rect 2800 55650 2810 55890
rect 3270 56010 3350 56020
rect 3458 56014 3658 56020
rect 3270 55950 3280 56010
rect 3340 55950 3350 56010
rect 3270 55900 3350 55950
rect 3270 55840 3280 55900
rect 3340 55840 3350 55900
rect 2960 55832 3160 55838
rect 2850 55800 2930 55820
rect 2850 55740 2860 55800
rect 2920 55788 2930 55800
rect 2960 55798 2972 55832
rect 3148 55830 3160 55832
rect 3270 55830 3350 55840
rect 3820 55970 3830 56210
rect 3870 55970 3890 56210
rect 3820 55890 3890 55970
rect 3458 55832 3658 55838
rect 3458 55830 3470 55832
rect 3148 55800 3470 55830
rect 3148 55798 3160 55800
rect 2960 55792 3160 55798
rect 3458 55798 3470 55800
rect 3646 55798 3658 55832
rect 3458 55792 3658 55798
rect 3690 55800 3770 55820
rect 2922 55754 2930 55788
rect 2920 55740 2930 55754
rect 2850 55720 2930 55740
rect 2960 55744 3160 55750
rect 2960 55710 2972 55744
rect 3148 55740 3160 55744
rect 3458 55744 3658 55750
rect 3458 55740 3470 55744
rect 3148 55730 3470 55740
rect 3148 55710 3280 55730
rect 2960 55704 3160 55710
rect 3270 55670 3280 55710
rect 3340 55710 3470 55730
rect 3646 55710 3658 55744
rect 3690 55740 3700 55800
rect 3760 55740 3770 55800
rect 3690 55720 3770 55740
rect 3340 55670 3350 55710
rect 3458 55704 3658 55710
rect 3270 55660 3350 55670
rect 2740 54500 2810 55650
rect 2740 54240 2760 54500
rect 2800 54240 2810 54500
rect 3820 55650 3830 55890
rect 3870 55650 3890 55890
rect 3820 54500 3890 55650
rect 3270 54470 3350 54480
rect 2960 54432 3160 54438
rect 2850 54400 2930 54420
rect 2850 54340 2860 54400
rect 2920 54388 2930 54400
rect 2960 54398 2972 54432
rect 3148 54430 3160 54432
rect 3270 54430 3280 54470
rect 3148 54410 3280 54430
rect 3340 54430 3350 54470
rect 3458 54432 3658 54438
rect 3458 54430 3470 54432
rect 3340 54410 3470 54430
rect 3148 54400 3470 54410
rect 3148 54398 3160 54400
rect 2960 54392 3160 54398
rect 3458 54398 3470 54400
rect 3646 54398 3658 54432
rect 3458 54392 3658 54398
rect 3690 54400 3770 54420
rect 2922 54354 2930 54388
rect 2920 54340 2930 54354
rect 2850 54320 2930 54340
rect 2960 54344 3160 54350
rect 2960 54310 2972 54344
rect 3148 54340 3160 54344
rect 3458 54344 3658 54350
rect 3458 54340 3470 54344
rect 3148 54310 3470 54340
rect 3646 54310 3658 54344
rect 3690 54340 3700 54400
rect 3760 54340 3770 54400
rect 3690 54320 3770 54340
rect 2960 54304 3160 54310
rect 2740 54180 2810 54240
rect 2740 53940 2760 54180
rect 2800 53940 2810 54180
rect 3270 54300 3350 54310
rect 3458 54304 3658 54310
rect 3270 54240 3280 54300
rect 3340 54240 3350 54300
rect 3270 54190 3350 54240
rect 3270 54130 3280 54190
rect 3340 54130 3350 54190
rect 2960 54122 3160 54128
rect 2850 54090 2930 54110
rect 2850 54030 2860 54090
rect 2920 54078 2930 54090
rect 2960 54088 2972 54122
rect 3148 54120 3160 54122
rect 3270 54120 3350 54130
rect 3820 54260 3830 54500
rect 3870 54260 3890 54500
rect 3820 54180 3890 54260
rect 3458 54122 3658 54128
rect 3458 54120 3470 54122
rect 3148 54090 3470 54120
rect 3148 54088 3160 54090
rect 2960 54082 3160 54088
rect 3458 54088 3470 54090
rect 3646 54088 3658 54122
rect 3458 54082 3658 54088
rect 3690 54090 3770 54110
rect 2922 54044 2930 54078
rect 2920 54030 2930 54044
rect 2850 54010 2930 54030
rect 2960 54034 3160 54040
rect 2960 54000 2972 54034
rect 3148 54030 3160 54034
rect 3458 54034 3658 54040
rect 3458 54030 3470 54034
rect 3148 54020 3470 54030
rect 3148 54000 3280 54020
rect 2960 53994 3160 54000
rect 3270 53960 3280 54000
rect 3340 54000 3470 54020
rect 3646 54000 3658 54034
rect 3690 54030 3700 54090
rect 3760 54030 3770 54090
rect 3690 54010 3770 54030
rect 3340 53960 3350 54000
rect 3458 53994 3658 54000
rect 3270 53950 3350 53960
rect 2740 52790 2810 53940
rect 2740 52530 2760 52790
rect 2800 52530 2810 52790
rect 3820 53940 3830 54180
rect 3870 53940 3890 54180
rect 3820 52790 3890 53940
rect 3270 52760 3350 52770
rect 2960 52722 3160 52728
rect 2850 52690 2930 52710
rect 2850 52630 2860 52690
rect 2920 52678 2930 52690
rect 2960 52688 2972 52722
rect 3148 52720 3160 52722
rect 3270 52720 3280 52760
rect 3148 52700 3280 52720
rect 3340 52720 3350 52760
rect 3458 52722 3658 52728
rect 3458 52720 3470 52722
rect 3340 52700 3470 52720
rect 3148 52690 3470 52700
rect 3148 52688 3160 52690
rect 2960 52682 3160 52688
rect 3458 52688 3470 52690
rect 3646 52688 3658 52722
rect 3458 52682 3658 52688
rect 3690 52690 3770 52710
rect 2922 52644 2930 52678
rect 2920 52630 2930 52644
rect 2850 52610 2930 52630
rect 2960 52634 3160 52640
rect 2960 52600 2972 52634
rect 3148 52630 3160 52634
rect 3458 52634 3658 52640
rect 3458 52630 3470 52634
rect 3148 52600 3470 52630
rect 3646 52600 3658 52634
rect 3690 52630 3700 52690
rect 3760 52630 3770 52690
rect 3690 52610 3770 52630
rect 2960 52594 3160 52600
rect 2740 52470 2810 52530
rect 2740 52230 2760 52470
rect 2800 52230 2810 52470
rect 3270 52590 3350 52600
rect 3458 52594 3658 52600
rect 3270 52530 3280 52590
rect 3340 52530 3350 52590
rect 3270 52480 3350 52530
rect 3270 52420 3280 52480
rect 3340 52420 3350 52480
rect 2960 52412 3160 52418
rect 2850 52380 2930 52400
rect 2850 52320 2860 52380
rect 2920 52368 2930 52380
rect 2960 52378 2972 52412
rect 3148 52410 3160 52412
rect 3270 52410 3350 52420
rect 3820 52550 3830 52790
rect 3870 52550 3890 52790
rect 3820 52470 3890 52550
rect 3458 52412 3658 52418
rect 3458 52410 3470 52412
rect 3148 52380 3470 52410
rect 3148 52378 3160 52380
rect 2960 52372 3160 52378
rect 3458 52378 3470 52380
rect 3646 52378 3658 52412
rect 3458 52372 3658 52378
rect 3690 52380 3770 52400
rect 2922 52334 2930 52368
rect 2920 52320 2930 52334
rect 2850 52300 2930 52320
rect 2960 52324 3160 52330
rect 2960 52290 2972 52324
rect 3148 52320 3160 52324
rect 3458 52324 3658 52330
rect 3458 52320 3470 52324
rect 3148 52310 3470 52320
rect 3148 52290 3280 52310
rect 2960 52284 3160 52290
rect 3270 52250 3280 52290
rect 3340 52290 3470 52310
rect 3646 52290 3658 52324
rect 3690 52320 3700 52380
rect 3760 52320 3770 52380
rect 3690 52300 3770 52320
rect 3340 52250 3350 52290
rect 3458 52284 3658 52290
rect 3270 52240 3350 52250
rect 2740 51080 2810 52230
rect 2740 50820 2760 51080
rect 2800 50820 2810 51080
rect 3820 52230 3830 52470
rect 3870 52230 3890 52470
rect 3820 51080 3890 52230
rect 3270 51050 3350 51060
rect 2960 51012 3160 51018
rect 2850 50980 2930 51000
rect 2850 50920 2860 50980
rect 2920 50968 2930 50980
rect 2960 50978 2972 51012
rect 3148 51010 3160 51012
rect 3270 51010 3280 51050
rect 3148 50990 3280 51010
rect 3340 51010 3350 51050
rect 3458 51012 3658 51018
rect 3458 51010 3470 51012
rect 3340 50990 3470 51010
rect 3148 50980 3470 50990
rect 3148 50978 3160 50980
rect 2960 50972 3160 50978
rect 3458 50978 3470 50980
rect 3646 50978 3658 51012
rect 3458 50972 3658 50978
rect 3690 50980 3770 51000
rect 2922 50934 2930 50968
rect 2920 50920 2930 50934
rect 2850 50900 2930 50920
rect 2960 50924 3160 50930
rect 2960 50890 2972 50924
rect 3148 50920 3160 50924
rect 3458 50924 3658 50930
rect 3458 50920 3470 50924
rect 3148 50890 3470 50920
rect 3646 50890 3658 50924
rect 3690 50920 3700 50980
rect 3760 50920 3770 50980
rect 3690 50900 3770 50920
rect 2960 50884 3160 50890
rect 2740 50760 2810 50820
rect 2740 50520 2760 50760
rect 2800 50520 2810 50760
rect 3270 50880 3350 50890
rect 3458 50884 3658 50890
rect 3270 50820 3280 50880
rect 3340 50820 3350 50880
rect 3270 50770 3350 50820
rect 3270 50710 3280 50770
rect 3340 50710 3350 50770
rect 2960 50702 3160 50708
rect 2850 50670 2930 50690
rect 2850 50610 2860 50670
rect 2920 50658 2930 50670
rect 2960 50668 2972 50702
rect 3148 50700 3160 50702
rect 3270 50700 3350 50710
rect 3820 50840 3830 51080
rect 3870 50840 3890 51080
rect 3820 50760 3890 50840
rect 3458 50702 3658 50708
rect 3458 50700 3470 50702
rect 3148 50670 3470 50700
rect 3148 50668 3160 50670
rect 2960 50662 3160 50668
rect 3458 50668 3470 50670
rect 3646 50668 3658 50702
rect 3458 50662 3658 50668
rect 3690 50670 3770 50690
rect 2922 50624 2930 50658
rect 2920 50610 2930 50624
rect 2850 50590 2930 50610
rect 2960 50614 3160 50620
rect 2960 50580 2972 50614
rect 3148 50610 3160 50614
rect 3458 50614 3658 50620
rect 3458 50610 3470 50614
rect 3148 50600 3470 50610
rect 3148 50580 3280 50600
rect 2960 50574 3160 50580
rect 3270 50540 3280 50580
rect 3340 50580 3470 50600
rect 3646 50580 3658 50614
rect 3690 50610 3700 50670
rect 3760 50610 3770 50670
rect 3690 50590 3770 50610
rect 3340 50540 3350 50580
rect 3458 50574 3658 50580
rect 3270 50530 3350 50540
rect 2740 49370 2810 50520
rect 2740 49110 2760 49370
rect 2800 49110 2810 49370
rect 3820 50520 3830 50760
rect 3870 50520 3890 50760
rect 3820 49370 3890 50520
rect 3270 49340 3350 49350
rect 2960 49302 3160 49308
rect 2850 49270 2930 49290
rect 2850 49210 2860 49270
rect 2920 49258 2930 49270
rect 2960 49268 2972 49302
rect 3148 49300 3160 49302
rect 3270 49300 3280 49340
rect 3148 49280 3280 49300
rect 3340 49300 3350 49340
rect 3458 49302 3658 49308
rect 3458 49300 3470 49302
rect 3340 49280 3470 49300
rect 3148 49270 3470 49280
rect 3148 49268 3160 49270
rect 2960 49262 3160 49268
rect 3458 49268 3470 49270
rect 3646 49268 3658 49302
rect 3458 49262 3658 49268
rect 3690 49270 3770 49290
rect 2922 49224 2930 49258
rect 2920 49210 2930 49224
rect 2850 49190 2930 49210
rect 2960 49214 3160 49220
rect 2960 49180 2972 49214
rect 3148 49210 3160 49214
rect 3458 49214 3658 49220
rect 3458 49210 3470 49214
rect 3148 49180 3470 49210
rect 3646 49180 3658 49214
rect 3690 49210 3700 49270
rect 3760 49210 3770 49270
rect 3690 49190 3770 49210
rect 2960 49174 3160 49180
rect 2740 49050 2810 49110
rect 2740 48810 2760 49050
rect 2800 48810 2810 49050
rect 3270 49170 3350 49180
rect 3458 49174 3658 49180
rect 3270 49110 3280 49170
rect 3340 49110 3350 49170
rect 3270 49060 3350 49110
rect 3270 49000 3280 49060
rect 3340 49000 3350 49060
rect 2960 48992 3160 48998
rect 2850 48960 2930 48980
rect 2850 48900 2860 48960
rect 2920 48948 2930 48960
rect 2960 48958 2972 48992
rect 3148 48990 3160 48992
rect 3270 48990 3350 49000
rect 3820 49130 3830 49370
rect 3870 49130 3890 49370
rect 3820 49050 3890 49130
rect 3458 48992 3658 48998
rect 3458 48990 3470 48992
rect 3148 48960 3470 48990
rect 3148 48958 3160 48960
rect 2960 48952 3160 48958
rect 3458 48958 3470 48960
rect 3646 48958 3658 48992
rect 3458 48952 3658 48958
rect 3690 48960 3770 48980
rect 2922 48914 2930 48948
rect 2920 48900 2930 48914
rect 2850 48880 2930 48900
rect 2960 48904 3160 48910
rect 2960 48870 2972 48904
rect 3148 48900 3160 48904
rect 3458 48904 3658 48910
rect 3458 48900 3470 48904
rect 3148 48890 3470 48900
rect 3148 48870 3280 48890
rect 2960 48864 3160 48870
rect 3270 48830 3280 48870
rect 3340 48870 3470 48890
rect 3646 48870 3658 48904
rect 3690 48900 3700 48960
rect 3760 48900 3770 48960
rect 3690 48880 3770 48900
rect 3340 48830 3350 48870
rect 3458 48864 3658 48870
rect 3270 48820 3350 48830
rect 2740 47660 2810 48810
rect 2740 47400 2760 47660
rect 2800 47400 2810 47660
rect 3820 48810 3830 49050
rect 3870 48810 3890 49050
rect 3820 47660 3890 48810
rect 3270 47630 3350 47640
rect 2960 47592 3160 47598
rect 2850 47560 2930 47580
rect 2850 47500 2860 47560
rect 2920 47548 2930 47560
rect 2960 47558 2972 47592
rect 3148 47590 3160 47592
rect 3270 47590 3280 47630
rect 3148 47570 3280 47590
rect 3340 47590 3350 47630
rect 3458 47592 3658 47598
rect 3458 47590 3470 47592
rect 3340 47570 3470 47590
rect 3148 47560 3470 47570
rect 3148 47558 3160 47560
rect 2960 47552 3160 47558
rect 3458 47558 3470 47560
rect 3646 47558 3658 47592
rect 3458 47552 3658 47558
rect 3690 47560 3770 47580
rect 2922 47514 2930 47548
rect 2920 47500 2930 47514
rect 2850 47480 2930 47500
rect 2960 47504 3160 47510
rect 2960 47470 2972 47504
rect 3148 47500 3160 47504
rect 3458 47504 3658 47510
rect 3458 47500 3470 47504
rect 3148 47470 3470 47500
rect 3646 47470 3658 47504
rect 3690 47500 3700 47560
rect 3760 47500 3770 47560
rect 3690 47480 3770 47500
rect 2960 47464 3160 47470
rect 2740 47340 2810 47400
rect 2740 47100 2760 47340
rect 2800 47100 2810 47340
rect 3270 47460 3350 47470
rect 3458 47464 3658 47470
rect 3270 47400 3280 47460
rect 3340 47400 3350 47460
rect 3270 47350 3350 47400
rect 3270 47290 3280 47350
rect 3340 47290 3350 47350
rect 2960 47282 3160 47288
rect 2850 47250 2930 47270
rect 2850 47190 2860 47250
rect 2920 47238 2930 47250
rect 2960 47248 2972 47282
rect 3148 47280 3160 47282
rect 3270 47280 3350 47290
rect 3820 47420 3830 47660
rect 3870 47420 3890 47660
rect 3820 47340 3890 47420
rect 3458 47282 3658 47288
rect 3458 47280 3470 47282
rect 3148 47250 3470 47280
rect 3148 47248 3160 47250
rect 2960 47242 3160 47248
rect 3458 47248 3470 47250
rect 3646 47248 3658 47282
rect 3458 47242 3658 47248
rect 3690 47250 3770 47270
rect 2922 47204 2930 47238
rect 2920 47190 2930 47204
rect 2850 47170 2930 47190
rect 2960 47194 3160 47200
rect 2960 47160 2972 47194
rect 3148 47190 3160 47194
rect 3458 47194 3658 47200
rect 3458 47190 3470 47194
rect 3148 47180 3470 47190
rect 3148 47160 3280 47180
rect 2960 47154 3160 47160
rect 3270 47120 3280 47160
rect 3340 47160 3470 47180
rect 3646 47160 3658 47194
rect 3690 47190 3700 47250
rect 3760 47190 3770 47250
rect 3690 47170 3770 47190
rect 3340 47120 3350 47160
rect 3458 47154 3658 47160
rect 3270 47110 3350 47120
rect 2740 45950 2810 47100
rect 2740 45690 2760 45950
rect 2800 45690 2810 45950
rect 3820 47100 3830 47340
rect 3870 47100 3890 47340
rect 3820 45950 3890 47100
rect 3270 45920 3350 45930
rect 2960 45882 3160 45888
rect 2850 45850 2930 45870
rect 2850 45790 2860 45850
rect 2920 45838 2930 45850
rect 2960 45848 2972 45882
rect 3148 45880 3160 45882
rect 3270 45880 3280 45920
rect 3148 45860 3280 45880
rect 3340 45880 3350 45920
rect 3458 45882 3658 45888
rect 3458 45880 3470 45882
rect 3340 45860 3470 45880
rect 3148 45850 3470 45860
rect 3148 45848 3160 45850
rect 2960 45842 3160 45848
rect 3458 45848 3470 45850
rect 3646 45848 3658 45882
rect 3458 45842 3658 45848
rect 3690 45850 3770 45870
rect 2922 45804 2930 45838
rect 2920 45790 2930 45804
rect 2850 45770 2930 45790
rect 2960 45794 3160 45800
rect 2960 45760 2972 45794
rect 3148 45790 3160 45794
rect 3458 45794 3658 45800
rect 3458 45790 3470 45794
rect 3148 45760 3470 45790
rect 3646 45760 3658 45794
rect 3690 45790 3700 45850
rect 3760 45790 3770 45850
rect 3690 45770 3770 45790
rect 2960 45754 3160 45760
rect 2740 45630 2810 45690
rect 2740 45390 2760 45630
rect 2800 45390 2810 45630
rect 3270 45750 3350 45760
rect 3458 45754 3658 45760
rect 3270 45690 3280 45750
rect 3340 45690 3350 45750
rect 3270 45640 3350 45690
rect 3270 45580 3280 45640
rect 3340 45580 3350 45640
rect 2960 45572 3160 45578
rect 2850 45540 2930 45560
rect 2850 45480 2860 45540
rect 2920 45528 2930 45540
rect 2960 45538 2972 45572
rect 3148 45570 3160 45572
rect 3270 45570 3350 45580
rect 3820 45710 3830 45950
rect 3870 45710 3890 45950
rect 3820 45630 3890 45710
rect 3458 45572 3658 45578
rect 3458 45570 3470 45572
rect 3148 45540 3470 45570
rect 3148 45538 3160 45540
rect 2960 45532 3160 45538
rect 3458 45538 3470 45540
rect 3646 45538 3658 45572
rect 3458 45532 3658 45538
rect 3690 45540 3770 45560
rect 2922 45494 2930 45528
rect 2920 45480 2930 45494
rect 2850 45460 2930 45480
rect 2960 45484 3160 45490
rect 2960 45450 2972 45484
rect 3148 45480 3160 45484
rect 3458 45484 3658 45490
rect 3458 45480 3470 45484
rect 3148 45470 3470 45480
rect 3148 45450 3280 45470
rect 2960 45444 3160 45450
rect 3270 45410 3280 45450
rect 3340 45450 3470 45470
rect 3646 45450 3658 45484
rect 3690 45480 3700 45540
rect 3760 45480 3770 45540
rect 3690 45460 3770 45480
rect 3340 45410 3350 45450
rect 3458 45444 3658 45450
rect 3270 45400 3350 45410
rect 2740 44240 2810 45390
rect 2740 43980 2760 44240
rect 2800 43980 2810 44240
rect 3820 45390 3830 45630
rect 3870 45390 3890 45630
rect 3820 44240 3890 45390
rect 3270 44210 3350 44220
rect 2960 44172 3160 44178
rect 2850 44140 2930 44160
rect 2850 44080 2860 44140
rect 2920 44128 2930 44140
rect 2960 44138 2972 44172
rect 3148 44170 3160 44172
rect 3270 44170 3280 44210
rect 3148 44150 3280 44170
rect 3340 44170 3350 44210
rect 3458 44172 3658 44178
rect 3458 44170 3470 44172
rect 3340 44150 3470 44170
rect 3148 44140 3470 44150
rect 3148 44138 3160 44140
rect 2960 44132 3160 44138
rect 3458 44138 3470 44140
rect 3646 44138 3658 44172
rect 3458 44132 3658 44138
rect 3690 44140 3770 44160
rect 2922 44094 2930 44128
rect 2920 44080 2930 44094
rect 2850 44060 2930 44080
rect 2960 44084 3160 44090
rect 2960 44050 2972 44084
rect 3148 44080 3160 44084
rect 3458 44084 3658 44090
rect 3458 44080 3470 44084
rect 3148 44050 3470 44080
rect 3646 44050 3658 44084
rect 3690 44080 3700 44140
rect 3760 44080 3770 44140
rect 3690 44060 3770 44080
rect 2960 44044 3160 44050
rect 2740 43920 2810 43980
rect 2740 43680 2760 43920
rect 2800 43680 2810 43920
rect 3270 44040 3350 44050
rect 3458 44044 3658 44050
rect 3270 43980 3280 44040
rect 3340 43980 3350 44040
rect 3270 43930 3350 43980
rect 3270 43870 3280 43930
rect 3340 43870 3350 43930
rect 2960 43862 3160 43868
rect 2850 43830 2930 43850
rect 2850 43770 2860 43830
rect 2920 43818 2930 43830
rect 2960 43828 2972 43862
rect 3148 43860 3160 43862
rect 3270 43860 3350 43870
rect 3820 44000 3830 44240
rect 3870 44000 3890 44240
rect 3820 43920 3890 44000
rect 3458 43862 3658 43868
rect 3458 43860 3470 43862
rect 3148 43830 3470 43860
rect 3148 43828 3160 43830
rect 2960 43822 3160 43828
rect 3458 43828 3470 43830
rect 3646 43828 3658 43862
rect 3458 43822 3658 43828
rect 3690 43830 3770 43850
rect 2922 43784 2930 43818
rect 2920 43770 2930 43784
rect 2850 43750 2930 43770
rect 2960 43774 3160 43780
rect 2960 43740 2972 43774
rect 3148 43770 3160 43774
rect 3458 43774 3658 43780
rect 3458 43770 3470 43774
rect 3148 43760 3470 43770
rect 3148 43740 3280 43760
rect 2960 43734 3160 43740
rect 3270 43700 3280 43740
rect 3340 43740 3470 43760
rect 3646 43740 3658 43774
rect 3690 43770 3700 43830
rect 3760 43770 3770 43830
rect 3690 43750 3770 43770
rect 3340 43700 3350 43740
rect 3458 43734 3658 43740
rect 3270 43690 3350 43700
rect 2740 42530 2810 43680
rect 2740 42270 2760 42530
rect 2800 42270 2810 42530
rect 3820 43680 3830 43920
rect 3870 43680 3890 43920
rect 3820 42530 3890 43680
rect 3270 42500 3350 42510
rect 2960 42462 3160 42468
rect 2850 42430 2930 42450
rect 2850 42370 2860 42430
rect 2920 42418 2930 42430
rect 2960 42428 2972 42462
rect 3148 42460 3160 42462
rect 3270 42460 3280 42500
rect 3148 42440 3280 42460
rect 3340 42460 3350 42500
rect 3458 42462 3658 42468
rect 3458 42460 3470 42462
rect 3340 42440 3470 42460
rect 3148 42430 3470 42440
rect 3148 42428 3160 42430
rect 2960 42422 3160 42428
rect 3458 42428 3470 42430
rect 3646 42428 3658 42462
rect 3458 42422 3658 42428
rect 3690 42430 3770 42450
rect 2922 42384 2930 42418
rect 2920 42370 2930 42384
rect 2850 42350 2930 42370
rect 2960 42374 3160 42380
rect 2960 42340 2972 42374
rect 3148 42370 3160 42374
rect 3458 42374 3658 42380
rect 3458 42370 3470 42374
rect 3148 42340 3470 42370
rect 3646 42340 3658 42374
rect 3690 42370 3700 42430
rect 3760 42370 3770 42430
rect 3690 42350 3770 42370
rect 2960 42334 3160 42340
rect 2740 42210 2810 42270
rect 2740 41970 2760 42210
rect 2800 41970 2810 42210
rect 3270 42330 3350 42340
rect 3458 42334 3658 42340
rect 3270 42270 3280 42330
rect 3340 42270 3350 42330
rect 3270 42220 3350 42270
rect 3270 42160 3280 42220
rect 3340 42160 3350 42220
rect 2960 42152 3160 42158
rect 2850 42120 2930 42140
rect 2850 42060 2860 42120
rect 2920 42108 2930 42120
rect 2960 42118 2972 42152
rect 3148 42150 3160 42152
rect 3270 42150 3350 42160
rect 3820 42290 3830 42530
rect 3870 42290 3890 42530
rect 3820 42210 3890 42290
rect 3458 42152 3658 42158
rect 3458 42150 3470 42152
rect 3148 42120 3470 42150
rect 3148 42118 3160 42120
rect 2960 42112 3160 42118
rect 3458 42118 3470 42120
rect 3646 42118 3658 42152
rect 3458 42112 3658 42118
rect 3690 42120 3770 42140
rect 2922 42074 2930 42108
rect 2920 42060 2930 42074
rect 2850 42040 2930 42060
rect 2960 42064 3160 42070
rect 2960 42030 2972 42064
rect 3148 42060 3160 42064
rect 3458 42064 3658 42070
rect 3458 42060 3470 42064
rect 3148 42050 3470 42060
rect 3148 42030 3280 42050
rect 2960 42024 3160 42030
rect 3270 41990 3280 42030
rect 3340 42030 3470 42050
rect 3646 42030 3658 42064
rect 3690 42060 3700 42120
rect 3760 42060 3770 42120
rect 3690 42040 3770 42060
rect 3340 41990 3350 42030
rect 3458 42024 3658 42030
rect 3270 41980 3350 41990
rect 2740 40820 2810 41970
rect 2740 40560 2760 40820
rect 2800 40560 2810 40820
rect 3820 41970 3830 42210
rect 3870 41970 3890 42210
rect 3820 40820 3890 41970
rect 3270 40790 3350 40800
rect 2960 40752 3160 40758
rect 2850 40720 2930 40740
rect 2850 40660 2860 40720
rect 2920 40708 2930 40720
rect 2960 40718 2972 40752
rect 3148 40750 3160 40752
rect 3270 40750 3280 40790
rect 3148 40730 3280 40750
rect 3340 40750 3350 40790
rect 3458 40752 3658 40758
rect 3458 40750 3470 40752
rect 3340 40730 3470 40750
rect 3148 40720 3470 40730
rect 3148 40718 3160 40720
rect 2960 40712 3160 40718
rect 3458 40718 3470 40720
rect 3646 40718 3658 40752
rect 3458 40712 3658 40718
rect 3690 40720 3770 40740
rect 2922 40674 2930 40708
rect 2920 40660 2930 40674
rect 2850 40640 2930 40660
rect 2960 40664 3160 40670
rect 2960 40630 2972 40664
rect 3148 40660 3160 40664
rect 3458 40664 3658 40670
rect 3458 40660 3470 40664
rect 3148 40630 3470 40660
rect 3646 40630 3658 40664
rect 3690 40660 3700 40720
rect 3760 40660 3770 40720
rect 3690 40640 3770 40660
rect 2960 40624 3160 40630
rect 2740 40500 2810 40560
rect 2740 40260 2760 40500
rect 2800 40260 2810 40500
rect 3270 40620 3350 40630
rect 3458 40624 3658 40630
rect 3270 40560 3280 40620
rect 3340 40560 3350 40620
rect 3270 40510 3350 40560
rect 3270 40450 3280 40510
rect 3340 40450 3350 40510
rect 2960 40442 3160 40448
rect 2850 40410 2930 40430
rect 2850 40350 2860 40410
rect 2920 40398 2930 40410
rect 2960 40408 2972 40442
rect 3148 40440 3160 40442
rect 3270 40440 3350 40450
rect 3820 40580 3830 40820
rect 3870 40580 3890 40820
rect 3820 40500 3890 40580
rect 3458 40442 3658 40448
rect 3458 40440 3470 40442
rect 3148 40410 3470 40440
rect 3148 40408 3160 40410
rect 2960 40402 3160 40408
rect 3458 40408 3470 40410
rect 3646 40408 3658 40442
rect 3458 40402 3658 40408
rect 3690 40410 3770 40430
rect 2922 40364 2930 40398
rect 2920 40350 2930 40364
rect 2850 40330 2930 40350
rect 2960 40354 3160 40360
rect 2960 40320 2972 40354
rect 3148 40350 3160 40354
rect 3458 40354 3658 40360
rect 3458 40350 3470 40354
rect 3148 40340 3470 40350
rect 3148 40320 3280 40340
rect 2960 40314 3160 40320
rect 3270 40280 3280 40320
rect 3340 40320 3470 40340
rect 3646 40320 3658 40354
rect 3690 40350 3700 40410
rect 3760 40350 3770 40410
rect 3690 40330 3770 40350
rect 3340 40280 3350 40320
rect 3458 40314 3658 40320
rect 3270 40270 3350 40280
rect 2740 39690 2810 40260
rect 3820 40260 3830 40500
rect 3870 40260 3890 40500
rect 3820 39690 3890 40260
rect 2740 39680 2820 39690
rect 2740 39620 2750 39680
rect 2810 39620 2820 39680
rect 3810 39680 3890 39690
rect 3810 39620 3820 39680
rect 3880 39620 3890 39680
rect 3810 39610 3890 39620
rect 3920 66480 3950 67050
rect 3920 66470 3980 66480
rect 3920 66400 3980 66410
rect 3920 64770 3950 66400
rect 4010 65950 4040 67050
rect 3980 65940 4040 65950
rect 3980 65870 4040 65880
rect 3920 64760 3980 64770
rect 3920 64690 3980 64700
rect 3920 63060 3950 64690
rect 4010 64240 4040 65870
rect 3980 64230 4040 64240
rect 3980 64160 4040 64170
rect 3920 63050 3980 63060
rect 3920 62980 3980 62990
rect 3920 61350 3950 62980
rect 4010 62530 4040 64160
rect 3980 62520 4040 62530
rect 3980 62450 4040 62460
rect 3920 61340 3980 61350
rect 3920 61270 3980 61280
rect 3920 59640 3950 61270
rect 4010 60820 4040 62450
rect 3980 60810 4040 60820
rect 3980 60740 4040 60750
rect 3920 59630 3980 59640
rect 3920 59560 3980 59570
rect 3920 57930 3950 59560
rect 4010 59110 4040 60740
rect 3980 59100 4040 59110
rect 3980 59030 4040 59040
rect 3920 57920 3980 57930
rect 3920 57850 3980 57860
rect 3920 56220 3950 57850
rect 4010 57400 4040 59030
rect 3980 57390 4040 57400
rect 3980 57320 4040 57330
rect 3920 56210 3980 56220
rect 3920 56140 3980 56150
rect 3920 54510 3950 56140
rect 4010 55690 4040 57320
rect 3980 55680 4040 55690
rect 3980 55610 4040 55620
rect 3920 54500 3980 54510
rect 3920 54430 3980 54440
rect 3920 52800 3950 54430
rect 4010 53980 4040 55610
rect 3980 53970 4040 53980
rect 3980 53900 4040 53910
rect 3920 52790 3980 52800
rect 3920 52720 3980 52730
rect 3920 51090 3950 52720
rect 4010 52270 4040 53900
rect 3980 52260 4040 52270
rect 3980 52190 4040 52200
rect 3920 51080 3980 51090
rect 3920 51010 3980 51020
rect 3920 49380 3950 51010
rect 4010 50560 4040 52190
rect 3980 50550 4040 50560
rect 3980 50480 4040 50490
rect 3920 49370 3980 49380
rect 3920 49300 3980 49310
rect 3920 47670 3950 49300
rect 4010 48850 4040 50480
rect 3980 48840 4040 48850
rect 3980 48770 4040 48780
rect 3920 47660 3980 47670
rect 3920 47590 3980 47600
rect 3920 45960 3950 47590
rect 4010 47140 4040 48770
rect 3980 47130 4040 47140
rect 3980 47060 4040 47070
rect 3920 45950 3980 45960
rect 3920 45880 3980 45890
rect 3920 44250 3950 45880
rect 4010 45430 4040 47060
rect 3980 45420 4040 45430
rect 3980 45350 4040 45360
rect 3920 44240 3980 44250
rect 3920 44170 3980 44180
rect 3920 42540 3950 44170
rect 4010 43720 4040 45350
rect 3980 43710 4040 43720
rect 3980 43640 4040 43650
rect 3920 42530 3980 42540
rect 3920 42460 3980 42470
rect 3920 40830 3950 42460
rect 4010 42010 4040 43640
rect 3980 42000 4040 42010
rect 3980 41930 4040 41940
rect 3920 40820 3980 40830
rect 3920 40750 3980 40760
rect 2450 39230 2710 39240
rect 2510 39210 2710 39230
rect 2450 39160 2510 39170
rect 3920 38840 3950 40750
rect 4010 40300 4040 41930
rect 3980 40290 4040 40300
rect 3980 40220 4040 40230
rect 4010 39690 4040 40220
rect 3980 39680 4040 39690
rect 3980 39610 4040 39620
rect 4070 66390 4100 67050
rect 4070 66380 4130 66390
rect 4070 66310 4130 66320
rect 4070 64680 4100 66310
rect 4070 64670 4130 64680
rect 4070 64600 4130 64610
rect 4070 62970 4100 64600
rect 4070 62960 4130 62970
rect 4070 62890 4130 62900
rect 4070 61260 4100 62890
rect 4070 61250 4130 61260
rect 4070 61180 4130 61190
rect 4070 59550 4100 61180
rect 4070 59540 4130 59550
rect 4070 59470 4130 59480
rect 4070 57840 4100 59470
rect 4070 57830 4130 57840
rect 4070 57760 4130 57770
rect 4070 56130 4100 57760
rect 4070 56120 4130 56130
rect 4070 56050 4130 56060
rect 4070 54420 4100 56050
rect 4070 54410 4130 54420
rect 4070 54340 4130 54350
rect 4070 52710 4100 54340
rect 4070 52700 4130 52710
rect 4070 52630 4130 52640
rect 4070 51000 4100 52630
rect 4070 50990 4130 51000
rect 4070 50920 4130 50930
rect 4070 49290 4100 50920
rect 4070 49280 4130 49290
rect 4070 49210 4130 49220
rect 4070 47580 4100 49210
rect 4070 47570 4130 47580
rect 4070 47500 4130 47510
rect 4070 45870 4100 47500
rect 4070 45860 4130 45870
rect 4070 45790 4130 45800
rect 4070 44160 4100 45790
rect 4070 44150 4130 44160
rect 4070 44080 4130 44090
rect 4070 42450 4100 44080
rect 4070 42440 4130 42450
rect 4070 42370 4130 42380
rect 4070 40740 4100 42370
rect 4070 40730 4130 40740
rect 4070 40660 4130 40670
rect 4070 39240 4100 40660
rect 4190 39690 4220 67050
rect 4310 39690 4340 67050
rect 4430 39690 4460 67050
rect 4550 39690 4580 67050
rect 4670 39690 4700 67050
rect 4790 39690 4820 67050
rect 6950 39690 6980 67050
rect 7070 39690 7100 67050
rect 7190 39690 7220 67050
rect 7310 39690 7340 67050
rect 7430 39690 7460 67050
rect 7550 39690 7580 67050
rect 7670 66390 7700 67050
rect 7640 66380 7700 66390
rect 7640 66310 7700 66320
rect 7670 64680 7700 66310
rect 7640 64670 7700 64680
rect 7640 64600 7700 64610
rect 7670 62970 7700 64600
rect 7640 62960 7700 62970
rect 7640 62890 7700 62900
rect 7670 61260 7700 62890
rect 7640 61250 7700 61260
rect 7640 61180 7700 61190
rect 7670 59550 7700 61180
rect 7640 59540 7700 59550
rect 7640 59470 7700 59480
rect 7670 57840 7700 59470
rect 7640 57830 7700 57840
rect 7640 57760 7700 57770
rect 7670 56130 7700 57760
rect 7640 56120 7700 56130
rect 7640 56050 7700 56060
rect 7670 54420 7700 56050
rect 7640 54410 7700 54420
rect 7640 54340 7700 54350
rect 7670 52710 7700 54340
rect 7640 52700 7700 52710
rect 7640 52630 7700 52640
rect 7670 51000 7700 52630
rect 7640 50990 7700 51000
rect 7640 50920 7700 50930
rect 7670 49290 7700 50920
rect 7640 49280 7700 49290
rect 7640 49210 7700 49220
rect 7670 47580 7700 49210
rect 7640 47570 7700 47580
rect 7640 47500 7700 47510
rect 7670 45870 7700 47500
rect 7640 45860 7700 45870
rect 7640 45790 7700 45800
rect 7670 44160 7700 45790
rect 7640 44150 7700 44160
rect 7640 44080 7700 44090
rect 7670 42450 7700 44080
rect 7640 42440 7700 42450
rect 7640 42370 7700 42380
rect 7670 40740 7700 42370
rect 7640 40730 7700 40740
rect 7640 40660 7700 40670
rect 7670 39240 7700 40660
rect 7730 66470 7800 67050
rect 7730 66210 7750 66470
rect 7790 66210 7800 66470
rect 8810 66470 8880 67050
rect 8260 66440 8340 66450
rect 7950 66402 8150 66408
rect 7840 66370 7920 66390
rect 7840 66310 7850 66370
rect 7910 66358 7920 66370
rect 7950 66368 7962 66402
rect 8138 66400 8150 66402
rect 8260 66400 8270 66440
rect 8138 66380 8270 66400
rect 8330 66400 8340 66440
rect 8448 66402 8648 66408
rect 8448 66400 8460 66402
rect 8330 66380 8460 66400
rect 8138 66370 8460 66380
rect 8138 66368 8150 66370
rect 7950 66362 8150 66368
rect 8448 66368 8460 66370
rect 8636 66368 8648 66402
rect 8448 66362 8648 66368
rect 8680 66370 8760 66390
rect 7912 66324 7920 66358
rect 7910 66310 7920 66324
rect 7840 66290 7920 66310
rect 7950 66314 8150 66320
rect 7950 66280 7962 66314
rect 8138 66310 8150 66314
rect 8448 66314 8648 66320
rect 8448 66310 8460 66314
rect 8138 66280 8460 66310
rect 8636 66280 8648 66314
rect 8680 66310 8690 66370
rect 8750 66310 8760 66370
rect 8680 66290 8760 66310
rect 7950 66274 8150 66280
rect 7730 66150 7800 66210
rect 7730 65910 7750 66150
rect 7790 65910 7800 66150
rect 8260 66270 8340 66280
rect 8448 66274 8648 66280
rect 8260 66210 8270 66270
rect 8330 66210 8340 66270
rect 8260 66160 8340 66210
rect 8260 66100 8270 66160
rect 8330 66100 8340 66160
rect 7950 66092 8150 66098
rect 7840 66060 7920 66080
rect 7840 66000 7850 66060
rect 7910 66048 7920 66060
rect 7950 66058 7962 66092
rect 8138 66090 8150 66092
rect 8260 66090 8340 66100
rect 8810 66230 8820 66470
rect 8860 66230 8880 66470
rect 8810 66150 8880 66230
rect 8448 66092 8648 66098
rect 8448 66090 8460 66092
rect 8138 66060 8460 66090
rect 8138 66058 8150 66060
rect 7950 66052 8150 66058
rect 8448 66058 8460 66060
rect 8636 66058 8648 66092
rect 8448 66052 8648 66058
rect 8680 66060 8760 66080
rect 7912 66014 7920 66048
rect 7910 66000 7920 66014
rect 7840 65980 7920 66000
rect 7950 66004 8150 66010
rect 7950 65970 7962 66004
rect 8138 66000 8150 66004
rect 8448 66004 8648 66010
rect 8448 66000 8460 66004
rect 8138 65990 8460 66000
rect 8138 65970 8270 65990
rect 7950 65964 8150 65970
rect 8260 65930 8270 65970
rect 8330 65970 8460 65990
rect 8636 65970 8648 66004
rect 8680 66000 8690 66060
rect 8750 66000 8760 66060
rect 8680 65980 8760 66000
rect 8330 65930 8340 65970
rect 8448 65964 8648 65970
rect 8260 65920 8340 65930
rect 7730 64760 7800 65910
rect 7730 64500 7750 64760
rect 7790 64500 7800 64760
rect 8810 65910 8820 66150
rect 8860 65910 8880 66150
rect 8810 64760 8880 65910
rect 8260 64730 8340 64740
rect 7950 64692 8150 64698
rect 7840 64660 7920 64680
rect 7840 64600 7850 64660
rect 7910 64648 7920 64660
rect 7950 64658 7962 64692
rect 8138 64690 8150 64692
rect 8260 64690 8270 64730
rect 8138 64670 8270 64690
rect 8330 64690 8340 64730
rect 8448 64692 8648 64698
rect 8448 64690 8460 64692
rect 8330 64670 8460 64690
rect 8138 64660 8460 64670
rect 8138 64658 8150 64660
rect 7950 64652 8150 64658
rect 8448 64658 8460 64660
rect 8636 64658 8648 64692
rect 8448 64652 8648 64658
rect 8680 64660 8760 64680
rect 7912 64614 7920 64648
rect 7910 64600 7920 64614
rect 7840 64580 7920 64600
rect 7950 64604 8150 64610
rect 7950 64570 7962 64604
rect 8138 64600 8150 64604
rect 8448 64604 8648 64610
rect 8448 64600 8460 64604
rect 8138 64570 8460 64600
rect 8636 64570 8648 64604
rect 8680 64600 8690 64660
rect 8750 64600 8760 64660
rect 8680 64580 8760 64600
rect 7950 64564 8150 64570
rect 7730 64440 7800 64500
rect 7730 64200 7750 64440
rect 7790 64200 7800 64440
rect 8260 64560 8340 64570
rect 8448 64564 8648 64570
rect 8260 64500 8270 64560
rect 8330 64500 8340 64560
rect 8260 64450 8340 64500
rect 8260 64390 8270 64450
rect 8330 64390 8340 64450
rect 7950 64382 8150 64388
rect 7840 64350 7920 64370
rect 7840 64290 7850 64350
rect 7910 64338 7920 64350
rect 7950 64348 7962 64382
rect 8138 64380 8150 64382
rect 8260 64380 8340 64390
rect 8810 64520 8820 64760
rect 8860 64520 8880 64760
rect 8810 64440 8880 64520
rect 8448 64382 8648 64388
rect 8448 64380 8460 64382
rect 8138 64350 8460 64380
rect 8138 64348 8150 64350
rect 7950 64342 8150 64348
rect 8448 64348 8460 64350
rect 8636 64348 8648 64382
rect 8448 64342 8648 64348
rect 8680 64350 8760 64370
rect 7912 64304 7920 64338
rect 7910 64290 7920 64304
rect 7840 64270 7920 64290
rect 7950 64294 8150 64300
rect 7950 64260 7962 64294
rect 8138 64290 8150 64294
rect 8448 64294 8648 64300
rect 8448 64290 8460 64294
rect 8138 64280 8460 64290
rect 8138 64260 8270 64280
rect 7950 64254 8150 64260
rect 8260 64220 8270 64260
rect 8330 64260 8460 64280
rect 8636 64260 8648 64294
rect 8680 64290 8690 64350
rect 8750 64290 8760 64350
rect 8680 64270 8760 64290
rect 8330 64220 8340 64260
rect 8448 64254 8648 64260
rect 8260 64210 8340 64220
rect 7730 63050 7800 64200
rect 7730 62790 7750 63050
rect 7790 62790 7800 63050
rect 8810 64200 8820 64440
rect 8860 64200 8880 64440
rect 8810 63050 8880 64200
rect 8260 63020 8340 63030
rect 7950 62982 8150 62988
rect 7840 62950 7920 62970
rect 7840 62890 7850 62950
rect 7910 62938 7920 62950
rect 7950 62948 7962 62982
rect 8138 62980 8150 62982
rect 8260 62980 8270 63020
rect 8138 62960 8270 62980
rect 8330 62980 8340 63020
rect 8448 62982 8648 62988
rect 8448 62980 8460 62982
rect 8330 62960 8460 62980
rect 8138 62950 8460 62960
rect 8138 62948 8150 62950
rect 7950 62942 8150 62948
rect 8448 62948 8460 62950
rect 8636 62948 8648 62982
rect 8448 62942 8648 62948
rect 8680 62950 8760 62970
rect 7912 62904 7920 62938
rect 7910 62890 7920 62904
rect 7840 62870 7920 62890
rect 7950 62894 8150 62900
rect 7950 62860 7962 62894
rect 8138 62890 8150 62894
rect 8448 62894 8648 62900
rect 8448 62890 8460 62894
rect 8138 62860 8460 62890
rect 8636 62860 8648 62894
rect 8680 62890 8690 62950
rect 8750 62890 8760 62950
rect 8680 62870 8760 62890
rect 7950 62854 8150 62860
rect 7730 62730 7800 62790
rect 7730 62490 7750 62730
rect 7790 62490 7800 62730
rect 8260 62850 8340 62860
rect 8448 62854 8648 62860
rect 8260 62790 8270 62850
rect 8330 62790 8340 62850
rect 8260 62740 8340 62790
rect 8260 62680 8270 62740
rect 8330 62680 8340 62740
rect 7950 62672 8150 62678
rect 7840 62640 7920 62660
rect 7840 62580 7850 62640
rect 7910 62628 7920 62640
rect 7950 62638 7962 62672
rect 8138 62670 8150 62672
rect 8260 62670 8340 62680
rect 8810 62810 8820 63050
rect 8860 62810 8880 63050
rect 8810 62730 8880 62810
rect 8448 62672 8648 62678
rect 8448 62670 8460 62672
rect 8138 62640 8460 62670
rect 8138 62638 8150 62640
rect 7950 62632 8150 62638
rect 8448 62638 8460 62640
rect 8636 62638 8648 62672
rect 8448 62632 8648 62638
rect 8680 62640 8760 62660
rect 7912 62594 7920 62628
rect 7910 62580 7920 62594
rect 7840 62560 7920 62580
rect 7950 62584 8150 62590
rect 7950 62550 7962 62584
rect 8138 62580 8150 62584
rect 8448 62584 8648 62590
rect 8448 62580 8460 62584
rect 8138 62570 8460 62580
rect 8138 62550 8270 62570
rect 7950 62544 8150 62550
rect 8260 62510 8270 62550
rect 8330 62550 8460 62570
rect 8636 62550 8648 62584
rect 8680 62580 8690 62640
rect 8750 62580 8760 62640
rect 8680 62560 8760 62580
rect 8330 62510 8340 62550
rect 8448 62544 8648 62550
rect 8260 62500 8340 62510
rect 7730 61340 7800 62490
rect 7730 61080 7750 61340
rect 7790 61080 7800 61340
rect 8810 62490 8820 62730
rect 8860 62490 8880 62730
rect 8810 61340 8880 62490
rect 8260 61310 8340 61320
rect 7950 61272 8150 61278
rect 7840 61240 7920 61260
rect 7840 61180 7850 61240
rect 7910 61228 7920 61240
rect 7950 61238 7962 61272
rect 8138 61270 8150 61272
rect 8260 61270 8270 61310
rect 8138 61250 8270 61270
rect 8330 61270 8340 61310
rect 8448 61272 8648 61278
rect 8448 61270 8460 61272
rect 8330 61250 8460 61270
rect 8138 61240 8460 61250
rect 8138 61238 8150 61240
rect 7950 61232 8150 61238
rect 8448 61238 8460 61240
rect 8636 61238 8648 61272
rect 8448 61232 8648 61238
rect 8680 61240 8760 61260
rect 7912 61194 7920 61228
rect 7910 61180 7920 61194
rect 7840 61160 7920 61180
rect 7950 61184 8150 61190
rect 7950 61150 7962 61184
rect 8138 61180 8150 61184
rect 8448 61184 8648 61190
rect 8448 61180 8460 61184
rect 8138 61150 8460 61180
rect 8636 61150 8648 61184
rect 8680 61180 8690 61240
rect 8750 61180 8760 61240
rect 8680 61160 8760 61180
rect 7950 61144 8150 61150
rect 7730 61020 7800 61080
rect 7730 60780 7750 61020
rect 7790 60780 7800 61020
rect 8260 61140 8340 61150
rect 8448 61144 8648 61150
rect 8260 61080 8270 61140
rect 8330 61080 8340 61140
rect 8260 61030 8340 61080
rect 8260 60970 8270 61030
rect 8330 60970 8340 61030
rect 7950 60962 8150 60968
rect 7840 60930 7920 60950
rect 7840 60870 7850 60930
rect 7910 60918 7920 60930
rect 7950 60928 7962 60962
rect 8138 60960 8150 60962
rect 8260 60960 8340 60970
rect 8810 61100 8820 61340
rect 8860 61100 8880 61340
rect 8810 61020 8880 61100
rect 8448 60962 8648 60968
rect 8448 60960 8460 60962
rect 8138 60930 8460 60960
rect 8138 60928 8150 60930
rect 7950 60922 8150 60928
rect 8448 60928 8460 60930
rect 8636 60928 8648 60962
rect 8448 60922 8648 60928
rect 8680 60930 8760 60950
rect 7912 60884 7920 60918
rect 7910 60870 7920 60884
rect 7840 60850 7920 60870
rect 7950 60874 8150 60880
rect 7950 60840 7962 60874
rect 8138 60870 8150 60874
rect 8448 60874 8648 60880
rect 8448 60870 8460 60874
rect 8138 60860 8460 60870
rect 8138 60840 8270 60860
rect 7950 60834 8150 60840
rect 8260 60800 8270 60840
rect 8330 60840 8460 60860
rect 8636 60840 8648 60874
rect 8680 60870 8690 60930
rect 8750 60870 8760 60930
rect 8680 60850 8760 60870
rect 8330 60800 8340 60840
rect 8448 60834 8648 60840
rect 8260 60790 8340 60800
rect 7730 59630 7800 60780
rect 7730 59370 7750 59630
rect 7790 59370 7800 59630
rect 8810 60780 8820 61020
rect 8860 60780 8880 61020
rect 8810 59630 8880 60780
rect 8260 59600 8340 59610
rect 7950 59562 8150 59568
rect 7840 59530 7920 59550
rect 7840 59470 7850 59530
rect 7910 59518 7920 59530
rect 7950 59528 7962 59562
rect 8138 59560 8150 59562
rect 8260 59560 8270 59600
rect 8138 59540 8270 59560
rect 8330 59560 8340 59600
rect 8448 59562 8648 59568
rect 8448 59560 8460 59562
rect 8330 59540 8460 59560
rect 8138 59530 8460 59540
rect 8138 59528 8150 59530
rect 7950 59522 8150 59528
rect 8448 59528 8460 59530
rect 8636 59528 8648 59562
rect 8448 59522 8648 59528
rect 8680 59530 8760 59550
rect 7912 59484 7920 59518
rect 7910 59470 7920 59484
rect 7840 59450 7920 59470
rect 7950 59474 8150 59480
rect 7950 59440 7962 59474
rect 8138 59470 8150 59474
rect 8448 59474 8648 59480
rect 8448 59470 8460 59474
rect 8138 59440 8460 59470
rect 8636 59440 8648 59474
rect 8680 59470 8690 59530
rect 8750 59470 8760 59530
rect 8680 59450 8760 59470
rect 7950 59434 8150 59440
rect 7730 59310 7800 59370
rect 7730 59070 7750 59310
rect 7790 59070 7800 59310
rect 8260 59430 8340 59440
rect 8448 59434 8648 59440
rect 8260 59370 8270 59430
rect 8330 59370 8340 59430
rect 8260 59320 8340 59370
rect 8260 59260 8270 59320
rect 8330 59260 8340 59320
rect 7950 59252 8150 59258
rect 7840 59220 7920 59240
rect 7840 59160 7850 59220
rect 7910 59208 7920 59220
rect 7950 59218 7962 59252
rect 8138 59250 8150 59252
rect 8260 59250 8340 59260
rect 8810 59390 8820 59630
rect 8860 59390 8880 59630
rect 8810 59310 8880 59390
rect 8448 59252 8648 59258
rect 8448 59250 8460 59252
rect 8138 59220 8460 59250
rect 8138 59218 8150 59220
rect 7950 59212 8150 59218
rect 8448 59218 8460 59220
rect 8636 59218 8648 59252
rect 8448 59212 8648 59218
rect 8680 59220 8760 59240
rect 7912 59174 7920 59208
rect 7910 59160 7920 59174
rect 7840 59140 7920 59160
rect 7950 59164 8150 59170
rect 7950 59130 7962 59164
rect 8138 59160 8150 59164
rect 8448 59164 8648 59170
rect 8448 59160 8460 59164
rect 8138 59150 8460 59160
rect 8138 59130 8270 59150
rect 7950 59124 8150 59130
rect 8260 59090 8270 59130
rect 8330 59130 8460 59150
rect 8636 59130 8648 59164
rect 8680 59160 8690 59220
rect 8750 59160 8760 59220
rect 8680 59140 8760 59160
rect 8330 59090 8340 59130
rect 8448 59124 8648 59130
rect 8260 59080 8340 59090
rect 7730 57920 7800 59070
rect 7730 57660 7750 57920
rect 7790 57660 7800 57920
rect 8810 59070 8820 59310
rect 8860 59070 8880 59310
rect 8810 57920 8880 59070
rect 8260 57890 8340 57900
rect 7950 57852 8150 57858
rect 7840 57820 7920 57840
rect 7840 57760 7850 57820
rect 7910 57808 7920 57820
rect 7950 57818 7962 57852
rect 8138 57850 8150 57852
rect 8260 57850 8270 57890
rect 8138 57830 8270 57850
rect 8330 57850 8340 57890
rect 8448 57852 8648 57858
rect 8448 57850 8460 57852
rect 8330 57830 8460 57850
rect 8138 57820 8460 57830
rect 8138 57818 8150 57820
rect 7950 57812 8150 57818
rect 8448 57818 8460 57820
rect 8636 57818 8648 57852
rect 8448 57812 8648 57818
rect 8680 57820 8760 57840
rect 7912 57774 7920 57808
rect 7910 57760 7920 57774
rect 7840 57740 7920 57760
rect 7950 57764 8150 57770
rect 7950 57730 7962 57764
rect 8138 57760 8150 57764
rect 8448 57764 8648 57770
rect 8448 57760 8460 57764
rect 8138 57730 8460 57760
rect 8636 57730 8648 57764
rect 8680 57760 8690 57820
rect 8750 57760 8760 57820
rect 8680 57740 8760 57760
rect 7950 57724 8150 57730
rect 7730 57600 7800 57660
rect 7730 57360 7750 57600
rect 7790 57360 7800 57600
rect 8260 57720 8340 57730
rect 8448 57724 8648 57730
rect 8260 57660 8270 57720
rect 8330 57660 8340 57720
rect 8260 57610 8340 57660
rect 8260 57550 8270 57610
rect 8330 57550 8340 57610
rect 7950 57542 8150 57548
rect 7840 57510 7920 57530
rect 7840 57450 7850 57510
rect 7910 57498 7920 57510
rect 7950 57508 7962 57542
rect 8138 57540 8150 57542
rect 8260 57540 8340 57550
rect 8810 57680 8820 57920
rect 8860 57680 8880 57920
rect 8810 57600 8880 57680
rect 8448 57542 8648 57548
rect 8448 57540 8460 57542
rect 8138 57510 8460 57540
rect 8138 57508 8150 57510
rect 7950 57502 8150 57508
rect 8448 57508 8460 57510
rect 8636 57508 8648 57542
rect 8448 57502 8648 57508
rect 8680 57510 8760 57530
rect 7912 57464 7920 57498
rect 7910 57450 7920 57464
rect 7840 57430 7920 57450
rect 7950 57454 8150 57460
rect 7950 57420 7962 57454
rect 8138 57450 8150 57454
rect 8448 57454 8648 57460
rect 8448 57450 8460 57454
rect 8138 57440 8460 57450
rect 8138 57420 8270 57440
rect 7950 57414 8150 57420
rect 8260 57380 8270 57420
rect 8330 57420 8460 57440
rect 8636 57420 8648 57454
rect 8680 57450 8690 57510
rect 8750 57450 8760 57510
rect 8680 57430 8760 57450
rect 8330 57380 8340 57420
rect 8448 57414 8648 57420
rect 8260 57370 8340 57380
rect 7730 56210 7800 57360
rect 7730 55950 7750 56210
rect 7790 55950 7800 56210
rect 8810 57360 8820 57600
rect 8860 57360 8880 57600
rect 8810 56210 8880 57360
rect 8260 56180 8340 56190
rect 7950 56142 8150 56148
rect 7840 56110 7920 56130
rect 7840 56050 7850 56110
rect 7910 56098 7920 56110
rect 7950 56108 7962 56142
rect 8138 56140 8150 56142
rect 8260 56140 8270 56180
rect 8138 56120 8270 56140
rect 8330 56140 8340 56180
rect 8448 56142 8648 56148
rect 8448 56140 8460 56142
rect 8330 56120 8460 56140
rect 8138 56110 8460 56120
rect 8138 56108 8150 56110
rect 7950 56102 8150 56108
rect 8448 56108 8460 56110
rect 8636 56108 8648 56142
rect 8448 56102 8648 56108
rect 8680 56110 8760 56130
rect 7912 56064 7920 56098
rect 7910 56050 7920 56064
rect 7840 56030 7920 56050
rect 7950 56054 8150 56060
rect 7950 56020 7962 56054
rect 8138 56050 8150 56054
rect 8448 56054 8648 56060
rect 8448 56050 8460 56054
rect 8138 56020 8460 56050
rect 8636 56020 8648 56054
rect 8680 56050 8690 56110
rect 8750 56050 8760 56110
rect 8680 56030 8760 56050
rect 7950 56014 8150 56020
rect 7730 55890 7800 55950
rect 7730 55650 7750 55890
rect 7790 55650 7800 55890
rect 8260 56010 8340 56020
rect 8448 56014 8648 56020
rect 8260 55950 8270 56010
rect 8330 55950 8340 56010
rect 8260 55900 8340 55950
rect 8260 55840 8270 55900
rect 8330 55840 8340 55900
rect 7950 55832 8150 55838
rect 7840 55800 7920 55820
rect 7840 55740 7850 55800
rect 7910 55788 7920 55800
rect 7950 55798 7962 55832
rect 8138 55830 8150 55832
rect 8260 55830 8340 55840
rect 8810 55970 8820 56210
rect 8860 55970 8880 56210
rect 8810 55890 8880 55970
rect 8448 55832 8648 55838
rect 8448 55830 8460 55832
rect 8138 55800 8460 55830
rect 8138 55798 8150 55800
rect 7950 55792 8150 55798
rect 8448 55798 8460 55800
rect 8636 55798 8648 55832
rect 8448 55792 8648 55798
rect 8680 55800 8760 55820
rect 7912 55754 7920 55788
rect 7910 55740 7920 55754
rect 7840 55720 7920 55740
rect 7950 55744 8150 55750
rect 7950 55710 7962 55744
rect 8138 55740 8150 55744
rect 8448 55744 8648 55750
rect 8448 55740 8460 55744
rect 8138 55730 8460 55740
rect 8138 55710 8270 55730
rect 7950 55704 8150 55710
rect 8260 55670 8270 55710
rect 8330 55710 8460 55730
rect 8636 55710 8648 55744
rect 8680 55740 8690 55800
rect 8750 55740 8760 55800
rect 8680 55720 8760 55740
rect 8330 55670 8340 55710
rect 8448 55704 8648 55710
rect 8260 55660 8340 55670
rect 7730 54500 7800 55650
rect 7730 54240 7750 54500
rect 7790 54240 7800 54500
rect 8810 55650 8820 55890
rect 8860 55650 8880 55890
rect 8810 54500 8880 55650
rect 8260 54470 8340 54480
rect 7950 54432 8150 54438
rect 7840 54400 7920 54420
rect 7840 54340 7850 54400
rect 7910 54388 7920 54400
rect 7950 54398 7962 54432
rect 8138 54430 8150 54432
rect 8260 54430 8270 54470
rect 8138 54410 8270 54430
rect 8330 54430 8340 54470
rect 8448 54432 8648 54438
rect 8448 54430 8460 54432
rect 8330 54410 8460 54430
rect 8138 54400 8460 54410
rect 8138 54398 8150 54400
rect 7950 54392 8150 54398
rect 8448 54398 8460 54400
rect 8636 54398 8648 54432
rect 8448 54392 8648 54398
rect 8680 54400 8760 54420
rect 7912 54354 7920 54388
rect 7910 54340 7920 54354
rect 7840 54320 7920 54340
rect 7950 54344 8150 54350
rect 7950 54310 7962 54344
rect 8138 54340 8150 54344
rect 8448 54344 8648 54350
rect 8448 54340 8460 54344
rect 8138 54310 8460 54340
rect 8636 54310 8648 54344
rect 8680 54340 8690 54400
rect 8750 54340 8760 54400
rect 8680 54320 8760 54340
rect 7950 54304 8150 54310
rect 7730 54180 7800 54240
rect 7730 53940 7750 54180
rect 7790 53940 7800 54180
rect 8260 54300 8340 54310
rect 8448 54304 8648 54310
rect 8260 54240 8270 54300
rect 8330 54240 8340 54300
rect 8260 54190 8340 54240
rect 8260 54130 8270 54190
rect 8330 54130 8340 54190
rect 7950 54122 8150 54128
rect 7840 54090 7920 54110
rect 7840 54030 7850 54090
rect 7910 54078 7920 54090
rect 7950 54088 7962 54122
rect 8138 54120 8150 54122
rect 8260 54120 8340 54130
rect 8810 54260 8820 54500
rect 8860 54260 8880 54500
rect 8810 54180 8880 54260
rect 8448 54122 8648 54128
rect 8448 54120 8460 54122
rect 8138 54090 8460 54120
rect 8138 54088 8150 54090
rect 7950 54082 8150 54088
rect 8448 54088 8460 54090
rect 8636 54088 8648 54122
rect 8448 54082 8648 54088
rect 8680 54090 8760 54110
rect 7912 54044 7920 54078
rect 7910 54030 7920 54044
rect 7840 54010 7920 54030
rect 7950 54034 8150 54040
rect 7950 54000 7962 54034
rect 8138 54030 8150 54034
rect 8448 54034 8648 54040
rect 8448 54030 8460 54034
rect 8138 54020 8460 54030
rect 8138 54000 8270 54020
rect 7950 53994 8150 54000
rect 8260 53960 8270 54000
rect 8330 54000 8460 54020
rect 8636 54000 8648 54034
rect 8680 54030 8690 54090
rect 8750 54030 8760 54090
rect 8680 54010 8760 54030
rect 8330 53960 8340 54000
rect 8448 53994 8648 54000
rect 8260 53950 8340 53960
rect 7730 52790 7800 53940
rect 7730 52530 7750 52790
rect 7790 52530 7800 52790
rect 8810 53940 8820 54180
rect 8860 53940 8880 54180
rect 8810 52790 8880 53940
rect 8260 52760 8340 52770
rect 7950 52722 8150 52728
rect 7840 52690 7920 52710
rect 7840 52630 7850 52690
rect 7910 52678 7920 52690
rect 7950 52688 7962 52722
rect 8138 52720 8150 52722
rect 8260 52720 8270 52760
rect 8138 52700 8270 52720
rect 8330 52720 8340 52760
rect 8448 52722 8648 52728
rect 8448 52720 8460 52722
rect 8330 52700 8460 52720
rect 8138 52690 8460 52700
rect 8138 52688 8150 52690
rect 7950 52682 8150 52688
rect 8448 52688 8460 52690
rect 8636 52688 8648 52722
rect 8448 52682 8648 52688
rect 8680 52690 8760 52710
rect 7912 52644 7920 52678
rect 7910 52630 7920 52644
rect 7840 52610 7920 52630
rect 7950 52634 8150 52640
rect 7950 52600 7962 52634
rect 8138 52630 8150 52634
rect 8448 52634 8648 52640
rect 8448 52630 8460 52634
rect 8138 52600 8460 52630
rect 8636 52600 8648 52634
rect 8680 52630 8690 52690
rect 8750 52630 8760 52690
rect 8680 52610 8760 52630
rect 7950 52594 8150 52600
rect 7730 52470 7800 52530
rect 7730 52230 7750 52470
rect 7790 52230 7800 52470
rect 8260 52590 8340 52600
rect 8448 52594 8648 52600
rect 8260 52530 8270 52590
rect 8330 52530 8340 52590
rect 8260 52480 8340 52530
rect 8260 52420 8270 52480
rect 8330 52420 8340 52480
rect 7950 52412 8150 52418
rect 7840 52380 7920 52400
rect 7840 52320 7850 52380
rect 7910 52368 7920 52380
rect 7950 52378 7962 52412
rect 8138 52410 8150 52412
rect 8260 52410 8340 52420
rect 8810 52550 8820 52790
rect 8860 52550 8880 52790
rect 8810 52470 8880 52550
rect 8448 52412 8648 52418
rect 8448 52410 8460 52412
rect 8138 52380 8460 52410
rect 8138 52378 8150 52380
rect 7950 52372 8150 52378
rect 8448 52378 8460 52380
rect 8636 52378 8648 52412
rect 8448 52372 8648 52378
rect 8680 52380 8760 52400
rect 7912 52334 7920 52368
rect 7910 52320 7920 52334
rect 7840 52300 7920 52320
rect 7950 52324 8150 52330
rect 7950 52290 7962 52324
rect 8138 52320 8150 52324
rect 8448 52324 8648 52330
rect 8448 52320 8460 52324
rect 8138 52310 8460 52320
rect 8138 52290 8270 52310
rect 7950 52284 8150 52290
rect 8260 52250 8270 52290
rect 8330 52290 8460 52310
rect 8636 52290 8648 52324
rect 8680 52320 8690 52380
rect 8750 52320 8760 52380
rect 8680 52300 8760 52320
rect 8330 52250 8340 52290
rect 8448 52284 8648 52290
rect 8260 52240 8340 52250
rect 7730 51080 7800 52230
rect 7730 50820 7750 51080
rect 7790 50820 7800 51080
rect 8810 52230 8820 52470
rect 8860 52230 8880 52470
rect 8810 51080 8880 52230
rect 8260 51050 8340 51060
rect 7950 51012 8150 51018
rect 7840 50980 7920 51000
rect 7840 50920 7850 50980
rect 7910 50968 7920 50980
rect 7950 50978 7962 51012
rect 8138 51010 8150 51012
rect 8260 51010 8270 51050
rect 8138 50990 8270 51010
rect 8330 51010 8340 51050
rect 8448 51012 8648 51018
rect 8448 51010 8460 51012
rect 8330 50990 8460 51010
rect 8138 50980 8460 50990
rect 8138 50978 8150 50980
rect 7950 50972 8150 50978
rect 8448 50978 8460 50980
rect 8636 50978 8648 51012
rect 8448 50972 8648 50978
rect 8680 50980 8760 51000
rect 7912 50934 7920 50968
rect 7910 50920 7920 50934
rect 7840 50900 7920 50920
rect 7950 50924 8150 50930
rect 7950 50890 7962 50924
rect 8138 50920 8150 50924
rect 8448 50924 8648 50930
rect 8448 50920 8460 50924
rect 8138 50890 8460 50920
rect 8636 50890 8648 50924
rect 8680 50920 8690 50980
rect 8750 50920 8760 50980
rect 8680 50900 8760 50920
rect 7950 50884 8150 50890
rect 7730 50760 7800 50820
rect 7730 50520 7750 50760
rect 7790 50520 7800 50760
rect 8260 50880 8340 50890
rect 8448 50884 8648 50890
rect 8260 50820 8270 50880
rect 8330 50820 8340 50880
rect 8260 50770 8340 50820
rect 8260 50710 8270 50770
rect 8330 50710 8340 50770
rect 7950 50702 8150 50708
rect 7840 50670 7920 50690
rect 7840 50610 7850 50670
rect 7910 50658 7920 50670
rect 7950 50668 7962 50702
rect 8138 50700 8150 50702
rect 8260 50700 8340 50710
rect 8810 50840 8820 51080
rect 8860 50840 8880 51080
rect 8810 50760 8880 50840
rect 8448 50702 8648 50708
rect 8448 50700 8460 50702
rect 8138 50670 8460 50700
rect 8138 50668 8150 50670
rect 7950 50662 8150 50668
rect 8448 50668 8460 50670
rect 8636 50668 8648 50702
rect 8448 50662 8648 50668
rect 8680 50670 8760 50690
rect 7912 50624 7920 50658
rect 7910 50610 7920 50624
rect 7840 50590 7920 50610
rect 7950 50614 8150 50620
rect 7950 50580 7962 50614
rect 8138 50610 8150 50614
rect 8448 50614 8648 50620
rect 8448 50610 8460 50614
rect 8138 50600 8460 50610
rect 8138 50580 8270 50600
rect 7950 50574 8150 50580
rect 8260 50540 8270 50580
rect 8330 50580 8460 50600
rect 8636 50580 8648 50614
rect 8680 50610 8690 50670
rect 8750 50610 8760 50670
rect 8680 50590 8760 50610
rect 8330 50540 8340 50580
rect 8448 50574 8648 50580
rect 8260 50530 8340 50540
rect 7730 49370 7800 50520
rect 7730 49110 7750 49370
rect 7790 49110 7800 49370
rect 8810 50520 8820 50760
rect 8860 50520 8880 50760
rect 8810 49370 8880 50520
rect 8260 49340 8340 49350
rect 7950 49302 8150 49308
rect 7840 49270 7920 49290
rect 7840 49210 7850 49270
rect 7910 49258 7920 49270
rect 7950 49268 7962 49302
rect 8138 49300 8150 49302
rect 8260 49300 8270 49340
rect 8138 49280 8270 49300
rect 8330 49300 8340 49340
rect 8448 49302 8648 49308
rect 8448 49300 8460 49302
rect 8330 49280 8460 49300
rect 8138 49270 8460 49280
rect 8138 49268 8150 49270
rect 7950 49262 8150 49268
rect 8448 49268 8460 49270
rect 8636 49268 8648 49302
rect 8448 49262 8648 49268
rect 8680 49270 8760 49290
rect 7912 49224 7920 49258
rect 7910 49210 7920 49224
rect 7840 49190 7920 49210
rect 7950 49214 8150 49220
rect 7950 49180 7962 49214
rect 8138 49210 8150 49214
rect 8448 49214 8648 49220
rect 8448 49210 8460 49214
rect 8138 49180 8460 49210
rect 8636 49180 8648 49214
rect 8680 49210 8690 49270
rect 8750 49210 8760 49270
rect 8680 49190 8760 49210
rect 7950 49174 8150 49180
rect 7730 49050 7800 49110
rect 7730 48810 7750 49050
rect 7790 48810 7800 49050
rect 8260 49170 8340 49180
rect 8448 49174 8648 49180
rect 8260 49110 8270 49170
rect 8330 49110 8340 49170
rect 8260 49060 8340 49110
rect 8260 49000 8270 49060
rect 8330 49000 8340 49060
rect 7950 48992 8150 48998
rect 7840 48960 7920 48980
rect 7840 48900 7850 48960
rect 7910 48948 7920 48960
rect 7950 48958 7962 48992
rect 8138 48990 8150 48992
rect 8260 48990 8340 49000
rect 8810 49130 8820 49370
rect 8860 49130 8880 49370
rect 8810 49050 8880 49130
rect 8448 48992 8648 48998
rect 8448 48990 8460 48992
rect 8138 48960 8460 48990
rect 8138 48958 8150 48960
rect 7950 48952 8150 48958
rect 8448 48958 8460 48960
rect 8636 48958 8648 48992
rect 8448 48952 8648 48958
rect 8680 48960 8760 48980
rect 7912 48914 7920 48948
rect 7910 48900 7920 48914
rect 7840 48880 7920 48900
rect 7950 48904 8150 48910
rect 7950 48870 7962 48904
rect 8138 48900 8150 48904
rect 8448 48904 8648 48910
rect 8448 48900 8460 48904
rect 8138 48890 8460 48900
rect 8138 48870 8270 48890
rect 7950 48864 8150 48870
rect 8260 48830 8270 48870
rect 8330 48870 8460 48890
rect 8636 48870 8648 48904
rect 8680 48900 8690 48960
rect 8750 48900 8760 48960
rect 8680 48880 8760 48900
rect 8330 48830 8340 48870
rect 8448 48864 8648 48870
rect 8260 48820 8340 48830
rect 7730 47660 7800 48810
rect 7730 47400 7750 47660
rect 7790 47400 7800 47660
rect 8810 48810 8820 49050
rect 8860 48810 8880 49050
rect 8810 47660 8880 48810
rect 8260 47630 8340 47640
rect 7950 47592 8150 47598
rect 7840 47560 7920 47580
rect 7840 47500 7850 47560
rect 7910 47548 7920 47560
rect 7950 47558 7962 47592
rect 8138 47590 8150 47592
rect 8260 47590 8270 47630
rect 8138 47570 8270 47590
rect 8330 47590 8340 47630
rect 8448 47592 8648 47598
rect 8448 47590 8460 47592
rect 8330 47570 8460 47590
rect 8138 47560 8460 47570
rect 8138 47558 8150 47560
rect 7950 47552 8150 47558
rect 8448 47558 8460 47560
rect 8636 47558 8648 47592
rect 8448 47552 8648 47558
rect 8680 47560 8760 47580
rect 7912 47514 7920 47548
rect 7910 47500 7920 47514
rect 7840 47480 7920 47500
rect 7950 47504 8150 47510
rect 7950 47470 7962 47504
rect 8138 47500 8150 47504
rect 8448 47504 8648 47510
rect 8448 47500 8460 47504
rect 8138 47470 8460 47500
rect 8636 47470 8648 47504
rect 8680 47500 8690 47560
rect 8750 47500 8760 47560
rect 8680 47480 8760 47500
rect 7950 47464 8150 47470
rect 7730 47340 7800 47400
rect 7730 47100 7750 47340
rect 7790 47100 7800 47340
rect 8260 47460 8340 47470
rect 8448 47464 8648 47470
rect 8260 47400 8270 47460
rect 8330 47400 8340 47460
rect 8260 47350 8340 47400
rect 8260 47290 8270 47350
rect 8330 47290 8340 47350
rect 7950 47282 8150 47288
rect 7840 47250 7920 47270
rect 7840 47190 7850 47250
rect 7910 47238 7920 47250
rect 7950 47248 7962 47282
rect 8138 47280 8150 47282
rect 8260 47280 8340 47290
rect 8810 47420 8820 47660
rect 8860 47420 8880 47660
rect 8810 47340 8880 47420
rect 8448 47282 8648 47288
rect 8448 47280 8460 47282
rect 8138 47250 8460 47280
rect 8138 47248 8150 47250
rect 7950 47242 8150 47248
rect 8448 47248 8460 47250
rect 8636 47248 8648 47282
rect 8448 47242 8648 47248
rect 8680 47250 8760 47270
rect 7912 47204 7920 47238
rect 7910 47190 7920 47204
rect 7840 47170 7920 47190
rect 7950 47194 8150 47200
rect 7950 47160 7962 47194
rect 8138 47190 8150 47194
rect 8448 47194 8648 47200
rect 8448 47190 8460 47194
rect 8138 47180 8460 47190
rect 8138 47160 8270 47180
rect 7950 47154 8150 47160
rect 8260 47120 8270 47160
rect 8330 47160 8460 47180
rect 8636 47160 8648 47194
rect 8680 47190 8690 47250
rect 8750 47190 8760 47250
rect 8680 47170 8760 47190
rect 8330 47120 8340 47160
rect 8448 47154 8648 47160
rect 8260 47110 8340 47120
rect 7730 45950 7800 47100
rect 7730 45690 7750 45950
rect 7790 45690 7800 45950
rect 8810 47100 8820 47340
rect 8860 47100 8880 47340
rect 8810 45950 8880 47100
rect 8260 45920 8340 45930
rect 7950 45882 8150 45888
rect 7840 45850 7920 45870
rect 7840 45790 7850 45850
rect 7910 45838 7920 45850
rect 7950 45848 7962 45882
rect 8138 45880 8150 45882
rect 8260 45880 8270 45920
rect 8138 45860 8270 45880
rect 8330 45880 8340 45920
rect 8448 45882 8648 45888
rect 8448 45880 8460 45882
rect 8330 45860 8460 45880
rect 8138 45850 8460 45860
rect 8138 45848 8150 45850
rect 7950 45842 8150 45848
rect 8448 45848 8460 45850
rect 8636 45848 8648 45882
rect 8448 45842 8648 45848
rect 8680 45850 8760 45870
rect 7912 45804 7920 45838
rect 7910 45790 7920 45804
rect 7840 45770 7920 45790
rect 7950 45794 8150 45800
rect 7950 45760 7962 45794
rect 8138 45790 8150 45794
rect 8448 45794 8648 45800
rect 8448 45790 8460 45794
rect 8138 45760 8460 45790
rect 8636 45760 8648 45794
rect 8680 45790 8690 45850
rect 8750 45790 8760 45850
rect 8680 45770 8760 45790
rect 7950 45754 8150 45760
rect 7730 45630 7800 45690
rect 7730 45390 7750 45630
rect 7790 45390 7800 45630
rect 8260 45750 8340 45760
rect 8448 45754 8648 45760
rect 8260 45690 8270 45750
rect 8330 45690 8340 45750
rect 8260 45640 8340 45690
rect 8260 45580 8270 45640
rect 8330 45580 8340 45640
rect 7950 45572 8150 45578
rect 7840 45540 7920 45560
rect 7840 45480 7850 45540
rect 7910 45528 7920 45540
rect 7950 45538 7962 45572
rect 8138 45570 8150 45572
rect 8260 45570 8340 45580
rect 8810 45710 8820 45950
rect 8860 45710 8880 45950
rect 8810 45630 8880 45710
rect 8448 45572 8648 45578
rect 8448 45570 8460 45572
rect 8138 45540 8460 45570
rect 8138 45538 8150 45540
rect 7950 45532 8150 45538
rect 8448 45538 8460 45540
rect 8636 45538 8648 45572
rect 8448 45532 8648 45538
rect 8680 45540 8760 45560
rect 7912 45494 7920 45528
rect 7910 45480 7920 45494
rect 7840 45460 7920 45480
rect 7950 45484 8150 45490
rect 7950 45450 7962 45484
rect 8138 45480 8150 45484
rect 8448 45484 8648 45490
rect 8448 45480 8460 45484
rect 8138 45470 8460 45480
rect 8138 45450 8270 45470
rect 7950 45444 8150 45450
rect 8260 45410 8270 45450
rect 8330 45450 8460 45470
rect 8636 45450 8648 45484
rect 8680 45480 8690 45540
rect 8750 45480 8760 45540
rect 8680 45460 8760 45480
rect 8330 45410 8340 45450
rect 8448 45444 8648 45450
rect 8260 45400 8340 45410
rect 7730 44240 7800 45390
rect 7730 43980 7750 44240
rect 7790 43980 7800 44240
rect 8810 45390 8820 45630
rect 8860 45390 8880 45630
rect 8810 44240 8880 45390
rect 8260 44210 8340 44220
rect 7950 44172 8150 44178
rect 7840 44140 7920 44160
rect 7840 44080 7850 44140
rect 7910 44128 7920 44140
rect 7950 44138 7962 44172
rect 8138 44170 8150 44172
rect 8260 44170 8270 44210
rect 8138 44150 8270 44170
rect 8330 44170 8340 44210
rect 8448 44172 8648 44178
rect 8448 44170 8460 44172
rect 8330 44150 8460 44170
rect 8138 44140 8460 44150
rect 8138 44138 8150 44140
rect 7950 44132 8150 44138
rect 8448 44138 8460 44140
rect 8636 44138 8648 44172
rect 8448 44132 8648 44138
rect 8680 44140 8760 44160
rect 7912 44094 7920 44128
rect 7910 44080 7920 44094
rect 7840 44060 7920 44080
rect 7950 44084 8150 44090
rect 7950 44050 7962 44084
rect 8138 44080 8150 44084
rect 8448 44084 8648 44090
rect 8448 44080 8460 44084
rect 8138 44050 8460 44080
rect 8636 44050 8648 44084
rect 8680 44080 8690 44140
rect 8750 44080 8760 44140
rect 8680 44060 8760 44080
rect 7950 44044 8150 44050
rect 7730 43920 7800 43980
rect 7730 43680 7750 43920
rect 7790 43680 7800 43920
rect 8260 44040 8340 44050
rect 8448 44044 8648 44050
rect 8260 43980 8270 44040
rect 8330 43980 8340 44040
rect 8260 43930 8340 43980
rect 8260 43870 8270 43930
rect 8330 43870 8340 43930
rect 7950 43862 8150 43868
rect 7840 43830 7920 43850
rect 7840 43770 7850 43830
rect 7910 43818 7920 43830
rect 7950 43828 7962 43862
rect 8138 43860 8150 43862
rect 8260 43860 8340 43870
rect 8810 44000 8820 44240
rect 8860 44000 8880 44240
rect 8810 43920 8880 44000
rect 8448 43862 8648 43868
rect 8448 43860 8460 43862
rect 8138 43830 8460 43860
rect 8138 43828 8150 43830
rect 7950 43822 8150 43828
rect 8448 43828 8460 43830
rect 8636 43828 8648 43862
rect 8448 43822 8648 43828
rect 8680 43830 8760 43850
rect 7912 43784 7920 43818
rect 7910 43770 7920 43784
rect 7840 43750 7920 43770
rect 7950 43774 8150 43780
rect 7950 43740 7962 43774
rect 8138 43770 8150 43774
rect 8448 43774 8648 43780
rect 8448 43770 8460 43774
rect 8138 43760 8460 43770
rect 8138 43740 8270 43760
rect 7950 43734 8150 43740
rect 8260 43700 8270 43740
rect 8330 43740 8460 43760
rect 8636 43740 8648 43774
rect 8680 43770 8690 43830
rect 8750 43770 8760 43830
rect 8680 43750 8760 43770
rect 8330 43700 8340 43740
rect 8448 43734 8648 43740
rect 8260 43690 8340 43700
rect 7730 42530 7800 43680
rect 7730 42270 7750 42530
rect 7790 42270 7800 42530
rect 8810 43680 8820 43920
rect 8860 43680 8880 43920
rect 8810 42530 8880 43680
rect 8260 42500 8340 42510
rect 7950 42462 8150 42468
rect 7840 42430 7920 42450
rect 7840 42370 7850 42430
rect 7910 42418 7920 42430
rect 7950 42428 7962 42462
rect 8138 42460 8150 42462
rect 8260 42460 8270 42500
rect 8138 42440 8270 42460
rect 8330 42460 8340 42500
rect 8448 42462 8648 42468
rect 8448 42460 8460 42462
rect 8330 42440 8460 42460
rect 8138 42430 8460 42440
rect 8138 42428 8150 42430
rect 7950 42422 8150 42428
rect 8448 42428 8460 42430
rect 8636 42428 8648 42462
rect 8448 42422 8648 42428
rect 8680 42430 8760 42450
rect 7912 42384 7920 42418
rect 7910 42370 7920 42384
rect 7840 42350 7920 42370
rect 7950 42374 8150 42380
rect 7950 42340 7962 42374
rect 8138 42370 8150 42374
rect 8448 42374 8648 42380
rect 8448 42370 8460 42374
rect 8138 42340 8460 42370
rect 8636 42340 8648 42374
rect 8680 42370 8690 42430
rect 8750 42370 8760 42430
rect 8680 42350 8760 42370
rect 7950 42334 8150 42340
rect 7730 42210 7800 42270
rect 7730 41970 7750 42210
rect 7790 41970 7800 42210
rect 8260 42330 8340 42340
rect 8448 42334 8648 42340
rect 8260 42270 8270 42330
rect 8330 42270 8340 42330
rect 8260 42220 8340 42270
rect 8260 42160 8270 42220
rect 8330 42160 8340 42220
rect 7950 42152 8150 42158
rect 7840 42120 7920 42140
rect 7840 42060 7850 42120
rect 7910 42108 7920 42120
rect 7950 42118 7962 42152
rect 8138 42150 8150 42152
rect 8260 42150 8340 42160
rect 8810 42290 8820 42530
rect 8860 42290 8880 42530
rect 8810 42210 8880 42290
rect 8448 42152 8648 42158
rect 8448 42150 8460 42152
rect 8138 42120 8460 42150
rect 8138 42118 8150 42120
rect 7950 42112 8150 42118
rect 8448 42118 8460 42120
rect 8636 42118 8648 42152
rect 8448 42112 8648 42118
rect 8680 42120 8760 42140
rect 7912 42074 7920 42108
rect 7910 42060 7920 42074
rect 7840 42040 7920 42060
rect 7950 42064 8150 42070
rect 7950 42030 7962 42064
rect 8138 42060 8150 42064
rect 8448 42064 8648 42070
rect 8448 42060 8460 42064
rect 8138 42050 8460 42060
rect 8138 42030 8270 42050
rect 7950 42024 8150 42030
rect 8260 41990 8270 42030
rect 8330 42030 8460 42050
rect 8636 42030 8648 42064
rect 8680 42060 8690 42120
rect 8750 42060 8760 42120
rect 8680 42040 8760 42060
rect 8330 41990 8340 42030
rect 8448 42024 8648 42030
rect 8260 41980 8340 41990
rect 7730 40820 7800 41970
rect 7730 40560 7750 40820
rect 7790 40560 7800 40820
rect 8810 41970 8820 42210
rect 8860 41970 8880 42210
rect 8810 40820 8880 41970
rect 8260 40790 8340 40800
rect 7950 40752 8150 40758
rect 7840 40720 7920 40740
rect 7840 40660 7850 40720
rect 7910 40708 7920 40720
rect 7950 40718 7962 40752
rect 8138 40750 8150 40752
rect 8260 40750 8270 40790
rect 8138 40730 8270 40750
rect 8330 40750 8340 40790
rect 8448 40752 8648 40758
rect 8448 40750 8460 40752
rect 8330 40730 8460 40750
rect 8138 40720 8460 40730
rect 8138 40718 8150 40720
rect 7950 40712 8150 40718
rect 8448 40718 8460 40720
rect 8636 40718 8648 40752
rect 8448 40712 8648 40718
rect 8680 40720 8760 40740
rect 7912 40674 7920 40708
rect 7910 40660 7920 40674
rect 7840 40640 7920 40660
rect 7950 40664 8150 40670
rect 7950 40630 7962 40664
rect 8138 40660 8150 40664
rect 8448 40664 8648 40670
rect 8448 40660 8460 40664
rect 8138 40630 8460 40660
rect 8636 40630 8648 40664
rect 8680 40660 8690 40720
rect 8750 40660 8760 40720
rect 8680 40640 8760 40660
rect 7950 40624 8150 40630
rect 7730 40500 7800 40560
rect 7730 40260 7750 40500
rect 7790 40260 7800 40500
rect 8260 40620 8340 40630
rect 8448 40624 8648 40630
rect 8260 40560 8270 40620
rect 8330 40560 8340 40620
rect 8260 40510 8340 40560
rect 8260 40450 8270 40510
rect 8330 40450 8340 40510
rect 7950 40442 8150 40448
rect 7840 40410 7920 40430
rect 7840 40350 7850 40410
rect 7910 40398 7920 40410
rect 7950 40408 7962 40442
rect 8138 40440 8150 40442
rect 8260 40440 8340 40450
rect 8810 40580 8820 40820
rect 8860 40580 8880 40820
rect 8810 40500 8880 40580
rect 8448 40442 8648 40448
rect 8448 40440 8460 40442
rect 8138 40410 8460 40440
rect 8138 40408 8150 40410
rect 7950 40402 8150 40408
rect 8448 40408 8460 40410
rect 8636 40408 8648 40442
rect 8448 40402 8648 40408
rect 8680 40410 8760 40430
rect 7912 40364 7920 40398
rect 7910 40350 7920 40364
rect 7840 40330 7920 40350
rect 7950 40354 8150 40360
rect 7950 40320 7962 40354
rect 8138 40350 8150 40354
rect 8448 40354 8648 40360
rect 8448 40350 8460 40354
rect 8138 40340 8460 40350
rect 8138 40320 8270 40340
rect 7950 40314 8150 40320
rect 8260 40280 8270 40320
rect 8330 40320 8460 40340
rect 8636 40320 8648 40354
rect 8680 40350 8690 40410
rect 8750 40350 8760 40410
rect 8680 40330 8760 40350
rect 8330 40280 8340 40320
rect 8448 40314 8648 40320
rect 8260 40270 8340 40280
rect 7730 39690 7800 40260
rect 8810 40260 8820 40500
rect 8860 40260 8880 40500
rect 8810 39690 8880 40260
rect 7730 39680 7810 39690
rect 7730 39620 7740 39680
rect 7800 39620 7810 39680
rect 8800 39680 8880 39690
rect 8800 39620 8810 39680
rect 8870 39620 8880 39680
rect 8800 39610 8880 39620
rect 8910 66480 8940 67050
rect 8910 66470 8970 66480
rect 8910 66400 8970 66410
rect 8910 64770 8940 66400
rect 9000 65950 9030 67050
rect 8970 65940 9030 65950
rect 8970 65870 9030 65880
rect 8910 64760 8970 64770
rect 8910 64690 8970 64700
rect 8910 63060 8940 64690
rect 9000 64240 9030 65870
rect 8970 64230 9030 64240
rect 8970 64160 9030 64170
rect 8910 63050 8970 63060
rect 8910 62980 8970 62990
rect 8910 61350 8940 62980
rect 9000 62530 9030 64160
rect 8970 62520 9030 62530
rect 8970 62450 9030 62460
rect 8910 61340 8970 61350
rect 8910 61270 8970 61280
rect 8910 59640 8940 61270
rect 9000 60820 9030 62450
rect 8970 60810 9030 60820
rect 8970 60740 9030 60750
rect 8910 59630 8970 59640
rect 8910 59560 8970 59570
rect 8910 57930 8940 59560
rect 9000 59110 9030 60740
rect 8970 59100 9030 59110
rect 8970 59030 9030 59040
rect 8910 57920 8970 57930
rect 8910 57850 8970 57860
rect 8910 56220 8940 57850
rect 9000 57400 9030 59030
rect 8970 57390 9030 57400
rect 8970 57320 9030 57330
rect 8910 56210 8970 56220
rect 8910 56140 8970 56150
rect 8910 54510 8940 56140
rect 9000 55690 9030 57320
rect 8970 55680 9030 55690
rect 8970 55610 9030 55620
rect 8910 54500 8970 54510
rect 8910 54430 8970 54440
rect 8910 52800 8940 54430
rect 9000 53980 9030 55610
rect 8970 53970 9030 53980
rect 8970 53900 9030 53910
rect 8910 52790 8970 52800
rect 8910 52720 8970 52730
rect 8910 51090 8940 52720
rect 9000 52270 9030 53900
rect 8970 52260 9030 52270
rect 8970 52190 9030 52200
rect 8910 51080 8970 51090
rect 8910 51010 8970 51020
rect 8910 49380 8940 51010
rect 9000 50560 9030 52190
rect 8970 50550 9030 50560
rect 8970 50480 9030 50490
rect 8910 49370 8970 49380
rect 8910 49300 8970 49310
rect 8910 47670 8940 49300
rect 9000 48850 9030 50480
rect 8970 48840 9030 48850
rect 8970 48770 9030 48780
rect 8910 47660 8970 47670
rect 8910 47590 8970 47600
rect 8910 45960 8940 47590
rect 9000 47140 9030 48770
rect 8970 47130 9030 47140
rect 8970 47060 9030 47070
rect 8910 45950 8970 45960
rect 8910 45880 8970 45890
rect 8910 44250 8940 45880
rect 9000 45430 9030 47060
rect 8970 45420 9030 45430
rect 8970 45350 9030 45360
rect 8910 44240 8970 44250
rect 8910 44170 8970 44180
rect 8910 42540 8940 44170
rect 9000 43720 9030 45350
rect 8970 43710 9030 43720
rect 8970 43640 9030 43650
rect 8910 42530 8970 42540
rect 8910 42460 8970 42470
rect 8910 40830 8940 42460
rect 9000 42010 9030 43640
rect 8970 42000 9030 42010
rect 8970 41930 9030 41940
rect 8910 40820 8970 40830
rect 8910 40750 8970 40760
rect 4070 39230 4330 39240
rect 4070 39210 4270 39230
rect 4270 39160 4330 39170
rect 7440 39230 7700 39240
rect 7500 39210 7700 39230
rect 7440 39160 7500 39170
rect 8910 38840 8940 40750
rect 9000 40300 9030 41930
rect 8970 40290 9030 40300
rect 8970 40220 9030 40230
rect 9000 39690 9030 40220
rect 8970 39680 9030 39690
rect 8970 39610 9030 39620
rect 9060 66390 9090 67050
rect 9060 66380 9120 66390
rect 9060 66310 9120 66320
rect 9060 64680 9090 66310
rect 9060 64670 9120 64680
rect 9060 64600 9120 64610
rect 9060 62970 9090 64600
rect 9060 62960 9120 62970
rect 9060 62890 9120 62900
rect 9060 61260 9090 62890
rect 9060 61250 9120 61260
rect 9060 61180 9120 61190
rect 9060 59550 9090 61180
rect 9060 59540 9120 59550
rect 9060 59470 9120 59480
rect 9060 57840 9090 59470
rect 9060 57830 9120 57840
rect 9060 57760 9120 57770
rect 9060 56130 9090 57760
rect 9060 56120 9120 56130
rect 9060 56050 9120 56060
rect 9060 54420 9090 56050
rect 9060 54410 9120 54420
rect 9060 54340 9120 54350
rect 9060 52710 9090 54340
rect 9060 52700 9120 52710
rect 9060 52630 9120 52640
rect 9060 51000 9090 52630
rect 9060 50990 9120 51000
rect 9060 50920 9120 50930
rect 9060 49290 9090 50920
rect 9060 49280 9120 49290
rect 9060 49210 9120 49220
rect 9060 47580 9090 49210
rect 9060 47570 9120 47580
rect 9060 47500 9120 47510
rect 9060 45870 9090 47500
rect 9060 45860 9120 45870
rect 9060 45790 9120 45800
rect 9060 44160 9090 45790
rect 9060 44150 9120 44160
rect 9060 44080 9120 44090
rect 9060 42450 9090 44080
rect 9060 42440 9120 42450
rect 9060 42370 9120 42380
rect 9060 40740 9090 42370
rect 9060 40730 9120 40740
rect 9060 40660 9120 40670
rect 9060 39240 9090 40660
rect 9180 39690 9210 67050
rect 9300 39690 9330 67050
rect 9420 39690 9450 67050
rect 9540 39690 9570 67050
rect 9660 39690 9690 67050
rect 9780 39690 9810 67050
rect 11940 39690 11970 67050
rect 12060 39690 12090 67050
rect 12180 39690 12210 67050
rect 12300 39690 12330 67050
rect 12420 39690 12450 67050
rect 12540 59550 12570 67050
rect 12660 66390 12690 67050
rect 12630 66380 12690 66390
rect 12630 66310 12690 66320
rect 12660 64680 12690 66310
rect 12630 64670 12690 64680
rect 12630 64600 12690 64610
rect 12660 62970 12690 64600
rect 12630 62960 12690 62970
rect 12630 62890 12690 62900
rect 12660 61260 12690 62890
rect 12630 61250 12690 61260
rect 12630 61180 12690 61190
rect 12510 59540 12570 59550
rect 12510 59470 12570 59480
rect 12540 57840 12570 59470
rect 12510 57830 12570 57840
rect 12510 57760 12570 57770
rect 12540 56130 12570 57760
rect 12510 56120 12570 56130
rect 12510 56050 12570 56060
rect 12540 54420 12570 56050
rect 12510 54410 12570 54420
rect 12510 54340 12570 54350
rect 12540 52710 12570 54340
rect 12510 52700 12570 52710
rect 12510 52630 12570 52640
rect 12540 51000 12570 52630
rect 12510 50990 12570 51000
rect 12510 50920 12570 50930
rect 12540 49290 12570 50920
rect 12510 49280 12570 49290
rect 12510 49210 12570 49220
rect 12540 47580 12570 49210
rect 12510 47570 12570 47580
rect 12510 47500 12570 47510
rect 12540 39300 12570 47500
rect 12660 45870 12690 61180
rect 12630 45860 12690 45870
rect 12630 45790 12690 45800
rect 12660 44160 12690 45790
rect 12630 44150 12690 44160
rect 12630 44080 12690 44090
rect 12660 42450 12690 44080
rect 12630 42440 12690 42450
rect 12630 42370 12690 42380
rect 12660 40740 12690 42370
rect 12630 40730 12690 40740
rect 12630 40660 12690 40670
rect 12250 39290 12570 39300
rect 9060 39230 9320 39240
rect 9060 39210 9260 39230
rect 12310 39270 12570 39290
rect 12660 39240 12690 40660
rect 12720 66470 12790 67050
rect 12720 66210 12740 66470
rect 12780 66210 12790 66470
rect 13800 66470 13870 67050
rect 13250 66440 13330 66450
rect 12940 66402 13140 66408
rect 12830 66370 12910 66390
rect 12830 66310 12840 66370
rect 12900 66358 12910 66370
rect 12940 66368 12952 66402
rect 13128 66400 13140 66402
rect 13250 66400 13260 66440
rect 13128 66380 13260 66400
rect 13320 66400 13330 66440
rect 13438 66402 13638 66408
rect 13438 66400 13450 66402
rect 13320 66380 13450 66400
rect 13128 66370 13450 66380
rect 13128 66368 13140 66370
rect 12940 66362 13140 66368
rect 13438 66368 13450 66370
rect 13626 66368 13638 66402
rect 13438 66362 13638 66368
rect 13670 66370 13750 66390
rect 12902 66324 12910 66358
rect 12900 66310 12910 66324
rect 12830 66290 12910 66310
rect 12940 66314 13140 66320
rect 12940 66280 12952 66314
rect 13128 66310 13140 66314
rect 13438 66314 13638 66320
rect 13438 66310 13450 66314
rect 13128 66280 13450 66310
rect 13626 66280 13638 66314
rect 13670 66310 13680 66370
rect 13740 66310 13750 66370
rect 13670 66290 13750 66310
rect 12940 66274 13140 66280
rect 12720 66150 12790 66210
rect 12720 65910 12740 66150
rect 12780 65910 12790 66150
rect 13250 66270 13330 66280
rect 13438 66274 13638 66280
rect 13250 66210 13260 66270
rect 13320 66210 13330 66270
rect 13250 66160 13330 66210
rect 13250 66100 13260 66160
rect 13320 66100 13330 66160
rect 12940 66092 13140 66098
rect 12830 66060 12910 66080
rect 12830 66000 12840 66060
rect 12900 66048 12910 66060
rect 12940 66058 12952 66092
rect 13128 66090 13140 66092
rect 13250 66090 13330 66100
rect 13800 66230 13810 66470
rect 13850 66230 13870 66470
rect 13800 66150 13870 66230
rect 13438 66092 13638 66098
rect 13438 66090 13450 66092
rect 13128 66060 13450 66090
rect 13128 66058 13140 66060
rect 12940 66052 13140 66058
rect 13438 66058 13450 66060
rect 13626 66058 13638 66092
rect 13438 66052 13638 66058
rect 13670 66060 13750 66080
rect 12902 66014 12910 66048
rect 12900 66000 12910 66014
rect 12830 65980 12910 66000
rect 12940 66004 13140 66010
rect 12940 65970 12952 66004
rect 13128 66000 13140 66004
rect 13438 66004 13638 66010
rect 13438 66000 13450 66004
rect 13128 65990 13450 66000
rect 13128 65970 13260 65990
rect 12940 65964 13140 65970
rect 13250 65930 13260 65970
rect 13320 65970 13450 65990
rect 13626 65970 13638 66004
rect 13670 66000 13680 66060
rect 13740 66000 13750 66060
rect 13670 65980 13750 66000
rect 13320 65930 13330 65970
rect 13438 65964 13638 65970
rect 13250 65920 13330 65930
rect 12720 64760 12790 65910
rect 12720 64500 12740 64760
rect 12780 64500 12790 64760
rect 13800 65910 13810 66150
rect 13850 65910 13870 66150
rect 13800 64760 13870 65910
rect 13250 64730 13330 64740
rect 12940 64692 13140 64698
rect 12830 64660 12910 64680
rect 12830 64600 12840 64660
rect 12900 64648 12910 64660
rect 12940 64658 12952 64692
rect 13128 64690 13140 64692
rect 13250 64690 13260 64730
rect 13128 64670 13260 64690
rect 13320 64690 13330 64730
rect 13438 64692 13638 64698
rect 13438 64690 13450 64692
rect 13320 64670 13450 64690
rect 13128 64660 13450 64670
rect 13128 64658 13140 64660
rect 12940 64652 13140 64658
rect 13438 64658 13450 64660
rect 13626 64658 13638 64692
rect 13438 64652 13638 64658
rect 13670 64660 13750 64680
rect 12902 64614 12910 64648
rect 12900 64600 12910 64614
rect 12830 64580 12910 64600
rect 12940 64604 13140 64610
rect 12940 64570 12952 64604
rect 13128 64600 13140 64604
rect 13438 64604 13638 64610
rect 13438 64600 13450 64604
rect 13128 64570 13450 64600
rect 13626 64570 13638 64604
rect 13670 64600 13680 64660
rect 13740 64600 13750 64660
rect 13670 64580 13750 64600
rect 12940 64564 13140 64570
rect 12720 64440 12790 64500
rect 12720 64200 12740 64440
rect 12780 64200 12790 64440
rect 13250 64560 13330 64570
rect 13438 64564 13638 64570
rect 13250 64500 13260 64560
rect 13320 64500 13330 64560
rect 13250 64450 13330 64500
rect 13250 64390 13260 64450
rect 13320 64390 13330 64450
rect 12940 64382 13140 64388
rect 12830 64350 12910 64370
rect 12830 64290 12840 64350
rect 12900 64338 12910 64350
rect 12940 64348 12952 64382
rect 13128 64380 13140 64382
rect 13250 64380 13330 64390
rect 13800 64520 13810 64760
rect 13850 64520 13870 64760
rect 13800 64440 13870 64520
rect 13438 64382 13638 64388
rect 13438 64380 13450 64382
rect 13128 64350 13450 64380
rect 13128 64348 13140 64350
rect 12940 64342 13140 64348
rect 13438 64348 13450 64350
rect 13626 64348 13638 64382
rect 13438 64342 13638 64348
rect 13670 64350 13750 64370
rect 12902 64304 12910 64338
rect 12900 64290 12910 64304
rect 12830 64270 12910 64290
rect 12940 64294 13140 64300
rect 12940 64260 12952 64294
rect 13128 64290 13140 64294
rect 13438 64294 13638 64300
rect 13438 64290 13450 64294
rect 13128 64280 13450 64290
rect 13128 64260 13260 64280
rect 12940 64254 13140 64260
rect 13250 64220 13260 64260
rect 13320 64260 13450 64280
rect 13626 64260 13638 64294
rect 13670 64290 13680 64350
rect 13740 64290 13750 64350
rect 13670 64270 13750 64290
rect 13320 64220 13330 64260
rect 13438 64254 13638 64260
rect 13250 64210 13330 64220
rect 12720 63050 12790 64200
rect 12720 62790 12740 63050
rect 12780 62790 12790 63050
rect 13800 64200 13810 64440
rect 13850 64200 13870 64440
rect 13800 63050 13870 64200
rect 13250 63020 13330 63030
rect 12940 62982 13140 62988
rect 12830 62950 12910 62970
rect 12830 62890 12840 62950
rect 12900 62938 12910 62950
rect 12940 62948 12952 62982
rect 13128 62980 13140 62982
rect 13250 62980 13260 63020
rect 13128 62960 13260 62980
rect 13320 62980 13330 63020
rect 13438 62982 13638 62988
rect 13438 62980 13450 62982
rect 13320 62960 13450 62980
rect 13128 62950 13450 62960
rect 13128 62948 13140 62950
rect 12940 62942 13140 62948
rect 13438 62948 13450 62950
rect 13626 62948 13638 62982
rect 13438 62942 13638 62948
rect 13670 62950 13750 62970
rect 12902 62904 12910 62938
rect 12900 62890 12910 62904
rect 12830 62870 12910 62890
rect 12940 62894 13140 62900
rect 12940 62860 12952 62894
rect 13128 62890 13140 62894
rect 13438 62894 13638 62900
rect 13438 62890 13450 62894
rect 13128 62860 13450 62890
rect 13626 62860 13638 62894
rect 13670 62890 13680 62950
rect 13740 62890 13750 62950
rect 13670 62870 13750 62890
rect 12940 62854 13140 62860
rect 12720 62730 12790 62790
rect 12720 62490 12740 62730
rect 12780 62490 12790 62730
rect 13250 62850 13330 62860
rect 13438 62854 13638 62860
rect 13250 62790 13260 62850
rect 13320 62790 13330 62850
rect 13250 62740 13330 62790
rect 13250 62680 13260 62740
rect 13320 62680 13330 62740
rect 12940 62672 13140 62678
rect 12830 62640 12910 62660
rect 12830 62580 12840 62640
rect 12900 62628 12910 62640
rect 12940 62638 12952 62672
rect 13128 62670 13140 62672
rect 13250 62670 13330 62680
rect 13800 62810 13810 63050
rect 13850 62810 13870 63050
rect 13800 62730 13870 62810
rect 13438 62672 13638 62678
rect 13438 62670 13450 62672
rect 13128 62640 13450 62670
rect 13128 62638 13140 62640
rect 12940 62632 13140 62638
rect 13438 62638 13450 62640
rect 13626 62638 13638 62672
rect 13438 62632 13638 62638
rect 13670 62640 13750 62660
rect 12902 62594 12910 62628
rect 12900 62580 12910 62594
rect 12830 62560 12910 62580
rect 12940 62584 13140 62590
rect 12940 62550 12952 62584
rect 13128 62580 13140 62584
rect 13438 62584 13638 62590
rect 13438 62580 13450 62584
rect 13128 62570 13450 62580
rect 13128 62550 13260 62570
rect 12940 62544 13140 62550
rect 13250 62510 13260 62550
rect 13320 62550 13450 62570
rect 13626 62550 13638 62584
rect 13670 62580 13680 62640
rect 13740 62580 13750 62640
rect 13670 62560 13750 62580
rect 13320 62510 13330 62550
rect 13438 62544 13638 62550
rect 13250 62500 13330 62510
rect 12720 61340 12790 62490
rect 12720 61080 12740 61340
rect 12780 61080 12790 61340
rect 13800 62490 13810 62730
rect 13850 62490 13870 62730
rect 13800 61340 13870 62490
rect 13250 61310 13330 61320
rect 12940 61272 13140 61278
rect 12830 61240 12910 61260
rect 12830 61180 12840 61240
rect 12900 61228 12910 61240
rect 12940 61238 12952 61272
rect 13128 61270 13140 61272
rect 13250 61270 13260 61310
rect 13128 61250 13260 61270
rect 13320 61270 13330 61310
rect 13438 61272 13638 61278
rect 13438 61270 13450 61272
rect 13320 61250 13450 61270
rect 13128 61240 13450 61250
rect 13128 61238 13140 61240
rect 12940 61232 13140 61238
rect 13438 61238 13450 61240
rect 13626 61238 13638 61272
rect 13438 61232 13638 61238
rect 13670 61240 13750 61260
rect 12902 61194 12910 61228
rect 12900 61180 12910 61194
rect 12830 61160 12910 61180
rect 12940 61184 13140 61190
rect 12940 61150 12952 61184
rect 13128 61180 13140 61184
rect 13438 61184 13638 61190
rect 13438 61180 13450 61184
rect 13128 61150 13450 61180
rect 13626 61150 13638 61184
rect 13670 61180 13680 61240
rect 13740 61180 13750 61240
rect 13670 61160 13750 61180
rect 12940 61144 13140 61150
rect 12720 61020 12790 61080
rect 12720 60780 12740 61020
rect 12780 60780 12790 61020
rect 13250 61140 13330 61150
rect 13438 61144 13638 61150
rect 13250 61080 13260 61140
rect 13320 61080 13330 61140
rect 13250 61030 13330 61080
rect 13250 60970 13260 61030
rect 13320 60970 13330 61030
rect 12940 60962 13140 60968
rect 12830 60930 12910 60950
rect 12830 60870 12840 60930
rect 12900 60918 12910 60930
rect 12940 60928 12952 60962
rect 13128 60960 13140 60962
rect 13250 60960 13330 60970
rect 13800 61100 13810 61340
rect 13850 61100 13870 61340
rect 13800 61020 13870 61100
rect 13438 60962 13638 60968
rect 13438 60960 13450 60962
rect 13128 60930 13450 60960
rect 13128 60928 13140 60930
rect 12940 60922 13140 60928
rect 13438 60928 13450 60930
rect 13626 60928 13638 60962
rect 13438 60922 13638 60928
rect 13670 60930 13750 60950
rect 12902 60884 12910 60918
rect 12900 60870 12910 60884
rect 12830 60850 12910 60870
rect 12940 60874 13140 60880
rect 12940 60840 12952 60874
rect 13128 60870 13140 60874
rect 13438 60874 13638 60880
rect 13438 60870 13450 60874
rect 13128 60860 13450 60870
rect 13128 60840 13260 60860
rect 12940 60834 13140 60840
rect 13250 60800 13260 60840
rect 13320 60840 13450 60860
rect 13626 60840 13638 60874
rect 13670 60870 13680 60930
rect 13740 60870 13750 60930
rect 13670 60850 13750 60870
rect 13320 60800 13330 60840
rect 13438 60834 13638 60840
rect 13250 60790 13330 60800
rect 12720 59630 12790 60780
rect 12720 59370 12740 59630
rect 12780 59370 12790 59630
rect 13800 60780 13810 61020
rect 13850 60780 13870 61020
rect 13800 59630 13870 60780
rect 13250 59600 13330 59610
rect 12940 59562 13140 59568
rect 12830 59530 12910 59550
rect 12830 59470 12840 59530
rect 12900 59518 12910 59530
rect 12940 59528 12952 59562
rect 13128 59560 13140 59562
rect 13250 59560 13260 59600
rect 13128 59540 13260 59560
rect 13320 59560 13330 59600
rect 13438 59562 13638 59568
rect 13438 59560 13450 59562
rect 13320 59540 13450 59560
rect 13128 59530 13450 59540
rect 13128 59528 13140 59530
rect 12940 59522 13140 59528
rect 13438 59528 13450 59530
rect 13626 59528 13638 59562
rect 13438 59522 13638 59528
rect 13670 59530 13750 59550
rect 12902 59484 12910 59518
rect 12900 59470 12910 59484
rect 12830 59450 12910 59470
rect 12940 59474 13140 59480
rect 12940 59440 12952 59474
rect 13128 59470 13140 59474
rect 13438 59474 13638 59480
rect 13438 59470 13450 59474
rect 13128 59440 13450 59470
rect 13626 59440 13638 59474
rect 13670 59470 13680 59530
rect 13740 59470 13750 59530
rect 13670 59450 13750 59470
rect 12940 59434 13140 59440
rect 12720 59310 12790 59370
rect 12720 59070 12740 59310
rect 12780 59070 12790 59310
rect 13250 59430 13330 59440
rect 13438 59434 13638 59440
rect 13250 59370 13260 59430
rect 13320 59370 13330 59430
rect 13250 59320 13330 59370
rect 13250 59260 13260 59320
rect 13320 59260 13330 59320
rect 12940 59252 13140 59258
rect 12830 59220 12910 59240
rect 12830 59160 12840 59220
rect 12900 59208 12910 59220
rect 12940 59218 12952 59252
rect 13128 59250 13140 59252
rect 13250 59250 13330 59260
rect 13800 59390 13810 59630
rect 13850 59390 13870 59630
rect 13800 59310 13870 59390
rect 13438 59252 13638 59258
rect 13438 59250 13450 59252
rect 13128 59220 13450 59250
rect 13128 59218 13140 59220
rect 12940 59212 13140 59218
rect 13438 59218 13450 59220
rect 13626 59218 13638 59252
rect 13438 59212 13638 59218
rect 13670 59220 13750 59240
rect 12902 59174 12910 59208
rect 12900 59160 12910 59174
rect 12830 59140 12910 59160
rect 12940 59164 13140 59170
rect 12940 59130 12952 59164
rect 13128 59160 13140 59164
rect 13438 59164 13638 59170
rect 13438 59160 13450 59164
rect 13128 59150 13450 59160
rect 13128 59130 13260 59150
rect 12940 59124 13140 59130
rect 13250 59090 13260 59130
rect 13320 59130 13450 59150
rect 13626 59130 13638 59164
rect 13670 59160 13680 59220
rect 13740 59160 13750 59220
rect 13670 59140 13750 59160
rect 13320 59090 13330 59130
rect 13438 59124 13638 59130
rect 13250 59080 13330 59090
rect 12720 57920 12790 59070
rect 12720 57660 12740 57920
rect 12780 57660 12790 57920
rect 13800 59070 13810 59310
rect 13850 59070 13870 59310
rect 13800 57920 13870 59070
rect 13250 57890 13330 57900
rect 12940 57852 13140 57858
rect 12830 57820 12910 57840
rect 12830 57760 12840 57820
rect 12900 57808 12910 57820
rect 12940 57818 12952 57852
rect 13128 57850 13140 57852
rect 13250 57850 13260 57890
rect 13128 57830 13260 57850
rect 13320 57850 13330 57890
rect 13438 57852 13638 57858
rect 13438 57850 13450 57852
rect 13320 57830 13450 57850
rect 13128 57820 13450 57830
rect 13128 57818 13140 57820
rect 12940 57812 13140 57818
rect 13438 57818 13450 57820
rect 13626 57818 13638 57852
rect 13438 57812 13638 57818
rect 13670 57820 13750 57840
rect 12902 57774 12910 57808
rect 12900 57760 12910 57774
rect 12830 57740 12910 57760
rect 12940 57764 13140 57770
rect 12940 57730 12952 57764
rect 13128 57760 13140 57764
rect 13438 57764 13638 57770
rect 13438 57760 13450 57764
rect 13128 57730 13450 57760
rect 13626 57730 13638 57764
rect 13670 57760 13680 57820
rect 13740 57760 13750 57820
rect 13670 57740 13750 57760
rect 12940 57724 13140 57730
rect 12720 57600 12790 57660
rect 12720 57360 12740 57600
rect 12780 57360 12790 57600
rect 13250 57720 13330 57730
rect 13438 57724 13638 57730
rect 13250 57660 13260 57720
rect 13320 57660 13330 57720
rect 13250 57610 13330 57660
rect 13250 57550 13260 57610
rect 13320 57550 13330 57610
rect 12940 57542 13140 57548
rect 12830 57510 12910 57530
rect 12830 57450 12840 57510
rect 12900 57498 12910 57510
rect 12940 57508 12952 57542
rect 13128 57540 13140 57542
rect 13250 57540 13330 57550
rect 13800 57680 13810 57920
rect 13850 57680 13870 57920
rect 13800 57600 13870 57680
rect 13438 57542 13638 57548
rect 13438 57540 13450 57542
rect 13128 57510 13450 57540
rect 13128 57508 13140 57510
rect 12940 57502 13140 57508
rect 13438 57508 13450 57510
rect 13626 57508 13638 57542
rect 13438 57502 13638 57508
rect 13670 57510 13750 57530
rect 12902 57464 12910 57498
rect 12900 57450 12910 57464
rect 12830 57430 12910 57450
rect 12940 57454 13140 57460
rect 12940 57420 12952 57454
rect 13128 57450 13140 57454
rect 13438 57454 13638 57460
rect 13438 57450 13450 57454
rect 13128 57440 13450 57450
rect 13128 57420 13260 57440
rect 12940 57414 13140 57420
rect 13250 57380 13260 57420
rect 13320 57420 13450 57440
rect 13626 57420 13638 57454
rect 13670 57450 13680 57510
rect 13740 57450 13750 57510
rect 13670 57430 13750 57450
rect 13320 57380 13330 57420
rect 13438 57414 13638 57420
rect 13250 57370 13330 57380
rect 12720 56210 12790 57360
rect 12720 55950 12740 56210
rect 12780 55950 12790 56210
rect 13800 57360 13810 57600
rect 13850 57360 13870 57600
rect 13800 56210 13870 57360
rect 13250 56180 13330 56190
rect 12940 56142 13140 56148
rect 12830 56110 12910 56130
rect 12830 56050 12840 56110
rect 12900 56098 12910 56110
rect 12940 56108 12952 56142
rect 13128 56140 13140 56142
rect 13250 56140 13260 56180
rect 13128 56120 13260 56140
rect 13320 56140 13330 56180
rect 13438 56142 13638 56148
rect 13438 56140 13450 56142
rect 13320 56120 13450 56140
rect 13128 56110 13450 56120
rect 13128 56108 13140 56110
rect 12940 56102 13140 56108
rect 13438 56108 13450 56110
rect 13626 56108 13638 56142
rect 13438 56102 13638 56108
rect 13670 56110 13750 56130
rect 12902 56064 12910 56098
rect 12900 56050 12910 56064
rect 12830 56030 12910 56050
rect 12940 56054 13140 56060
rect 12940 56020 12952 56054
rect 13128 56050 13140 56054
rect 13438 56054 13638 56060
rect 13438 56050 13450 56054
rect 13128 56020 13450 56050
rect 13626 56020 13638 56054
rect 13670 56050 13680 56110
rect 13740 56050 13750 56110
rect 13670 56030 13750 56050
rect 12940 56014 13140 56020
rect 12720 55890 12790 55950
rect 12720 55650 12740 55890
rect 12780 55650 12790 55890
rect 13250 56010 13330 56020
rect 13438 56014 13638 56020
rect 13250 55950 13260 56010
rect 13320 55950 13330 56010
rect 13250 55900 13330 55950
rect 13250 55840 13260 55900
rect 13320 55840 13330 55900
rect 12940 55832 13140 55838
rect 12830 55800 12910 55820
rect 12830 55740 12840 55800
rect 12900 55788 12910 55800
rect 12940 55798 12952 55832
rect 13128 55830 13140 55832
rect 13250 55830 13330 55840
rect 13800 55970 13810 56210
rect 13850 55970 13870 56210
rect 13800 55890 13870 55970
rect 13438 55832 13638 55838
rect 13438 55830 13450 55832
rect 13128 55800 13450 55830
rect 13128 55798 13140 55800
rect 12940 55792 13140 55798
rect 13438 55798 13450 55800
rect 13626 55798 13638 55832
rect 13438 55792 13638 55798
rect 13670 55800 13750 55820
rect 12902 55754 12910 55788
rect 12900 55740 12910 55754
rect 12830 55720 12910 55740
rect 12940 55744 13140 55750
rect 12940 55710 12952 55744
rect 13128 55740 13140 55744
rect 13438 55744 13638 55750
rect 13438 55740 13450 55744
rect 13128 55730 13450 55740
rect 13128 55710 13260 55730
rect 12940 55704 13140 55710
rect 13250 55670 13260 55710
rect 13320 55710 13450 55730
rect 13626 55710 13638 55744
rect 13670 55740 13680 55800
rect 13740 55740 13750 55800
rect 13670 55720 13750 55740
rect 13320 55670 13330 55710
rect 13438 55704 13638 55710
rect 13250 55660 13330 55670
rect 12720 54500 12790 55650
rect 12720 54240 12740 54500
rect 12780 54240 12790 54500
rect 13800 55650 13810 55890
rect 13850 55650 13870 55890
rect 13800 54500 13870 55650
rect 13250 54470 13330 54480
rect 12940 54432 13140 54438
rect 12830 54400 12910 54420
rect 12830 54340 12840 54400
rect 12900 54388 12910 54400
rect 12940 54398 12952 54432
rect 13128 54430 13140 54432
rect 13250 54430 13260 54470
rect 13128 54410 13260 54430
rect 13320 54430 13330 54470
rect 13438 54432 13638 54438
rect 13438 54430 13450 54432
rect 13320 54410 13450 54430
rect 13128 54400 13450 54410
rect 13128 54398 13140 54400
rect 12940 54392 13140 54398
rect 13438 54398 13450 54400
rect 13626 54398 13638 54432
rect 13438 54392 13638 54398
rect 13670 54400 13750 54420
rect 12902 54354 12910 54388
rect 12900 54340 12910 54354
rect 12830 54320 12910 54340
rect 12940 54344 13140 54350
rect 12940 54310 12952 54344
rect 13128 54340 13140 54344
rect 13438 54344 13638 54350
rect 13438 54340 13450 54344
rect 13128 54310 13450 54340
rect 13626 54310 13638 54344
rect 13670 54340 13680 54400
rect 13740 54340 13750 54400
rect 13670 54320 13750 54340
rect 12940 54304 13140 54310
rect 12720 54180 12790 54240
rect 12720 53940 12740 54180
rect 12780 53940 12790 54180
rect 13250 54300 13330 54310
rect 13438 54304 13638 54310
rect 13250 54240 13260 54300
rect 13320 54240 13330 54300
rect 13250 54190 13330 54240
rect 13250 54130 13260 54190
rect 13320 54130 13330 54190
rect 12940 54122 13140 54128
rect 12830 54090 12910 54110
rect 12830 54030 12840 54090
rect 12900 54078 12910 54090
rect 12940 54088 12952 54122
rect 13128 54120 13140 54122
rect 13250 54120 13330 54130
rect 13800 54260 13810 54500
rect 13850 54260 13870 54500
rect 13800 54180 13870 54260
rect 13438 54122 13638 54128
rect 13438 54120 13450 54122
rect 13128 54090 13450 54120
rect 13128 54088 13140 54090
rect 12940 54082 13140 54088
rect 13438 54088 13450 54090
rect 13626 54088 13638 54122
rect 13438 54082 13638 54088
rect 13670 54090 13750 54110
rect 12902 54044 12910 54078
rect 12900 54030 12910 54044
rect 12830 54010 12910 54030
rect 12940 54034 13140 54040
rect 12940 54000 12952 54034
rect 13128 54030 13140 54034
rect 13438 54034 13638 54040
rect 13438 54030 13450 54034
rect 13128 54020 13450 54030
rect 13128 54000 13260 54020
rect 12940 53994 13140 54000
rect 13250 53960 13260 54000
rect 13320 54000 13450 54020
rect 13626 54000 13638 54034
rect 13670 54030 13680 54090
rect 13740 54030 13750 54090
rect 13670 54010 13750 54030
rect 13320 53960 13330 54000
rect 13438 53994 13638 54000
rect 13250 53950 13330 53960
rect 12720 52790 12790 53940
rect 12720 52530 12740 52790
rect 12780 52530 12790 52790
rect 13800 53940 13810 54180
rect 13850 53940 13870 54180
rect 13800 52790 13870 53940
rect 13250 52760 13330 52770
rect 12940 52722 13140 52728
rect 12830 52690 12910 52710
rect 12830 52630 12840 52690
rect 12900 52678 12910 52690
rect 12940 52688 12952 52722
rect 13128 52720 13140 52722
rect 13250 52720 13260 52760
rect 13128 52700 13260 52720
rect 13320 52720 13330 52760
rect 13438 52722 13638 52728
rect 13438 52720 13450 52722
rect 13320 52700 13450 52720
rect 13128 52690 13450 52700
rect 13128 52688 13140 52690
rect 12940 52682 13140 52688
rect 13438 52688 13450 52690
rect 13626 52688 13638 52722
rect 13438 52682 13638 52688
rect 13670 52690 13750 52710
rect 12902 52644 12910 52678
rect 12900 52630 12910 52644
rect 12830 52610 12910 52630
rect 12940 52634 13140 52640
rect 12940 52600 12952 52634
rect 13128 52630 13140 52634
rect 13438 52634 13638 52640
rect 13438 52630 13450 52634
rect 13128 52600 13450 52630
rect 13626 52600 13638 52634
rect 13670 52630 13680 52690
rect 13740 52630 13750 52690
rect 13670 52610 13750 52630
rect 12940 52594 13140 52600
rect 12720 52470 12790 52530
rect 12720 52230 12740 52470
rect 12780 52230 12790 52470
rect 13250 52590 13330 52600
rect 13438 52594 13638 52600
rect 13250 52530 13260 52590
rect 13320 52530 13330 52590
rect 13250 52480 13330 52530
rect 13250 52420 13260 52480
rect 13320 52420 13330 52480
rect 12940 52412 13140 52418
rect 12830 52380 12910 52400
rect 12830 52320 12840 52380
rect 12900 52368 12910 52380
rect 12940 52378 12952 52412
rect 13128 52410 13140 52412
rect 13250 52410 13330 52420
rect 13800 52550 13810 52790
rect 13850 52550 13870 52790
rect 13800 52470 13870 52550
rect 13438 52412 13638 52418
rect 13438 52410 13450 52412
rect 13128 52380 13450 52410
rect 13128 52378 13140 52380
rect 12940 52372 13140 52378
rect 13438 52378 13450 52380
rect 13626 52378 13638 52412
rect 13438 52372 13638 52378
rect 13670 52380 13750 52400
rect 12902 52334 12910 52368
rect 12900 52320 12910 52334
rect 12830 52300 12910 52320
rect 12940 52324 13140 52330
rect 12940 52290 12952 52324
rect 13128 52320 13140 52324
rect 13438 52324 13638 52330
rect 13438 52320 13450 52324
rect 13128 52310 13450 52320
rect 13128 52290 13260 52310
rect 12940 52284 13140 52290
rect 13250 52250 13260 52290
rect 13320 52290 13450 52310
rect 13626 52290 13638 52324
rect 13670 52320 13680 52380
rect 13740 52320 13750 52380
rect 13670 52300 13750 52320
rect 13320 52250 13330 52290
rect 13438 52284 13638 52290
rect 13250 52240 13330 52250
rect 12720 51080 12790 52230
rect 12720 50820 12740 51080
rect 12780 50820 12790 51080
rect 13800 52230 13810 52470
rect 13850 52230 13870 52470
rect 13800 51080 13870 52230
rect 13250 51050 13330 51060
rect 12940 51012 13140 51018
rect 12830 50980 12910 51000
rect 12830 50920 12840 50980
rect 12900 50968 12910 50980
rect 12940 50978 12952 51012
rect 13128 51010 13140 51012
rect 13250 51010 13260 51050
rect 13128 50990 13260 51010
rect 13320 51010 13330 51050
rect 13438 51012 13638 51018
rect 13438 51010 13450 51012
rect 13320 50990 13450 51010
rect 13128 50980 13450 50990
rect 13128 50978 13140 50980
rect 12940 50972 13140 50978
rect 13438 50978 13450 50980
rect 13626 50978 13638 51012
rect 13438 50972 13638 50978
rect 13670 50980 13750 51000
rect 12902 50934 12910 50968
rect 12900 50920 12910 50934
rect 12830 50900 12910 50920
rect 12940 50924 13140 50930
rect 12940 50890 12952 50924
rect 13128 50920 13140 50924
rect 13438 50924 13638 50930
rect 13438 50920 13450 50924
rect 13128 50890 13450 50920
rect 13626 50890 13638 50924
rect 13670 50920 13680 50980
rect 13740 50920 13750 50980
rect 13670 50900 13750 50920
rect 12940 50884 13140 50890
rect 12720 50760 12790 50820
rect 12720 50520 12740 50760
rect 12780 50520 12790 50760
rect 13250 50880 13330 50890
rect 13438 50884 13638 50890
rect 13250 50820 13260 50880
rect 13320 50820 13330 50880
rect 13250 50770 13330 50820
rect 13250 50710 13260 50770
rect 13320 50710 13330 50770
rect 12940 50702 13140 50708
rect 12830 50670 12910 50690
rect 12830 50610 12840 50670
rect 12900 50658 12910 50670
rect 12940 50668 12952 50702
rect 13128 50700 13140 50702
rect 13250 50700 13330 50710
rect 13800 50840 13810 51080
rect 13850 50840 13870 51080
rect 13800 50760 13870 50840
rect 13438 50702 13638 50708
rect 13438 50700 13450 50702
rect 13128 50670 13450 50700
rect 13128 50668 13140 50670
rect 12940 50662 13140 50668
rect 13438 50668 13450 50670
rect 13626 50668 13638 50702
rect 13438 50662 13638 50668
rect 13670 50670 13750 50690
rect 12902 50624 12910 50658
rect 12900 50610 12910 50624
rect 12830 50590 12910 50610
rect 12940 50614 13140 50620
rect 12940 50580 12952 50614
rect 13128 50610 13140 50614
rect 13438 50614 13638 50620
rect 13438 50610 13450 50614
rect 13128 50600 13450 50610
rect 13128 50580 13260 50600
rect 12940 50574 13140 50580
rect 13250 50540 13260 50580
rect 13320 50580 13450 50600
rect 13626 50580 13638 50614
rect 13670 50610 13680 50670
rect 13740 50610 13750 50670
rect 13670 50590 13750 50610
rect 13320 50540 13330 50580
rect 13438 50574 13638 50580
rect 13250 50530 13330 50540
rect 12720 49370 12790 50520
rect 12720 49110 12740 49370
rect 12780 49110 12790 49370
rect 13800 50520 13810 50760
rect 13850 50520 13870 50760
rect 13800 49370 13870 50520
rect 13250 49340 13330 49350
rect 12940 49302 13140 49308
rect 12830 49270 12910 49290
rect 12830 49210 12840 49270
rect 12900 49258 12910 49270
rect 12940 49268 12952 49302
rect 13128 49300 13140 49302
rect 13250 49300 13260 49340
rect 13128 49280 13260 49300
rect 13320 49300 13330 49340
rect 13438 49302 13638 49308
rect 13438 49300 13450 49302
rect 13320 49280 13450 49300
rect 13128 49270 13450 49280
rect 13128 49268 13140 49270
rect 12940 49262 13140 49268
rect 13438 49268 13450 49270
rect 13626 49268 13638 49302
rect 13438 49262 13638 49268
rect 13670 49270 13750 49290
rect 12902 49224 12910 49258
rect 12900 49210 12910 49224
rect 12830 49190 12910 49210
rect 12940 49214 13140 49220
rect 12940 49180 12952 49214
rect 13128 49210 13140 49214
rect 13438 49214 13638 49220
rect 13438 49210 13450 49214
rect 13128 49180 13450 49210
rect 13626 49180 13638 49214
rect 13670 49210 13680 49270
rect 13740 49210 13750 49270
rect 13670 49190 13750 49210
rect 12940 49174 13140 49180
rect 12720 49050 12790 49110
rect 12720 48810 12740 49050
rect 12780 48810 12790 49050
rect 13250 49170 13330 49180
rect 13438 49174 13638 49180
rect 13250 49110 13260 49170
rect 13320 49110 13330 49170
rect 13250 49060 13330 49110
rect 13250 49000 13260 49060
rect 13320 49000 13330 49060
rect 12940 48992 13140 48998
rect 12830 48960 12910 48980
rect 12830 48900 12840 48960
rect 12900 48948 12910 48960
rect 12940 48958 12952 48992
rect 13128 48990 13140 48992
rect 13250 48990 13330 49000
rect 13800 49130 13810 49370
rect 13850 49130 13870 49370
rect 13800 49050 13870 49130
rect 13438 48992 13638 48998
rect 13438 48990 13450 48992
rect 13128 48960 13450 48990
rect 13128 48958 13140 48960
rect 12940 48952 13140 48958
rect 13438 48958 13450 48960
rect 13626 48958 13638 48992
rect 13438 48952 13638 48958
rect 13670 48960 13750 48980
rect 12902 48914 12910 48948
rect 12900 48900 12910 48914
rect 12830 48880 12910 48900
rect 12940 48904 13140 48910
rect 12940 48870 12952 48904
rect 13128 48900 13140 48904
rect 13438 48904 13638 48910
rect 13438 48900 13450 48904
rect 13128 48890 13450 48900
rect 13128 48870 13260 48890
rect 12940 48864 13140 48870
rect 13250 48830 13260 48870
rect 13320 48870 13450 48890
rect 13626 48870 13638 48904
rect 13670 48900 13680 48960
rect 13740 48900 13750 48960
rect 13670 48880 13750 48900
rect 13320 48830 13330 48870
rect 13438 48864 13638 48870
rect 13250 48820 13330 48830
rect 12720 47660 12790 48810
rect 12720 47400 12740 47660
rect 12780 47400 12790 47660
rect 13800 48810 13810 49050
rect 13850 48810 13870 49050
rect 13800 47660 13870 48810
rect 13250 47630 13330 47640
rect 12940 47592 13140 47598
rect 12830 47560 12910 47580
rect 12830 47500 12840 47560
rect 12900 47548 12910 47560
rect 12940 47558 12952 47592
rect 13128 47590 13140 47592
rect 13250 47590 13260 47630
rect 13128 47570 13260 47590
rect 13320 47590 13330 47630
rect 13438 47592 13638 47598
rect 13438 47590 13450 47592
rect 13320 47570 13450 47590
rect 13128 47560 13450 47570
rect 13128 47558 13140 47560
rect 12940 47552 13140 47558
rect 13438 47558 13450 47560
rect 13626 47558 13638 47592
rect 13438 47552 13638 47558
rect 13670 47560 13750 47580
rect 12902 47514 12910 47548
rect 12900 47500 12910 47514
rect 12830 47480 12910 47500
rect 12940 47504 13140 47510
rect 12940 47470 12952 47504
rect 13128 47500 13140 47504
rect 13438 47504 13638 47510
rect 13438 47500 13450 47504
rect 13128 47470 13450 47500
rect 13626 47470 13638 47504
rect 13670 47500 13680 47560
rect 13740 47500 13750 47560
rect 13670 47480 13750 47500
rect 12940 47464 13140 47470
rect 12720 47340 12790 47400
rect 12720 47100 12740 47340
rect 12780 47100 12790 47340
rect 13250 47460 13330 47470
rect 13438 47464 13638 47470
rect 13250 47400 13260 47460
rect 13320 47400 13330 47460
rect 13250 47350 13330 47400
rect 13250 47290 13260 47350
rect 13320 47290 13330 47350
rect 12940 47282 13140 47288
rect 12830 47250 12910 47270
rect 12830 47190 12840 47250
rect 12900 47238 12910 47250
rect 12940 47248 12952 47282
rect 13128 47280 13140 47282
rect 13250 47280 13330 47290
rect 13800 47420 13810 47660
rect 13850 47420 13870 47660
rect 13800 47340 13870 47420
rect 13438 47282 13638 47288
rect 13438 47280 13450 47282
rect 13128 47250 13450 47280
rect 13128 47248 13140 47250
rect 12940 47242 13140 47248
rect 13438 47248 13450 47250
rect 13626 47248 13638 47282
rect 13438 47242 13638 47248
rect 13670 47250 13750 47270
rect 12902 47204 12910 47238
rect 12900 47190 12910 47204
rect 12830 47170 12910 47190
rect 12940 47194 13140 47200
rect 12940 47160 12952 47194
rect 13128 47190 13140 47194
rect 13438 47194 13638 47200
rect 13438 47190 13450 47194
rect 13128 47180 13450 47190
rect 13128 47160 13260 47180
rect 12940 47154 13140 47160
rect 13250 47120 13260 47160
rect 13320 47160 13450 47180
rect 13626 47160 13638 47194
rect 13670 47190 13680 47250
rect 13740 47190 13750 47250
rect 13670 47170 13750 47190
rect 13320 47120 13330 47160
rect 13438 47154 13638 47160
rect 13250 47110 13330 47120
rect 12720 45950 12790 47100
rect 12720 45690 12740 45950
rect 12780 45690 12790 45950
rect 13800 47100 13810 47340
rect 13850 47100 13870 47340
rect 13800 45950 13870 47100
rect 13250 45920 13330 45930
rect 12940 45882 13140 45888
rect 12830 45850 12910 45870
rect 12830 45790 12840 45850
rect 12900 45838 12910 45850
rect 12940 45848 12952 45882
rect 13128 45880 13140 45882
rect 13250 45880 13260 45920
rect 13128 45860 13260 45880
rect 13320 45880 13330 45920
rect 13438 45882 13638 45888
rect 13438 45880 13450 45882
rect 13320 45860 13450 45880
rect 13128 45850 13450 45860
rect 13128 45848 13140 45850
rect 12940 45842 13140 45848
rect 13438 45848 13450 45850
rect 13626 45848 13638 45882
rect 13438 45842 13638 45848
rect 13670 45850 13750 45870
rect 12902 45804 12910 45838
rect 12900 45790 12910 45804
rect 12830 45770 12910 45790
rect 12940 45794 13140 45800
rect 12940 45760 12952 45794
rect 13128 45790 13140 45794
rect 13438 45794 13638 45800
rect 13438 45790 13450 45794
rect 13128 45760 13450 45790
rect 13626 45760 13638 45794
rect 13670 45790 13680 45850
rect 13740 45790 13750 45850
rect 13670 45770 13750 45790
rect 12940 45754 13140 45760
rect 12720 45630 12790 45690
rect 12720 45390 12740 45630
rect 12780 45390 12790 45630
rect 13250 45750 13330 45760
rect 13438 45754 13638 45760
rect 13250 45690 13260 45750
rect 13320 45690 13330 45750
rect 13250 45640 13330 45690
rect 13250 45580 13260 45640
rect 13320 45580 13330 45640
rect 12940 45572 13140 45578
rect 12830 45540 12910 45560
rect 12830 45480 12840 45540
rect 12900 45528 12910 45540
rect 12940 45538 12952 45572
rect 13128 45570 13140 45572
rect 13250 45570 13330 45580
rect 13800 45710 13810 45950
rect 13850 45710 13870 45950
rect 13800 45630 13870 45710
rect 13438 45572 13638 45578
rect 13438 45570 13450 45572
rect 13128 45540 13450 45570
rect 13128 45538 13140 45540
rect 12940 45532 13140 45538
rect 13438 45538 13450 45540
rect 13626 45538 13638 45572
rect 13438 45532 13638 45538
rect 13670 45540 13750 45560
rect 12902 45494 12910 45528
rect 12900 45480 12910 45494
rect 12830 45460 12910 45480
rect 12940 45484 13140 45490
rect 12940 45450 12952 45484
rect 13128 45480 13140 45484
rect 13438 45484 13638 45490
rect 13438 45480 13450 45484
rect 13128 45470 13450 45480
rect 13128 45450 13260 45470
rect 12940 45444 13140 45450
rect 13250 45410 13260 45450
rect 13320 45450 13450 45470
rect 13626 45450 13638 45484
rect 13670 45480 13680 45540
rect 13740 45480 13750 45540
rect 13670 45460 13750 45480
rect 13320 45410 13330 45450
rect 13438 45444 13638 45450
rect 13250 45400 13330 45410
rect 12720 44240 12790 45390
rect 12720 43980 12740 44240
rect 12780 43980 12790 44240
rect 13800 45390 13810 45630
rect 13850 45390 13870 45630
rect 13800 44240 13870 45390
rect 13250 44210 13330 44220
rect 12940 44172 13140 44178
rect 12830 44140 12910 44160
rect 12830 44080 12840 44140
rect 12900 44128 12910 44140
rect 12940 44138 12952 44172
rect 13128 44170 13140 44172
rect 13250 44170 13260 44210
rect 13128 44150 13260 44170
rect 13320 44170 13330 44210
rect 13438 44172 13638 44178
rect 13438 44170 13450 44172
rect 13320 44150 13450 44170
rect 13128 44140 13450 44150
rect 13128 44138 13140 44140
rect 12940 44132 13140 44138
rect 13438 44138 13450 44140
rect 13626 44138 13638 44172
rect 13438 44132 13638 44138
rect 13670 44140 13750 44160
rect 12902 44094 12910 44128
rect 12900 44080 12910 44094
rect 12830 44060 12910 44080
rect 12940 44084 13140 44090
rect 12940 44050 12952 44084
rect 13128 44080 13140 44084
rect 13438 44084 13638 44090
rect 13438 44080 13450 44084
rect 13128 44050 13450 44080
rect 13626 44050 13638 44084
rect 13670 44080 13680 44140
rect 13740 44080 13750 44140
rect 13670 44060 13750 44080
rect 12940 44044 13140 44050
rect 12720 43920 12790 43980
rect 12720 43680 12740 43920
rect 12780 43680 12790 43920
rect 13250 44040 13330 44050
rect 13438 44044 13638 44050
rect 13250 43980 13260 44040
rect 13320 43980 13330 44040
rect 13250 43930 13330 43980
rect 13250 43870 13260 43930
rect 13320 43870 13330 43930
rect 12940 43862 13140 43868
rect 12830 43830 12910 43850
rect 12830 43770 12840 43830
rect 12900 43818 12910 43830
rect 12940 43828 12952 43862
rect 13128 43860 13140 43862
rect 13250 43860 13330 43870
rect 13800 44000 13810 44240
rect 13850 44000 13870 44240
rect 13800 43920 13870 44000
rect 13438 43862 13638 43868
rect 13438 43860 13450 43862
rect 13128 43830 13450 43860
rect 13128 43828 13140 43830
rect 12940 43822 13140 43828
rect 13438 43828 13450 43830
rect 13626 43828 13638 43862
rect 13438 43822 13638 43828
rect 13670 43830 13750 43850
rect 12902 43784 12910 43818
rect 12900 43770 12910 43784
rect 12830 43750 12910 43770
rect 12940 43774 13140 43780
rect 12940 43740 12952 43774
rect 13128 43770 13140 43774
rect 13438 43774 13638 43780
rect 13438 43770 13450 43774
rect 13128 43760 13450 43770
rect 13128 43740 13260 43760
rect 12940 43734 13140 43740
rect 13250 43700 13260 43740
rect 13320 43740 13450 43760
rect 13626 43740 13638 43774
rect 13670 43770 13680 43830
rect 13740 43770 13750 43830
rect 13670 43750 13750 43770
rect 13320 43700 13330 43740
rect 13438 43734 13638 43740
rect 13250 43690 13330 43700
rect 12720 42530 12790 43680
rect 12720 42270 12740 42530
rect 12780 42270 12790 42530
rect 13800 43680 13810 43920
rect 13850 43680 13870 43920
rect 13800 42530 13870 43680
rect 13250 42500 13330 42510
rect 12940 42462 13140 42468
rect 12830 42430 12910 42450
rect 12830 42370 12840 42430
rect 12900 42418 12910 42430
rect 12940 42428 12952 42462
rect 13128 42460 13140 42462
rect 13250 42460 13260 42500
rect 13128 42440 13260 42460
rect 13320 42460 13330 42500
rect 13438 42462 13638 42468
rect 13438 42460 13450 42462
rect 13320 42440 13450 42460
rect 13128 42430 13450 42440
rect 13128 42428 13140 42430
rect 12940 42422 13140 42428
rect 13438 42428 13450 42430
rect 13626 42428 13638 42462
rect 13438 42422 13638 42428
rect 13670 42430 13750 42450
rect 12902 42384 12910 42418
rect 12900 42370 12910 42384
rect 12830 42350 12910 42370
rect 12940 42374 13140 42380
rect 12940 42340 12952 42374
rect 13128 42370 13140 42374
rect 13438 42374 13638 42380
rect 13438 42370 13450 42374
rect 13128 42340 13450 42370
rect 13626 42340 13638 42374
rect 13670 42370 13680 42430
rect 13740 42370 13750 42430
rect 13670 42350 13750 42370
rect 12940 42334 13140 42340
rect 12720 42210 12790 42270
rect 12720 41970 12740 42210
rect 12780 41970 12790 42210
rect 13250 42330 13330 42340
rect 13438 42334 13638 42340
rect 13250 42270 13260 42330
rect 13320 42270 13330 42330
rect 13250 42220 13330 42270
rect 13250 42160 13260 42220
rect 13320 42160 13330 42220
rect 12940 42152 13140 42158
rect 12830 42120 12910 42140
rect 12830 42060 12840 42120
rect 12900 42108 12910 42120
rect 12940 42118 12952 42152
rect 13128 42150 13140 42152
rect 13250 42150 13330 42160
rect 13800 42290 13810 42530
rect 13850 42290 13870 42530
rect 13800 42210 13870 42290
rect 13438 42152 13638 42158
rect 13438 42150 13450 42152
rect 13128 42120 13450 42150
rect 13128 42118 13140 42120
rect 12940 42112 13140 42118
rect 13438 42118 13450 42120
rect 13626 42118 13638 42152
rect 13438 42112 13638 42118
rect 13670 42120 13750 42140
rect 12902 42074 12910 42108
rect 12900 42060 12910 42074
rect 12830 42040 12910 42060
rect 12940 42064 13140 42070
rect 12940 42030 12952 42064
rect 13128 42060 13140 42064
rect 13438 42064 13638 42070
rect 13438 42060 13450 42064
rect 13128 42050 13450 42060
rect 13128 42030 13260 42050
rect 12940 42024 13140 42030
rect 13250 41990 13260 42030
rect 13320 42030 13450 42050
rect 13626 42030 13638 42064
rect 13670 42060 13680 42120
rect 13740 42060 13750 42120
rect 13670 42040 13750 42060
rect 13320 41990 13330 42030
rect 13438 42024 13638 42030
rect 13250 41980 13330 41990
rect 12720 40820 12790 41970
rect 12720 40560 12740 40820
rect 12780 40560 12790 40820
rect 13800 41970 13810 42210
rect 13850 41970 13870 42210
rect 13800 40820 13870 41970
rect 13250 40790 13330 40800
rect 12940 40752 13140 40758
rect 12830 40720 12910 40740
rect 12830 40660 12840 40720
rect 12900 40708 12910 40720
rect 12940 40718 12952 40752
rect 13128 40750 13140 40752
rect 13250 40750 13260 40790
rect 13128 40730 13260 40750
rect 13320 40750 13330 40790
rect 13438 40752 13638 40758
rect 13438 40750 13450 40752
rect 13320 40730 13450 40750
rect 13128 40720 13450 40730
rect 13128 40718 13140 40720
rect 12940 40712 13140 40718
rect 13438 40718 13450 40720
rect 13626 40718 13638 40752
rect 13438 40712 13638 40718
rect 13670 40720 13750 40740
rect 12902 40674 12910 40708
rect 12900 40660 12910 40674
rect 12830 40640 12910 40660
rect 12940 40664 13140 40670
rect 12940 40630 12952 40664
rect 13128 40660 13140 40664
rect 13438 40664 13638 40670
rect 13438 40660 13450 40664
rect 13128 40630 13450 40660
rect 13626 40630 13638 40664
rect 13670 40660 13680 40720
rect 13740 40660 13750 40720
rect 13670 40640 13750 40660
rect 12940 40624 13140 40630
rect 12720 40500 12790 40560
rect 12720 40260 12740 40500
rect 12780 40260 12790 40500
rect 13250 40620 13330 40630
rect 13438 40624 13638 40630
rect 13250 40560 13260 40620
rect 13320 40560 13330 40620
rect 13250 40510 13330 40560
rect 13250 40450 13260 40510
rect 13320 40450 13330 40510
rect 12940 40442 13140 40448
rect 12830 40410 12910 40430
rect 12830 40350 12840 40410
rect 12900 40398 12910 40410
rect 12940 40408 12952 40442
rect 13128 40440 13140 40442
rect 13250 40440 13330 40450
rect 13800 40580 13810 40820
rect 13850 40580 13870 40820
rect 13800 40500 13870 40580
rect 13438 40442 13638 40448
rect 13438 40440 13450 40442
rect 13128 40410 13450 40440
rect 13128 40408 13140 40410
rect 12940 40402 13140 40408
rect 13438 40408 13450 40410
rect 13626 40408 13638 40442
rect 13438 40402 13638 40408
rect 13670 40410 13750 40430
rect 12902 40364 12910 40398
rect 12900 40350 12910 40364
rect 12830 40330 12910 40350
rect 12940 40354 13140 40360
rect 12940 40320 12952 40354
rect 13128 40350 13140 40354
rect 13438 40354 13638 40360
rect 13438 40350 13450 40354
rect 13128 40340 13450 40350
rect 13128 40320 13260 40340
rect 12940 40314 13140 40320
rect 13250 40280 13260 40320
rect 13320 40320 13450 40340
rect 13626 40320 13638 40354
rect 13670 40350 13680 40410
rect 13740 40350 13750 40410
rect 13670 40330 13750 40350
rect 13320 40280 13330 40320
rect 13438 40314 13638 40320
rect 13250 40270 13330 40280
rect 12720 39690 12790 40260
rect 13800 40260 13810 40500
rect 13850 40260 13870 40500
rect 13800 39690 13870 40260
rect 12720 39680 12800 39690
rect 12720 39620 12730 39680
rect 12790 39620 12800 39680
rect 13790 39680 13870 39690
rect 13790 39620 13800 39680
rect 13860 39620 13870 39680
rect 13790 39610 13870 39620
rect 13900 66480 13930 67050
rect 13900 66470 13960 66480
rect 13900 66400 13960 66410
rect 13900 64770 13930 66400
rect 13990 65950 14020 67050
rect 13960 65940 14020 65950
rect 13960 65870 14020 65880
rect 13900 64760 13960 64770
rect 13900 64690 13960 64700
rect 13900 63060 13930 64690
rect 13990 64240 14020 65870
rect 13960 64230 14020 64240
rect 13960 64160 14020 64170
rect 13900 63050 13960 63060
rect 13900 62980 13960 62990
rect 13900 61350 13930 62980
rect 13990 62530 14020 64160
rect 13960 62520 14020 62530
rect 13960 62450 14020 62460
rect 13900 61340 13960 61350
rect 13900 61270 13960 61280
rect 13900 59640 13930 61270
rect 13990 60820 14020 62450
rect 13960 60810 14020 60820
rect 13960 60740 14020 60750
rect 13900 59630 13960 59640
rect 13900 59560 13960 59570
rect 13900 57930 13930 59560
rect 13990 59110 14020 60740
rect 13960 59100 14020 59110
rect 13960 59030 14020 59040
rect 13900 57920 13960 57930
rect 13900 57850 13960 57860
rect 13900 56220 13930 57850
rect 13990 57400 14020 59030
rect 13960 57390 14020 57400
rect 13960 57320 14020 57330
rect 13900 56210 13960 56220
rect 13900 56140 13960 56150
rect 13900 54510 13930 56140
rect 13990 55690 14020 57320
rect 13960 55680 14020 55690
rect 13960 55610 14020 55620
rect 13900 54500 13960 54510
rect 13900 54430 13960 54440
rect 13900 52800 13930 54430
rect 13990 53980 14020 55610
rect 13960 53970 14020 53980
rect 13960 53900 14020 53910
rect 13900 52790 13960 52800
rect 13900 52720 13960 52730
rect 13900 51090 13930 52720
rect 13990 52270 14020 53900
rect 13960 52260 14020 52270
rect 13960 52190 14020 52200
rect 13900 51080 13960 51090
rect 13900 51010 13960 51020
rect 13900 49380 13930 51010
rect 13990 50560 14020 52190
rect 13960 50550 14020 50560
rect 13960 50480 14020 50490
rect 13900 49370 13960 49380
rect 13900 49300 13960 49310
rect 13900 47670 13930 49300
rect 13990 48850 14020 50480
rect 13960 48840 14020 48850
rect 13960 48770 14020 48780
rect 13900 47660 13960 47670
rect 13900 47590 13960 47600
rect 13900 45960 13930 47590
rect 13990 47140 14020 48770
rect 13960 47130 14020 47140
rect 13960 47060 14020 47070
rect 13900 45950 13960 45960
rect 13900 45880 13960 45890
rect 13900 44250 13930 45880
rect 13990 45430 14020 47060
rect 13960 45420 14020 45430
rect 13960 45350 14020 45360
rect 13900 44240 13960 44250
rect 13900 44170 13960 44180
rect 13900 42540 13930 44170
rect 13990 43720 14020 45350
rect 13960 43710 14020 43720
rect 13960 43640 14020 43650
rect 13900 42530 13960 42540
rect 13900 42460 13960 42470
rect 13900 40830 13930 42460
rect 13990 42010 14020 43640
rect 13960 42000 14020 42010
rect 13960 41930 14020 41940
rect 13900 40820 13960 40830
rect 13900 40750 13960 40760
rect 12250 39220 12310 39230
rect 12430 39230 12690 39240
rect 9260 39160 9320 39170
rect 12490 39210 12690 39230
rect 12430 39160 12490 39170
rect 13900 38840 13930 40750
rect 13990 40300 14020 41930
rect 13960 40290 14020 40300
rect 13960 40220 14020 40230
rect 13990 39690 14020 40220
rect 13960 39680 14020 39690
rect 13960 39610 14020 39620
rect 14050 66390 14080 67050
rect 14050 66380 14110 66390
rect 14050 66310 14110 66320
rect 14050 64680 14080 66310
rect 14050 64670 14110 64680
rect 14050 64600 14110 64610
rect 14050 62970 14080 64600
rect 14050 62960 14110 62970
rect 14050 62890 14110 62900
rect 14050 61260 14080 62890
rect 14050 61250 14110 61260
rect 14050 61180 14110 61190
rect 14050 45870 14080 61180
rect 14170 59550 14200 67050
rect 14170 59540 14230 59550
rect 14170 59470 14230 59480
rect 14170 57840 14200 59470
rect 14170 57830 14230 57840
rect 14170 57760 14230 57770
rect 14170 56130 14200 57760
rect 14170 56120 14230 56130
rect 14170 56050 14230 56060
rect 14170 54420 14200 56050
rect 14170 54410 14230 54420
rect 14170 54340 14230 54350
rect 14170 52710 14200 54340
rect 14170 52700 14230 52710
rect 14170 52630 14230 52640
rect 14170 51000 14200 52630
rect 14170 50990 14230 51000
rect 14170 50920 14230 50930
rect 14170 49290 14200 50920
rect 14170 49280 14230 49290
rect 14170 49210 14230 49220
rect 14170 47580 14200 49210
rect 14170 47570 14230 47580
rect 14170 47500 14230 47510
rect 14050 45860 14110 45870
rect 14050 45790 14110 45800
rect 14050 44160 14080 45790
rect 14050 44150 14110 44160
rect 14050 44080 14110 44090
rect 14050 42450 14080 44080
rect 14050 42440 14110 42450
rect 14050 42370 14110 42380
rect 14050 40740 14080 42370
rect 14050 40730 14110 40740
rect 14050 40660 14110 40670
rect 14050 39240 14080 40660
rect 14170 39300 14200 47500
rect 14290 39690 14320 67050
rect 14410 39690 14440 67050
rect 14530 39690 14560 67050
rect 14650 39690 14680 67050
rect 14770 39690 14800 67050
rect 16930 39690 16960 67050
rect 17050 39690 17080 67050
rect 17170 39690 17200 67050
rect 17290 39690 17320 67050
rect 17410 39690 17440 67050
rect 17530 59550 17560 67050
rect 17650 66390 17680 67050
rect 17620 66380 17680 66390
rect 17620 66310 17680 66320
rect 17650 64680 17680 66310
rect 17620 64670 17680 64680
rect 17620 64600 17680 64610
rect 17650 62970 17680 64600
rect 17620 62960 17680 62970
rect 17620 62890 17680 62900
rect 17650 61260 17680 62890
rect 17620 61250 17680 61260
rect 17620 61180 17680 61190
rect 17500 59540 17560 59550
rect 17500 59470 17560 59480
rect 17530 57840 17560 59470
rect 17500 57830 17560 57840
rect 17500 57760 17560 57770
rect 17530 56130 17560 57760
rect 17500 56120 17560 56130
rect 17500 56050 17560 56060
rect 17530 54420 17560 56050
rect 17500 54410 17560 54420
rect 17500 54340 17560 54350
rect 17530 52710 17560 54340
rect 17500 52700 17560 52710
rect 17500 52630 17560 52640
rect 17530 51000 17560 52630
rect 17500 50990 17560 51000
rect 17500 50920 17560 50930
rect 17530 49290 17560 50920
rect 17500 49280 17560 49290
rect 17500 49210 17560 49220
rect 17530 47580 17560 49210
rect 17500 47570 17560 47580
rect 17500 47500 17560 47510
rect 17530 39300 17560 47500
rect 17650 45870 17680 61180
rect 17620 45860 17680 45870
rect 17620 45790 17680 45800
rect 17650 44160 17680 45790
rect 17620 44150 17680 44160
rect 17620 44080 17680 44090
rect 17650 42450 17680 44080
rect 17620 42440 17680 42450
rect 17620 42370 17680 42380
rect 17650 40740 17680 42370
rect 17620 40730 17680 40740
rect 17620 40660 17680 40670
rect 14170 39290 14490 39300
rect 14170 39270 14430 39290
rect 14050 39230 14310 39240
rect 14050 39210 14250 39230
rect 14430 39220 14490 39230
rect 17240 39290 17560 39300
rect 17300 39270 17560 39290
rect 17650 39240 17680 40660
rect 17710 66470 17780 67050
rect 17710 66210 17730 66470
rect 17770 66210 17780 66470
rect 18790 66470 18860 67050
rect 18240 66440 18320 66450
rect 17930 66402 18130 66408
rect 17820 66370 17900 66390
rect 17820 66310 17830 66370
rect 17890 66358 17900 66370
rect 17930 66368 17942 66402
rect 18118 66400 18130 66402
rect 18240 66400 18250 66440
rect 18118 66380 18250 66400
rect 18310 66400 18320 66440
rect 18428 66402 18628 66408
rect 18428 66400 18440 66402
rect 18310 66380 18440 66400
rect 18118 66370 18440 66380
rect 18118 66368 18130 66370
rect 17930 66362 18130 66368
rect 18428 66368 18440 66370
rect 18616 66368 18628 66402
rect 18428 66362 18628 66368
rect 18660 66370 18740 66390
rect 17892 66324 17900 66358
rect 17890 66310 17900 66324
rect 17820 66290 17900 66310
rect 17930 66314 18130 66320
rect 17930 66280 17942 66314
rect 18118 66310 18130 66314
rect 18428 66314 18628 66320
rect 18428 66310 18440 66314
rect 18118 66280 18440 66310
rect 18616 66280 18628 66314
rect 18660 66310 18670 66370
rect 18730 66310 18740 66370
rect 18660 66290 18740 66310
rect 17930 66274 18130 66280
rect 17710 66150 17780 66210
rect 17710 65910 17730 66150
rect 17770 65910 17780 66150
rect 18240 66270 18320 66280
rect 18428 66274 18628 66280
rect 18240 66210 18250 66270
rect 18310 66210 18320 66270
rect 18240 66160 18320 66210
rect 18240 66100 18250 66160
rect 18310 66100 18320 66160
rect 17930 66092 18130 66098
rect 17820 66060 17900 66080
rect 17820 66000 17830 66060
rect 17890 66048 17900 66060
rect 17930 66058 17942 66092
rect 18118 66090 18130 66092
rect 18240 66090 18320 66100
rect 18790 66230 18800 66470
rect 18840 66230 18860 66470
rect 18790 66150 18860 66230
rect 18428 66092 18628 66098
rect 18428 66090 18440 66092
rect 18118 66060 18440 66090
rect 18118 66058 18130 66060
rect 17930 66052 18130 66058
rect 18428 66058 18440 66060
rect 18616 66058 18628 66092
rect 18428 66052 18628 66058
rect 18660 66060 18740 66080
rect 17892 66014 17900 66048
rect 17890 66000 17900 66014
rect 17820 65980 17900 66000
rect 17930 66004 18130 66010
rect 17930 65970 17942 66004
rect 18118 66000 18130 66004
rect 18428 66004 18628 66010
rect 18428 66000 18440 66004
rect 18118 65990 18440 66000
rect 18118 65970 18250 65990
rect 17930 65964 18130 65970
rect 18240 65930 18250 65970
rect 18310 65970 18440 65990
rect 18616 65970 18628 66004
rect 18660 66000 18670 66060
rect 18730 66000 18740 66060
rect 18660 65980 18740 66000
rect 18310 65930 18320 65970
rect 18428 65964 18628 65970
rect 18240 65920 18320 65930
rect 17710 64760 17780 65910
rect 17710 64500 17730 64760
rect 17770 64500 17780 64760
rect 18790 65910 18800 66150
rect 18840 65910 18860 66150
rect 18790 64760 18860 65910
rect 18240 64730 18320 64740
rect 17930 64692 18130 64698
rect 17820 64660 17900 64680
rect 17820 64600 17830 64660
rect 17890 64648 17900 64660
rect 17930 64658 17942 64692
rect 18118 64690 18130 64692
rect 18240 64690 18250 64730
rect 18118 64670 18250 64690
rect 18310 64690 18320 64730
rect 18428 64692 18628 64698
rect 18428 64690 18440 64692
rect 18310 64670 18440 64690
rect 18118 64660 18440 64670
rect 18118 64658 18130 64660
rect 17930 64652 18130 64658
rect 18428 64658 18440 64660
rect 18616 64658 18628 64692
rect 18428 64652 18628 64658
rect 18660 64660 18740 64680
rect 17892 64614 17900 64648
rect 17890 64600 17900 64614
rect 17820 64580 17900 64600
rect 17930 64604 18130 64610
rect 17930 64570 17942 64604
rect 18118 64600 18130 64604
rect 18428 64604 18628 64610
rect 18428 64600 18440 64604
rect 18118 64570 18440 64600
rect 18616 64570 18628 64604
rect 18660 64600 18670 64660
rect 18730 64600 18740 64660
rect 18660 64580 18740 64600
rect 17930 64564 18130 64570
rect 17710 64440 17780 64500
rect 17710 64200 17730 64440
rect 17770 64200 17780 64440
rect 18240 64560 18320 64570
rect 18428 64564 18628 64570
rect 18240 64500 18250 64560
rect 18310 64500 18320 64560
rect 18240 64450 18320 64500
rect 18240 64390 18250 64450
rect 18310 64390 18320 64450
rect 17930 64382 18130 64388
rect 17820 64350 17900 64370
rect 17820 64290 17830 64350
rect 17890 64338 17900 64350
rect 17930 64348 17942 64382
rect 18118 64380 18130 64382
rect 18240 64380 18320 64390
rect 18790 64520 18800 64760
rect 18840 64520 18860 64760
rect 18790 64440 18860 64520
rect 18428 64382 18628 64388
rect 18428 64380 18440 64382
rect 18118 64350 18440 64380
rect 18118 64348 18130 64350
rect 17930 64342 18130 64348
rect 18428 64348 18440 64350
rect 18616 64348 18628 64382
rect 18428 64342 18628 64348
rect 18660 64350 18740 64370
rect 17892 64304 17900 64338
rect 17890 64290 17900 64304
rect 17820 64270 17900 64290
rect 17930 64294 18130 64300
rect 17930 64260 17942 64294
rect 18118 64290 18130 64294
rect 18428 64294 18628 64300
rect 18428 64290 18440 64294
rect 18118 64280 18440 64290
rect 18118 64260 18250 64280
rect 17930 64254 18130 64260
rect 18240 64220 18250 64260
rect 18310 64260 18440 64280
rect 18616 64260 18628 64294
rect 18660 64290 18670 64350
rect 18730 64290 18740 64350
rect 18660 64270 18740 64290
rect 18310 64220 18320 64260
rect 18428 64254 18628 64260
rect 18240 64210 18320 64220
rect 17710 63050 17780 64200
rect 17710 62790 17730 63050
rect 17770 62790 17780 63050
rect 18790 64200 18800 64440
rect 18840 64200 18860 64440
rect 18790 63050 18860 64200
rect 18240 63020 18320 63030
rect 17930 62982 18130 62988
rect 17820 62950 17900 62970
rect 17820 62890 17830 62950
rect 17890 62938 17900 62950
rect 17930 62948 17942 62982
rect 18118 62980 18130 62982
rect 18240 62980 18250 63020
rect 18118 62960 18250 62980
rect 18310 62980 18320 63020
rect 18428 62982 18628 62988
rect 18428 62980 18440 62982
rect 18310 62960 18440 62980
rect 18118 62950 18440 62960
rect 18118 62948 18130 62950
rect 17930 62942 18130 62948
rect 18428 62948 18440 62950
rect 18616 62948 18628 62982
rect 18428 62942 18628 62948
rect 18660 62950 18740 62970
rect 17892 62904 17900 62938
rect 17890 62890 17900 62904
rect 17820 62870 17900 62890
rect 17930 62894 18130 62900
rect 17930 62860 17942 62894
rect 18118 62890 18130 62894
rect 18428 62894 18628 62900
rect 18428 62890 18440 62894
rect 18118 62860 18440 62890
rect 18616 62860 18628 62894
rect 18660 62890 18670 62950
rect 18730 62890 18740 62950
rect 18660 62870 18740 62890
rect 17930 62854 18130 62860
rect 17710 62730 17780 62790
rect 17710 62490 17730 62730
rect 17770 62490 17780 62730
rect 18240 62850 18320 62860
rect 18428 62854 18628 62860
rect 18240 62790 18250 62850
rect 18310 62790 18320 62850
rect 18240 62740 18320 62790
rect 18240 62680 18250 62740
rect 18310 62680 18320 62740
rect 17930 62672 18130 62678
rect 17820 62640 17900 62660
rect 17820 62580 17830 62640
rect 17890 62628 17900 62640
rect 17930 62638 17942 62672
rect 18118 62670 18130 62672
rect 18240 62670 18320 62680
rect 18790 62810 18800 63050
rect 18840 62810 18860 63050
rect 18790 62730 18860 62810
rect 18428 62672 18628 62678
rect 18428 62670 18440 62672
rect 18118 62640 18440 62670
rect 18118 62638 18130 62640
rect 17930 62632 18130 62638
rect 18428 62638 18440 62640
rect 18616 62638 18628 62672
rect 18428 62632 18628 62638
rect 18660 62640 18740 62660
rect 17892 62594 17900 62628
rect 17890 62580 17900 62594
rect 17820 62560 17900 62580
rect 17930 62584 18130 62590
rect 17930 62550 17942 62584
rect 18118 62580 18130 62584
rect 18428 62584 18628 62590
rect 18428 62580 18440 62584
rect 18118 62570 18440 62580
rect 18118 62550 18250 62570
rect 17930 62544 18130 62550
rect 18240 62510 18250 62550
rect 18310 62550 18440 62570
rect 18616 62550 18628 62584
rect 18660 62580 18670 62640
rect 18730 62580 18740 62640
rect 18660 62560 18740 62580
rect 18310 62510 18320 62550
rect 18428 62544 18628 62550
rect 18240 62500 18320 62510
rect 17710 61340 17780 62490
rect 17710 61080 17730 61340
rect 17770 61080 17780 61340
rect 18790 62490 18800 62730
rect 18840 62490 18860 62730
rect 18790 61340 18860 62490
rect 18240 61310 18320 61320
rect 17930 61272 18130 61278
rect 17820 61240 17900 61260
rect 17820 61180 17830 61240
rect 17890 61228 17900 61240
rect 17930 61238 17942 61272
rect 18118 61270 18130 61272
rect 18240 61270 18250 61310
rect 18118 61250 18250 61270
rect 18310 61270 18320 61310
rect 18428 61272 18628 61278
rect 18428 61270 18440 61272
rect 18310 61250 18440 61270
rect 18118 61240 18440 61250
rect 18118 61238 18130 61240
rect 17930 61232 18130 61238
rect 18428 61238 18440 61240
rect 18616 61238 18628 61272
rect 18428 61232 18628 61238
rect 18660 61240 18740 61260
rect 17892 61194 17900 61228
rect 17890 61180 17900 61194
rect 17820 61160 17900 61180
rect 17930 61184 18130 61190
rect 17930 61150 17942 61184
rect 18118 61180 18130 61184
rect 18428 61184 18628 61190
rect 18428 61180 18440 61184
rect 18118 61150 18440 61180
rect 18616 61150 18628 61184
rect 18660 61180 18670 61240
rect 18730 61180 18740 61240
rect 18660 61160 18740 61180
rect 17930 61144 18130 61150
rect 17710 61020 17780 61080
rect 17710 60780 17730 61020
rect 17770 60780 17780 61020
rect 18240 61140 18320 61150
rect 18428 61144 18628 61150
rect 18240 61080 18250 61140
rect 18310 61080 18320 61140
rect 18240 61030 18320 61080
rect 18240 60970 18250 61030
rect 18310 60970 18320 61030
rect 17930 60962 18130 60968
rect 17820 60930 17900 60950
rect 17820 60870 17830 60930
rect 17890 60918 17900 60930
rect 17930 60928 17942 60962
rect 18118 60960 18130 60962
rect 18240 60960 18320 60970
rect 18790 61100 18800 61340
rect 18840 61100 18860 61340
rect 18790 61020 18860 61100
rect 18428 60962 18628 60968
rect 18428 60960 18440 60962
rect 18118 60930 18440 60960
rect 18118 60928 18130 60930
rect 17930 60922 18130 60928
rect 18428 60928 18440 60930
rect 18616 60928 18628 60962
rect 18428 60922 18628 60928
rect 18660 60930 18740 60950
rect 17892 60884 17900 60918
rect 17890 60870 17900 60884
rect 17820 60850 17900 60870
rect 17930 60874 18130 60880
rect 17930 60840 17942 60874
rect 18118 60870 18130 60874
rect 18428 60874 18628 60880
rect 18428 60870 18440 60874
rect 18118 60860 18440 60870
rect 18118 60840 18250 60860
rect 17930 60834 18130 60840
rect 18240 60800 18250 60840
rect 18310 60840 18440 60860
rect 18616 60840 18628 60874
rect 18660 60870 18670 60930
rect 18730 60870 18740 60930
rect 18660 60850 18740 60870
rect 18310 60800 18320 60840
rect 18428 60834 18628 60840
rect 18240 60790 18320 60800
rect 17710 59630 17780 60780
rect 17710 59370 17730 59630
rect 17770 59370 17780 59630
rect 18790 60780 18800 61020
rect 18840 60780 18860 61020
rect 18790 59630 18860 60780
rect 18240 59600 18320 59610
rect 17930 59562 18130 59568
rect 17820 59530 17900 59550
rect 17820 59470 17830 59530
rect 17890 59518 17900 59530
rect 17930 59528 17942 59562
rect 18118 59560 18130 59562
rect 18240 59560 18250 59600
rect 18118 59540 18250 59560
rect 18310 59560 18320 59600
rect 18428 59562 18628 59568
rect 18428 59560 18440 59562
rect 18310 59540 18440 59560
rect 18118 59530 18440 59540
rect 18118 59528 18130 59530
rect 17930 59522 18130 59528
rect 18428 59528 18440 59530
rect 18616 59528 18628 59562
rect 18428 59522 18628 59528
rect 18660 59530 18740 59550
rect 17892 59484 17900 59518
rect 17890 59470 17900 59484
rect 17820 59450 17900 59470
rect 17930 59474 18130 59480
rect 17930 59440 17942 59474
rect 18118 59470 18130 59474
rect 18428 59474 18628 59480
rect 18428 59470 18440 59474
rect 18118 59440 18440 59470
rect 18616 59440 18628 59474
rect 18660 59470 18670 59530
rect 18730 59470 18740 59530
rect 18660 59450 18740 59470
rect 17930 59434 18130 59440
rect 17710 59310 17780 59370
rect 17710 59070 17730 59310
rect 17770 59070 17780 59310
rect 18240 59430 18320 59440
rect 18428 59434 18628 59440
rect 18240 59370 18250 59430
rect 18310 59370 18320 59430
rect 18240 59320 18320 59370
rect 18240 59260 18250 59320
rect 18310 59260 18320 59320
rect 17930 59252 18130 59258
rect 17820 59220 17900 59240
rect 17820 59160 17830 59220
rect 17890 59208 17900 59220
rect 17930 59218 17942 59252
rect 18118 59250 18130 59252
rect 18240 59250 18320 59260
rect 18790 59390 18800 59630
rect 18840 59390 18860 59630
rect 18790 59310 18860 59390
rect 18428 59252 18628 59258
rect 18428 59250 18440 59252
rect 18118 59220 18440 59250
rect 18118 59218 18130 59220
rect 17930 59212 18130 59218
rect 18428 59218 18440 59220
rect 18616 59218 18628 59252
rect 18428 59212 18628 59218
rect 18660 59220 18740 59240
rect 17892 59174 17900 59208
rect 17890 59160 17900 59174
rect 17820 59140 17900 59160
rect 17930 59164 18130 59170
rect 17930 59130 17942 59164
rect 18118 59160 18130 59164
rect 18428 59164 18628 59170
rect 18428 59160 18440 59164
rect 18118 59150 18440 59160
rect 18118 59130 18250 59150
rect 17930 59124 18130 59130
rect 18240 59090 18250 59130
rect 18310 59130 18440 59150
rect 18616 59130 18628 59164
rect 18660 59160 18670 59220
rect 18730 59160 18740 59220
rect 18660 59140 18740 59160
rect 18310 59090 18320 59130
rect 18428 59124 18628 59130
rect 18240 59080 18320 59090
rect 17710 57920 17780 59070
rect 17710 57660 17730 57920
rect 17770 57660 17780 57920
rect 18790 59070 18800 59310
rect 18840 59070 18860 59310
rect 18790 57920 18860 59070
rect 18240 57890 18320 57900
rect 17930 57852 18130 57858
rect 17820 57820 17900 57840
rect 17820 57760 17830 57820
rect 17890 57808 17900 57820
rect 17930 57818 17942 57852
rect 18118 57850 18130 57852
rect 18240 57850 18250 57890
rect 18118 57830 18250 57850
rect 18310 57850 18320 57890
rect 18428 57852 18628 57858
rect 18428 57850 18440 57852
rect 18310 57830 18440 57850
rect 18118 57820 18440 57830
rect 18118 57818 18130 57820
rect 17930 57812 18130 57818
rect 18428 57818 18440 57820
rect 18616 57818 18628 57852
rect 18428 57812 18628 57818
rect 18660 57820 18740 57840
rect 17892 57774 17900 57808
rect 17890 57760 17900 57774
rect 17820 57740 17900 57760
rect 17930 57764 18130 57770
rect 17930 57730 17942 57764
rect 18118 57760 18130 57764
rect 18428 57764 18628 57770
rect 18428 57760 18440 57764
rect 18118 57730 18440 57760
rect 18616 57730 18628 57764
rect 18660 57760 18670 57820
rect 18730 57760 18740 57820
rect 18660 57740 18740 57760
rect 17930 57724 18130 57730
rect 17710 57600 17780 57660
rect 17710 57360 17730 57600
rect 17770 57360 17780 57600
rect 18240 57720 18320 57730
rect 18428 57724 18628 57730
rect 18240 57660 18250 57720
rect 18310 57660 18320 57720
rect 18240 57610 18320 57660
rect 18240 57550 18250 57610
rect 18310 57550 18320 57610
rect 17930 57542 18130 57548
rect 17820 57510 17900 57530
rect 17820 57450 17830 57510
rect 17890 57498 17900 57510
rect 17930 57508 17942 57542
rect 18118 57540 18130 57542
rect 18240 57540 18320 57550
rect 18790 57680 18800 57920
rect 18840 57680 18860 57920
rect 18790 57600 18860 57680
rect 18428 57542 18628 57548
rect 18428 57540 18440 57542
rect 18118 57510 18440 57540
rect 18118 57508 18130 57510
rect 17930 57502 18130 57508
rect 18428 57508 18440 57510
rect 18616 57508 18628 57542
rect 18428 57502 18628 57508
rect 18660 57510 18740 57530
rect 17892 57464 17900 57498
rect 17890 57450 17900 57464
rect 17820 57430 17900 57450
rect 17930 57454 18130 57460
rect 17930 57420 17942 57454
rect 18118 57450 18130 57454
rect 18428 57454 18628 57460
rect 18428 57450 18440 57454
rect 18118 57440 18440 57450
rect 18118 57420 18250 57440
rect 17930 57414 18130 57420
rect 18240 57380 18250 57420
rect 18310 57420 18440 57440
rect 18616 57420 18628 57454
rect 18660 57450 18670 57510
rect 18730 57450 18740 57510
rect 18660 57430 18740 57450
rect 18310 57380 18320 57420
rect 18428 57414 18628 57420
rect 18240 57370 18320 57380
rect 17710 56210 17780 57360
rect 17710 55950 17730 56210
rect 17770 55950 17780 56210
rect 18790 57360 18800 57600
rect 18840 57360 18860 57600
rect 18790 56210 18860 57360
rect 18240 56180 18320 56190
rect 17930 56142 18130 56148
rect 17820 56110 17900 56130
rect 17820 56050 17830 56110
rect 17890 56098 17900 56110
rect 17930 56108 17942 56142
rect 18118 56140 18130 56142
rect 18240 56140 18250 56180
rect 18118 56120 18250 56140
rect 18310 56140 18320 56180
rect 18428 56142 18628 56148
rect 18428 56140 18440 56142
rect 18310 56120 18440 56140
rect 18118 56110 18440 56120
rect 18118 56108 18130 56110
rect 17930 56102 18130 56108
rect 18428 56108 18440 56110
rect 18616 56108 18628 56142
rect 18428 56102 18628 56108
rect 18660 56110 18740 56130
rect 17892 56064 17900 56098
rect 17890 56050 17900 56064
rect 17820 56030 17900 56050
rect 17930 56054 18130 56060
rect 17930 56020 17942 56054
rect 18118 56050 18130 56054
rect 18428 56054 18628 56060
rect 18428 56050 18440 56054
rect 18118 56020 18440 56050
rect 18616 56020 18628 56054
rect 18660 56050 18670 56110
rect 18730 56050 18740 56110
rect 18660 56030 18740 56050
rect 17930 56014 18130 56020
rect 17710 55890 17780 55950
rect 17710 55650 17730 55890
rect 17770 55650 17780 55890
rect 18240 56010 18320 56020
rect 18428 56014 18628 56020
rect 18240 55950 18250 56010
rect 18310 55950 18320 56010
rect 18240 55900 18320 55950
rect 18240 55840 18250 55900
rect 18310 55840 18320 55900
rect 17930 55832 18130 55838
rect 17820 55800 17900 55820
rect 17820 55740 17830 55800
rect 17890 55788 17900 55800
rect 17930 55798 17942 55832
rect 18118 55830 18130 55832
rect 18240 55830 18320 55840
rect 18790 55970 18800 56210
rect 18840 55970 18860 56210
rect 18790 55890 18860 55970
rect 18428 55832 18628 55838
rect 18428 55830 18440 55832
rect 18118 55800 18440 55830
rect 18118 55798 18130 55800
rect 17930 55792 18130 55798
rect 18428 55798 18440 55800
rect 18616 55798 18628 55832
rect 18428 55792 18628 55798
rect 18660 55800 18740 55820
rect 17892 55754 17900 55788
rect 17890 55740 17900 55754
rect 17820 55720 17900 55740
rect 17930 55744 18130 55750
rect 17930 55710 17942 55744
rect 18118 55740 18130 55744
rect 18428 55744 18628 55750
rect 18428 55740 18440 55744
rect 18118 55730 18440 55740
rect 18118 55710 18250 55730
rect 17930 55704 18130 55710
rect 18240 55670 18250 55710
rect 18310 55710 18440 55730
rect 18616 55710 18628 55744
rect 18660 55740 18670 55800
rect 18730 55740 18740 55800
rect 18660 55720 18740 55740
rect 18310 55670 18320 55710
rect 18428 55704 18628 55710
rect 18240 55660 18320 55670
rect 17710 54500 17780 55650
rect 17710 54240 17730 54500
rect 17770 54240 17780 54500
rect 18790 55650 18800 55890
rect 18840 55650 18860 55890
rect 18790 54500 18860 55650
rect 18240 54470 18320 54480
rect 17930 54432 18130 54438
rect 17820 54400 17900 54420
rect 17820 54340 17830 54400
rect 17890 54388 17900 54400
rect 17930 54398 17942 54432
rect 18118 54430 18130 54432
rect 18240 54430 18250 54470
rect 18118 54410 18250 54430
rect 18310 54430 18320 54470
rect 18428 54432 18628 54438
rect 18428 54430 18440 54432
rect 18310 54410 18440 54430
rect 18118 54400 18440 54410
rect 18118 54398 18130 54400
rect 17930 54392 18130 54398
rect 18428 54398 18440 54400
rect 18616 54398 18628 54432
rect 18428 54392 18628 54398
rect 18660 54400 18740 54420
rect 17892 54354 17900 54388
rect 17890 54340 17900 54354
rect 17820 54320 17900 54340
rect 17930 54344 18130 54350
rect 17930 54310 17942 54344
rect 18118 54340 18130 54344
rect 18428 54344 18628 54350
rect 18428 54340 18440 54344
rect 18118 54310 18440 54340
rect 18616 54310 18628 54344
rect 18660 54340 18670 54400
rect 18730 54340 18740 54400
rect 18660 54320 18740 54340
rect 17930 54304 18130 54310
rect 17710 54180 17780 54240
rect 17710 53940 17730 54180
rect 17770 53940 17780 54180
rect 18240 54300 18320 54310
rect 18428 54304 18628 54310
rect 18240 54240 18250 54300
rect 18310 54240 18320 54300
rect 18240 54190 18320 54240
rect 18240 54130 18250 54190
rect 18310 54130 18320 54190
rect 17930 54122 18130 54128
rect 17820 54090 17900 54110
rect 17820 54030 17830 54090
rect 17890 54078 17900 54090
rect 17930 54088 17942 54122
rect 18118 54120 18130 54122
rect 18240 54120 18320 54130
rect 18790 54260 18800 54500
rect 18840 54260 18860 54500
rect 18790 54180 18860 54260
rect 18428 54122 18628 54128
rect 18428 54120 18440 54122
rect 18118 54090 18440 54120
rect 18118 54088 18130 54090
rect 17930 54082 18130 54088
rect 18428 54088 18440 54090
rect 18616 54088 18628 54122
rect 18428 54082 18628 54088
rect 18660 54090 18740 54110
rect 17892 54044 17900 54078
rect 17890 54030 17900 54044
rect 17820 54010 17900 54030
rect 17930 54034 18130 54040
rect 17930 54000 17942 54034
rect 18118 54030 18130 54034
rect 18428 54034 18628 54040
rect 18428 54030 18440 54034
rect 18118 54020 18440 54030
rect 18118 54000 18250 54020
rect 17930 53994 18130 54000
rect 18240 53960 18250 54000
rect 18310 54000 18440 54020
rect 18616 54000 18628 54034
rect 18660 54030 18670 54090
rect 18730 54030 18740 54090
rect 18660 54010 18740 54030
rect 18310 53960 18320 54000
rect 18428 53994 18628 54000
rect 18240 53950 18320 53960
rect 17710 52790 17780 53940
rect 17710 52530 17730 52790
rect 17770 52530 17780 52790
rect 18790 53940 18800 54180
rect 18840 53940 18860 54180
rect 18790 52790 18860 53940
rect 18240 52760 18320 52770
rect 17930 52722 18130 52728
rect 17820 52690 17900 52710
rect 17820 52630 17830 52690
rect 17890 52678 17900 52690
rect 17930 52688 17942 52722
rect 18118 52720 18130 52722
rect 18240 52720 18250 52760
rect 18118 52700 18250 52720
rect 18310 52720 18320 52760
rect 18428 52722 18628 52728
rect 18428 52720 18440 52722
rect 18310 52700 18440 52720
rect 18118 52690 18440 52700
rect 18118 52688 18130 52690
rect 17930 52682 18130 52688
rect 18428 52688 18440 52690
rect 18616 52688 18628 52722
rect 18428 52682 18628 52688
rect 18660 52690 18740 52710
rect 17892 52644 17900 52678
rect 17890 52630 17900 52644
rect 17820 52610 17900 52630
rect 17930 52634 18130 52640
rect 17930 52600 17942 52634
rect 18118 52630 18130 52634
rect 18428 52634 18628 52640
rect 18428 52630 18440 52634
rect 18118 52600 18440 52630
rect 18616 52600 18628 52634
rect 18660 52630 18670 52690
rect 18730 52630 18740 52690
rect 18660 52610 18740 52630
rect 17930 52594 18130 52600
rect 17710 52470 17780 52530
rect 17710 52230 17730 52470
rect 17770 52230 17780 52470
rect 18240 52590 18320 52600
rect 18428 52594 18628 52600
rect 18240 52530 18250 52590
rect 18310 52530 18320 52590
rect 18240 52480 18320 52530
rect 18240 52420 18250 52480
rect 18310 52420 18320 52480
rect 17930 52412 18130 52418
rect 17820 52380 17900 52400
rect 17820 52320 17830 52380
rect 17890 52368 17900 52380
rect 17930 52378 17942 52412
rect 18118 52410 18130 52412
rect 18240 52410 18320 52420
rect 18790 52550 18800 52790
rect 18840 52550 18860 52790
rect 18790 52470 18860 52550
rect 18428 52412 18628 52418
rect 18428 52410 18440 52412
rect 18118 52380 18440 52410
rect 18118 52378 18130 52380
rect 17930 52372 18130 52378
rect 18428 52378 18440 52380
rect 18616 52378 18628 52412
rect 18428 52372 18628 52378
rect 18660 52380 18740 52400
rect 17892 52334 17900 52368
rect 17890 52320 17900 52334
rect 17820 52300 17900 52320
rect 17930 52324 18130 52330
rect 17930 52290 17942 52324
rect 18118 52320 18130 52324
rect 18428 52324 18628 52330
rect 18428 52320 18440 52324
rect 18118 52310 18440 52320
rect 18118 52290 18250 52310
rect 17930 52284 18130 52290
rect 18240 52250 18250 52290
rect 18310 52290 18440 52310
rect 18616 52290 18628 52324
rect 18660 52320 18670 52380
rect 18730 52320 18740 52380
rect 18660 52300 18740 52320
rect 18310 52250 18320 52290
rect 18428 52284 18628 52290
rect 18240 52240 18320 52250
rect 17710 51080 17780 52230
rect 17710 50820 17730 51080
rect 17770 50820 17780 51080
rect 18790 52230 18800 52470
rect 18840 52230 18860 52470
rect 18790 51080 18860 52230
rect 18240 51050 18320 51060
rect 17930 51012 18130 51018
rect 17820 50980 17900 51000
rect 17820 50920 17830 50980
rect 17890 50968 17900 50980
rect 17930 50978 17942 51012
rect 18118 51010 18130 51012
rect 18240 51010 18250 51050
rect 18118 50990 18250 51010
rect 18310 51010 18320 51050
rect 18428 51012 18628 51018
rect 18428 51010 18440 51012
rect 18310 50990 18440 51010
rect 18118 50980 18440 50990
rect 18118 50978 18130 50980
rect 17930 50972 18130 50978
rect 18428 50978 18440 50980
rect 18616 50978 18628 51012
rect 18428 50972 18628 50978
rect 18660 50980 18740 51000
rect 17892 50934 17900 50968
rect 17890 50920 17900 50934
rect 17820 50900 17900 50920
rect 17930 50924 18130 50930
rect 17930 50890 17942 50924
rect 18118 50920 18130 50924
rect 18428 50924 18628 50930
rect 18428 50920 18440 50924
rect 18118 50890 18440 50920
rect 18616 50890 18628 50924
rect 18660 50920 18670 50980
rect 18730 50920 18740 50980
rect 18660 50900 18740 50920
rect 17930 50884 18130 50890
rect 17710 50760 17780 50820
rect 17710 50520 17730 50760
rect 17770 50520 17780 50760
rect 18240 50880 18320 50890
rect 18428 50884 18628 50890
rect 18240 50820 18250 50880
rect 18310 50820 18320 50880
rect 18240 50770 18320 50820
rect 18240 50710 18250 50770
rect 18310 50710 18320 50770
rect 17930 50702 18130 50708
rect 17820 50670 17900 50690
rect 17820 50610 17830 50670
rect 17890 50658 17900 50670
rect 17930 50668 17942 50702
rect 18118 50700 18130 50702
rect 18240 50700 18320 50710
rect 18790 50840 18800 51080
rect 18840 50840 18860 51080
rect 18790 50760 18860 50840
rect 18428 50702 18628 50708
rect 18428 50700 18440 50702
rect 18118 50670 18440 50700
rect 18118 50668 18130 50670
rect 17930 50662 18130 50668
rect 18428 50668 18440 50670
rect 18616 50668 18628 50702
rect 18428 50662 18628 50668
rect 18660 50670 18740 50690
rect 17892 50624 17900 50658
rect 17890 50610 17900 50624
rect 17820 50590 17900 50610
rect 17930 50614 18130 50620
rect 17930 50580 17942 50614
rect 18118 50610 18130 50614
rect 18428 50614 18628 50620
rect 18428 50610 18440 50614
rect 18118 50600 18440 50610
rect 18118 50580 18250 50600
rect 17930 50574 18130 50580
rect 18240 50540 18250 50580
rect 18310 50580 18440 50600
rect 18616 50580 18628 50614
rect 18660 50610 18670 50670
rect 18730 50610 18740 50670
rect 18660 50590 18740 50610
rect 18310 50540 18320 50580
rect 18428 50574 18628 50580
rect 18240 50530 18320 50540
rect 17710 49370 17780 50520
rect 17710 49110 17730 49370
rect 17770 49110 17780 49370
rect 18790 50520 18800 50760
rect 18840 50520 18860 50760
rect 18790 49370 18860 50520
rect 18240 49340 18320 49350
rect 17930 49302 18130 49308
rect 17820 49270 17900 49290
rect 17820 49210 17830 49270
rect 17890 49258 17900 49270
rect 17930 49268 17942 49302
rect 18118 49300 18130 49302
rect 18240 49300 18250 49340
rect 18118 49280 18250 49300
rect 18310 49300 18320 49340
rect 18428 49302 18628 49308
rect 18428 49300 18440 49302
rect 18310 49280 18440 49300
rect 18118 49270 18440 49280
rect 18118 49268 18130 49270
rect 17930 49262 18130 49268
rect 18428 49268 18440 49270
rect 18616 49268 18628 49302
rect 18428 49262 18628 49268
rect 18660 49270 18740 49290
rect 17892 49224 17900 49258
rect 17890 49210 17900 49224
rect 17820 49190 17900 49210
rect 17930 49214 18130 49220
rect 17930 49180 17942 49214
rect 18118 49210 18130 49214
rect 18428 49214 18628 49220
rect 18428 49210 18440 49214
rect 18118 49180 18440 49210
rect 18616 49180 18628 49214
rect 18660 49210 18670 49270
rect 18730 49210 18740 49270
rect 18660 49190 18740 49210
rect 17930 49174 18130 49180
rect 17710 49050 17780 49110
rect 17710 48810 17730 49050
rect 17770 48810 17780 49050
rect 18240 49170 18320 49180
rect 18428 49174 18628 49180
rect 18240 49110 18250 49170
rect 18310 49110 18320 49170
rect 18240 49060 18320 49110
rect 18240 49000 18250 49060
rect 18310 49000 18320 49060
rect 17930 48992 18130 48998
rect 17820 48960 17900 48980
rect 17820 48900 17830 48960
rect 17890 48948 17900 48960
rect 17930 48958 17942 48992
rect 18118 48990 18130 48992
rect 18240 48990 18320 49000
rect 18790 49130 18800 49370
rect 18840 49130 18860 49370
rect 18790 49050 18860 49130
rect 18428 48992 18628 48998
rect 18428 48990 18440 48992
rect 18118 48960 18440 48990
rect 18118 48958 18130 48960
rect 17930 48952 18130 48958
rect 18428 48958 18440 48960
rect 18616 48958 18628 48992
rect 18428 48952 18628 48958
rect 18660 48960 18740 48980
rect 17892 48914 17900 48948
rect 17890 48900 17900 48914
rect 17820 48880 17900 48900
rect 17930 48904 18130 48910
rect 17930 48870 17942 48904
rect 18118 48900 18130 48904
rect 18428 48904 18628 48910
rect 18428 48900 18440 48904
rect 18118 48890 18440 48900
rect 18118 48870 18250 48890
rect 17930 48864 18130 48870
rect 18240 48830 18250 48870
rect 18310 48870 18440 48890
rect 18616 48870 18628 48904
rect 18660 48900 18670 48960
rect 18730 48900 18740 48960
rect 18660 48880 18740 48900
rect 18310 48830 18320 48870
rect 18428 48864 18628 48870
rect 18240 48820 18320 48830
rect 17710 47660 17780 48810
rect 17710 47400 17730 47660
rect 17770 47400 17780 47660
rect 18790 48810 18800 49050
rect 18840 48810 18860 49050
rect 18790 47660 18860 48810
rect 18240 47630 18320 47640
rect 17930 47592 18130 47598
rect 17820 47560 17900 47580
rect 17820 47500 17830 47560
rect 17890 47548 17900 47560
rect 17930 47558 17942 47592
rect 18118 47590 18130 47592
rect 18240 47590 18250 47630
rect 18118 47570 18250 47590
rect 18310 47590 18320 47630
rect 18428 47592 18628 47598
rect 18428 47590 18440 47592
rect 18310 47570 18440 47590
rect 18118 47560 18440 47570
rect 18118 47558 18130 47560
rect 17930 47552 18130 47558
rect 18428 47558 18440 47560
rect 18616 47558 18628 47592
rect 18428 47552 18628 47558
rect 18660 47560 18740 47580
rect 17892 47514 17900 47548
rect 17890 47500 17900 47514
rect 17820 47480 17900 47500
rect 17930 47504 18130 47510
rect 17930 47470 17942 47504
rect 18118 47500 18130 47504
rect 18428 47504 18628 47510
rect 18428 47500 18440 47504
rect 18118 47470 18440 47500
rect 18616 47470 18628 47504
rect 18660 47500 18670 47560
rect 18730 47500 18740 47560
rect 18660 47480 18740 47500
rect 17930 47464 18130 47470
rect 17710 47340 17780 47400
rect 17710 47100 17730 47340
rect 17770 47100 17780 47340
rect 18240 47460 18320 47470
rect 18428 47464 18628 47470
rect 18240 47400 18250 47460
rect 18310 47400 18320 47460
rect 18240 47350 18320 47400
rect 18240 47290 18250 47350
rect 18310 47290 18320 47350
rect 17930 47282 18130 47288
rect 17820 47250 17900 47270
rect 17820 47190 17830 47250
rect 17890 47238 17900 47250
rect 17930 47248 17942 47282
rect 18118 47280 18130 47282
rect 18240 47280 18320 47290
rect 18790 47420 18800 47660
rect 18840 47420 18860 47660
rect 18790 47340 18860 47420
rect 18428 47282 18628 47288
rect 18428 47280 18440 47282
rect 18118 47250 18440 47280
rect 18118 47248 18130 47250
rect 17930 47242 18130 47248
rect 18428 47248 18440 47250
rect 18616 47248 18628 47282
rect 18428 47242 18628 47248
rect 18660 47250 18740 47270
rect 17892 47204 17900 47238
rect 17890 47190 17900 47204
rect 17820 47170 17900 47190
rect 17930 47194 18130 47200
rect 17930 47160 17942 47194
rect 18118 47190 18130 47194
rect 18428 47194 18628 47200
rect 18428 47190 18440 47194
rect 18118 47180 18440 47190
rect 18118 47160 18250 47180
rect 17930 47154 18130 47160
rect 18240 47120 18250 47160
rect 18310 47160 18440 47180
rect 18616 47160 18628 47194
rect 18660 47190 18670 47250
rect 18730 47190 18740 47250
rect 18660 47170 18740 47190
rect 18310 47120 18320 47160
rect 18428 47154 18628 47160
rect 18240 47110 18320 47120
rect 17710 45950 17780 47100
rect 17710 45690 17730 45950
rect 17770 45690 17780 45950
rect 18790 47100 18800 47340
rect 18840 47100 18860 47340
rect 18790 45950 18860 47100
rect 18240 45920 18320 45930
rect 17930 45882 18130 45888
rect 17820 45850 17900 45870
rect 17820 45790 17830 45850
rect 17890 45838 17900 45850
rect 17930 45848 17942 45882
rect 18118 45880 18130 45882
rect 18240 45880 18250 45920
rect 18118 45860 18250 45880
rect 18310 45880 18320 45920
rect 18428 45882 18628 45888
rect 18428 45880 18440 45882
rect 18310 45860 18440 45880
rect 18118 45850 18440 45860
rect 18118 45848 18130 45850
rect 17930 45842 18130 45848
rect 18428 45848 18440 45850
rect 18616 45848 18628 45882
rect 18428 45842 18628 45848
rect 18660 45850 18740 45870
rect 17892 45804 17900 45838
rect 17890 45790 17900 45804
rect 17820 45770 17900 45790
rect 17930 45794 18130 45800
rect 17930 45760 17942 45794
rect 18118 45790 18130 45794
rect 18428 45794 18628 45800
rect 18428 45790 18440 45794
rect 18118 45760 18440 45790
rect 18616 45760 18628 45794
rect 18660 45790 18670 45850
rect 18730 45790 18740 45850
rect 18660 45770 18740 45790
rect 17930 45754 18130 45760
rect 17710 45630 17780 45690
rect 17710 45390 17730 45630
rect 17770 45390 17780 45630
rect 18240 45750 18320 45760
rect 18428 45754 18628 45760
rect 18240 45690 18250 45750
rect 18310 45690 18320 45750
rect 18240 45640 18320 45690
rect 18240 45580 18250 45640
rect 18310 45580 18320 45640
rect 17930 45572 18130 45578
rect 17820 45540 17900 45560
rect 17820 45480 17830 45540
rect 17890 45528 17900 45540
rect 17930 45538 17942 45572
rect 18118 45570 18130 45572
rect 18240 45570 18320 45580
rect 18790 45710 18800 45950
rect 18840 45710 18860 45950
rect 18790 45630 18860 45710
rect 18428 45572 18628 45578
rect 18428 45570 18440 45572
rect 18118 45540 18440 45570
rect 18118 45538 18130 45540
rect 17930 45532 18130 45538
rect 18428 45538 18440 45540
rect 18616 45538 18628 45572
rect 18428 45532 18628 45538
rect 18660 45540 18740 45560
rect 17892 45494 17900 45528
rect 17890 45480 17900 45494
rect 17820 45460 17900 45480
rect 17930 45484 18130 45490
rect 17930 45450 17942 45484
rect 18118 45480 18130 45484
rect 18428 45484 18628 45490
rect 18428 45480 18440 45484
rect 18118 45470 18440 45480
rect 18118 45450 18250 45470
rect 17930 45444 18130 45450
rect 18240 45410 18250 45450
rect 18310 45450 18440 45470
rect 18616 45450 18628 45484
rect 18660 45480 18670 45540
rect 18730 45480 18740 45540
rect 18660 45460 18740 45480
rect 18310 45410 18320 45450
rect 18428 45444 18628 45450
rect 18240 45400 18320 45410
rect 17710 44240 17780 45390
rect 17710 43980 17730 44240
rect 17770 43980 17780 44240
rect 18790 45390 18800 45630
rect 18840 45390 18860 45630
rect 18790 44240 18860 45390
rect 18240 44210 18320 44220
rect 17930 44172 18130 44178
rect 17820 44140 17900 44160
rect 17820 44080 17830 44140
rect 17890 44128 17900 44140
rect 17930 44138 17942 44172
rect 18118 44170 18130 44172
rect 18240 44170 18250 44210
rect 18118 44150 18250 44170
rect 18310 44170 18320 44210
rect 18428 44172 18628 44178
rect 18428 44170 18440 44172
rect 18310 44150 18440 44170
rect 18118 44140 18440 44150
rect 18118 44138 18130 44140
rect 17930 44132 18130 44138
rect 18428 44138 18440 44140
rect 18616 44138 18628 44172
rect 18428 44132 18628 44138
rect 18660 44140 18740 44160
rect 17892 44094 17900 44128
rect 17890 44080 17900 44094
rect 17820 44060 17900 44080
rect 17930 44084 18130 44090
rect 17930 44050 17942 44084
rect 18118 44080 18130 44084
rect 18428 44084 18628 44090
rect 18428 44080 18440 44084
rect 18118 44050 18440 44080
rect 18616 44050 18628 44084
rect 18660 44080 18670 44140
rect 18730 44080 18740 44140
rect 18660 44060 18740 44080
rect 17930 44044 18130 44050
rect 17710 43920 17780 43980
rect 17710 43680 17730 43920
rect 17770 43680 17780 43920
rect 18240 44040 18320 44050
rect 18428 44044 18628 44050
rect 18240 43980 18250 44040
rect 18310 43980 18320 44040
rect 18240 43930 18320 43980
rect 18240 43870 18250 43930
rect 18310 43870 18320 43930
rect 17930 43862 18130 43868
rect 17820 43830 17900 43850
rect 17820 43770 17830 43830
rect 17890 43818 17900 43830
rect 17930 43828 17942 43862
rect 18118 43860 18130 43862
rect 18240 43860 18320 43870
rect 18790 44000 18800 44240
rect 18840 44000 18860 44240
rect 18790 43920 18860 44000
rect 18428 43862 18628 43868
rect 18428 43860 18440 43862
rect 18118 43830 18440 43860
rect 18118 43828 18130 43830
rect 17930 43822 18130 43828
rect 18428 43828 18440 43830
rect 18616 43828 18628 43862
rect 18428 43822 18628 43828
rect 18660 43830 18740 43850
rect 17892 43784 17900 43818
rect 17890 43770 17900 43784
rect 17820 43750 17900 43770
rect 17930 43774 18130 43780
rect 17930 43740 17942 43774
rect 18118 43770 18130 43774
rect 18428 43774 18628 43780
rect 18428 43770 18440 43774
rect 18118 43760 18440 43770
rect 18118 43740 18250 43760
rect 17930 43734 18130 43740
rect 18240 43700 18250 43740
rect 18310 43740 18440 43760
rect 18616 43740 18628 43774
rect 18660 43770 18670 43830
rect 18730 43770 18740 43830
rect 18660 43750 18740 43770
rect 18310 43700 18320 43740
rect 18428 43734 18628 43740
rect 18240 43690 18320 43700
rect 17710 42530 17780 43680
rect 17710 42270 17730 42530
rect 17770 42270 17780 42530
rect 18790 43680 18800 43920
rect 18840 43680 18860 43920
rect 18790 42530 18860 43680
rect 18240 42500 18320 42510
rect 17930 42462 18130 42468
rect 17820 42430 17900 42450
rect 17820 42370 17830 42430
rect 17890 42418 17900 42430
rect 17930 42428 17942 42462
rect 18118 42460 18130 42462
rect 18240 42460 18250 42500
rect 18118 42440 18250 42460
rect 18310 42460 18320 42500
rect 18428 42462 18628 42468
rect 18428 42460 18440 42462
rect 18310 42440 18440 42460
rect 18118 42430 18440 42440
rect 18118 42428 18130 42430
rect 17930 42422 18130 42428
rect 18428 42428 18440 42430
rect 18616 42428 18628 42462
rect 18428 42422 18628 42428
rect 18660 42430 18740 42450
rect 17892 42384 17900 42418
rect 17890 42370 17900 42384
rect 17820 42350 17900 42370
rect 17930 42374 18130 42380
rect 17930 42340 17942 42374
rect 18118 42370 18130 42374
rect 18428 42374 18628 42380
rect 18428 42370 18440 42374
rect 18118 42340 18440 42370
rect 18616 42340 18628 42374
rect 18660 42370 18670 42430
rect 18730 42370 18740 42430
rect 18660 42350 18740 42370
rect 17930 42334 18130 42340
rect 17710 42210 17780 42270
rect 17710 41970 17730 42210
rect 17770 41970 17780 42210
rect 18240 42330 18320 42340
rect 18428 42334 18628 42340
rect 18240 42270 18250 42330
rect 18310 42270 18320 42330
rect 18240 42220 18320 42270
rect 18240 42160 18250 42220
rect 18310 42160 18320 42220
rect 17930 42152 18130 42158
rect 17820 42120 17900 42140
rect 17820 42060 17830 42120
rect 17890 42108 17900 42120
rect 17930 42118 17942 42152
rect 18118 42150 18130 42152
rect 18240 42150 18320 42160
rect 18790 42290 18800 42530
rect 18840 42290 18860 42530
rect 18790 42210 18860 42290
rect 18428 42152 18628 42158
rect 18428 42150 18440 42152
rect 18118 42120 18440 42150
rect 18118 42118 18130 42120
rect 17930 42112 18130 42118
rect 18428 42118 18440 42120
rect 18616 42118 18628 42152
rect 18428 42112 18628 42118
rect 18660 42120 18740 42140
rect 17892 42074 17900 42108
rect 17890 42060 17900 42074
rect 17820 42040 17900 42060
rect 17930 42064 18130 42070
rect 17930 42030 17942 42064
rect 18118 42060 18130 42064
rect 18428 42064 18628 42070
rect 18428 42060 18440 42064
rect 18118 42050 18440 42060
rect 18118 42030 18250 42050
rect 17930 42024 18130 42030
rect 18240 41990 18250 42030
rect 18310 42030 18440 42050
rect 18616 42030 18628 42064
rect 18660 42060 18670 42120
rect 18730 42060 18740 42120
rect 18660 42040 18740 42060
rect 18310 41990 18320 42030
rect 18428 42024 18628 42030
rect 18240 41980 18320 41990
rect 17710 40820 17780 41970
rect 17710 40560 17730 40820
rect 17770 40560 17780 40820
rect 18790 41970 18800 42210
rect 18840 41970 18860 42210
rect 18790 40820 18860 41970
rect 18240 40790 18320 40800
rect 17930 40752 18130 40758
rect 17820 40720 17900 40740
rect 17820 40660 17830 40720
rect 17890 40708 17900 40720
rect 17930 40718 17942 40752
rect 18118 40750 18130 40752
rect 18240 40750 18250 40790
rect 18118 40730 18250 40750
rect 18310 40750 18320 40790
rect 18428 40752 18628 40758
rect 18428 40750 18440 40752
rect 18310 40730 18440 40750
rect 18118 40720 18440 40730
rect 18118 40718 18130 40720
rect 17930 40712 18130 40718
rect 18428 40718 18440 40720
rect 18616 40718 18628 40752
rect 18428 40712 18628 40718
rect 18660 40720 18740 40740
rect 17892 40674 17900 40708
rect 17890 40660 17900 40674
rect 17820 40640 17900 40660
rect 17930 40664 18130 40670
rect 17930 40630 17942 40664
rect 18118 40660 18130 40664
rect 18428 40664 18628 40670
rect 18428 40660 18440 40664
rect 18118 40630 18440 40660
rect 18616 40630 18628 40664
rect 18660 40660 18670 40720
rect 18730 40660 18740 40720
rect 18660 40640 18740 40660
rect 17930 40624 18130 40630
rect 17710 40500 17780 40560
rect 17710 40260 17730 40500
rect 17770 40260 17780 40500
rect 18240 40620 18320 40630
rect 18428 40624 18628 40630
rect 18240 40560 18250 40620
rect 18310 40560 18320 40620
rect 18240 40510 18320 40560
rect 18240 40450 18250 40510
rect 18310 40450 18320 40510
rect 17930 40442 18130 40448
rect 17820 40410 17900 40430
rect 17820 40350 17830 40410
rect 17890 40398 17900 40410
rect 17930 40408 17942 40442
rect 18118 40440 18130 40442
rect 18240 40440 18320 40450
rect 18790 40580 18800 40820
rect 18840 40580 18860 40820
rect 18790 40500 18860 40580
rect 18428 40442 18628 40448
rect 18428 40440 18440 40442
rect 18118 40410 18440 40440
rect 18118 40408 18130 40410
rect 17930 40402 18130 40408
rect 18428 40408 18440 40410
rect 18616 40408 18628 40442
rect 18428 40402 18628 40408
rect 18660 40410 18740 40430
rect 17892 40364 17900 40398
rect 17890 40350 17900 40364
rect 17820 40330 17900 40350
rect 17930 40354 18130 40360
rect 17930 40320 17942 40354
rect 18118 40350 18130 40354
rect 18428 40354 18628 40360
rect 18428 40350 18440 40354
rect 18118 40340 18440 40350
rect 18118 40320 18250 40340
rect 17930 40314 18130 40320
rect 18240 40280 18250 40320
rect 18310 40320 18440 40340
rect 18616 40320 18628 40354
rect 18660 40350 18670 40410
rect 18730 40350 18740 40410
rect 18660 40330 18740 40350
rect 18310 40280 18320 40320
rect 18428 40314 18628 40320
rect 18240 40270 18320 40280
rect 17710 39690 17780 40260
rect 18790 40260 18800 40500
rect 18840 40260 18860 40500
rect 18790 39690 18860 40260
rect 17710 39680 17790 39690
rect 17710 39620 17720 39680
rect 17780 39620 17790 39680
rect 18780 39680 18860 39690
rect 18780 39620 18790 39680
rect 18850 39620 18860 39680
rect 18780 39610 18860 39620
rect 18890 66480 18920 67050
rect 18890 66470 18950 66480
rect 18890 66400 18950 66410
rect 18890 64770 18920 66400
rect 18980 65950 19010 67050
rect 18950 65940 19010 65950
rect 18950 65870 19010 65880
rect 18890 64760 18950 64770
rect 18890 64690 18950 64700
rect 18890 63060 18920 64690
rect 18980 64240 19010 65870
rect 18950 64230 19010 64240
rect 18950 64160 19010 64170
rect 18890 63050 18950 63060
rect 18890 62980 18950 62990
rect 18890 61350 18920 62980
rect 18980 62530 19010 64160
rect 18950 62520 19010 62530
rect 18950 62450 19010 62460
rect 18890 61340 18950 61350
rect 18890 61270 18950 61280
rect 18890 59640 18920 61270
rect 18980 60820 19010 62450
rect 18950 60810 19010 60820
rect 18950 60740 19010 60750
rect 18890 59630 18950 59640
rect 18890 59560 18950 59570
rect 18890 57930 18920 59560
rect 18980 59110 19010 60740
rect 18950 59100 19010 59110
rect 18950 59030 19010 59040
rect 18890 57920 18950 57930
rect 18890 57850 18950 57860
rect 18890 56220 18920 57850
rect 18980 57400 19010 59030
rect 18950 57390 19010 57400
rect 18950 57320 19010 57330
rect 18890 56210 18950 56220
rect 18890 56140 18950 56150
rect 18890 54510 18920 56140
rect 18980 55690 19010 57320
rect 18950 55680 19010 55690
rect 18950 55610 19010 55620
rect 18890 54500 18950 54510
rect 18890 54430 18950 54440
rect 18890 52800 18920 54430
rect 18980 53980 19010 55610
rect 18950 53970 19010 53980
rect 18950 53900 19010 53910
rect 18890 52790 18950 52800
rect 18890 52720 18950 52730
rect 18890 51090 18920 52720
rect 18980 52270 19010 53900
rect 18950 52260 19010 52270
rect 18950 52190 19010 52200
rect 18890 51080 18950 51090
rect 18890 51010 18950 51020
rect 18890 49380 18920 51010
rect 18980 50560 19010 52190
rect 18950 50550 19010 50560
rect 18950 50480 19010 50490
rect 18890 49370 18950 49380
rect 18890 49300 18950 49310
rect 18890 47670 18920 49300
rect 18980 48850 19010 50480
rect 18950 48840 19010 48850
rect 18950 48770 19010 48780
rect 18890 47660 18950 47670
rect 18890 47590 18950 47600
rect 18890 45960 18920 47590
rect 18980 47140 19010 48770
rect 18950 47130 19010 47140
rect 18950 47060 19010 47070
rect 18890 45950 18950 45960
rect 18890 45880 18950 45890
rect 18890 44250 18920 45880
rect 18980 45430 19010 47060
rect 18950 45420 19010 45430
rect 18950 45350 19010 45360
rect 18890 44240 18950 44250
rect 18890 44170 18950 44180
rect 18890 42540 18920 44170
rect 18980 43720 19010 45350
rect 18950 43710 19010 43720
rect 18950 43640 19010 43650
rect 18890 42530 18950 42540
rect 18890 42460 18950 42470
rect 18890 40830 18920 42460
rect 18980 42010 19010 43640
rect 18950 42000 19010 42010
rect 18950 41930 19010 41940
rect 18890 40820 18950 40830
rect 18890 40750 18950 40760
rect 17240 39220 17300 39230
rect 17420 39230 17680 39240
rect 14250 39160 14310 39170
rect 17480 39210 17680 39230
rect 17420 39160 17480 39170
rect 18890 38840 18920 40750
rect 18980 40300 19010 41930
rect 18950 40290 19010 40300
rect 18950 40220 19010 40230
rect 18980 39690 19010 40220
rect 18950 39680 19010 39690
rect 18950 39610 19010 39620
rect 19040 66390 19070 67050
rect 19040 66380 19100 66390
rect 19040 66310 19100 66320
rect 19040 64680 19070 66310
rect 19040 64670 19100 64680
rect 19040 64600 19100 64610
rect 19040 62970 19070 64600
rect 19040 62960 19100 62970
rect 19040 62890 19100 62900
rect 19040 61260 19070 62890
rect 19040 61250 19100 61260
rect 19040 61180 19100 61190
rect 19040 45870 19070 61180
rect 19160 59550 19190 67050
rect 19160 59540 19220 59550
rect 19160 59470 19220 59480
rect 19160 57840 19190 59470
rect 19160 57830 19220 57840
rect 19160 57760 19220 57770
rect 19160 56130 19190 57760
rect 19160 56120 19220 56130
rect 19160 56050 19220 56060
rect 19160 54420 19190 56050
rect 19160 54410 19220 54420
rect 19160 54340 19220 54350
rect 19160 52710 19190 54340
rect 19160 52700 19220 52710
rect 19160 52630 19220 52640
rect 19160 51000 19190 52630
rect 19160 50990 19220 51000
rect 19160 50920 19220 50930
rect 19160 49290 19190 50920
rect 19160 49280 19220 49290
rect 19160 49210 19220 49220
rect 19160 47580 19190 49210
rect 19160 47570 19220 47580
rect 19160 47500 19220 47510
rect 19040 45860 19100 45870
rect 19040 45790 19100 45800
rect 19040 44160 19070 45790
rect 19040 44150 19100 44160
rect 19040 44080 19100 44090
rect 19040 42450 19070 44080
rect 19040 42440 19100 42450
rect 19040 42370 19100 42380
rect 19040 40740 19070 42370
rect 19040 40730 19100 40740
rect 19040 40660 19100 40670
rect 19040 39240 19070 40660
rect 19160 39300 19190 47500
rect 19280 39690 19310 67050
rect 19400 39690 19430 67050
rect 19520 39690 19550 67050
rect 19640 39690 19670 67050
rect 19760 39690 19790 67050
rect 21920 39690 21950 67050
rect 22040 39690 22070 67050
rect 22160 39690 22190 67050
rect 22280 57840 22310 67050
rect 22400 59550 22430 67050
rect 22520 62970 22550 67050
rect 22640 66390 22670 67050
rect 22610 66380 22670 66390
rect 22610 66310 22670 66320
rect 22640 64680 22670 66310
rect 22610 64670 22670 64680
rect 22610 64600 22670 64610
rect 22490 62960 22550 62970
rect 22490 62890 22550 62900
rect 22520 61250 22550 62890
rect 22490 61240 22550 61250
rect 22490 61170 22550 61180
rect 22370 59540 22430 59550
rect 22370 59470 22430 59480
rect 22250 57830 22310 57840
rect 22250 57760 22310 57770
rect 22280 56130 22310 57760
rect 22250 56120 22310 56130
rect 22250 56050 22310 56060
rect 22280 54420 22310 56050
rect 22250 54410 22310 54420
rect 22250 54340 22310 54350
rect 22280 52710 22310 54340
rect 22250 52700 22310 52710
rect 22250 52630 22310 52640
rect 22280 51000 22310 52630
rect 22250 50990 22310 51000
rect 22250 50920 22310 50930
rect 22280 49290 22310 50920
rect 22250 49280 22310 49290
rect 22250 49210 22310 49220
rect 22280 39420 22310 49210
rect 22400 47580 22430 59470
rect 22370 47570 22430 47580
rect 22370 47500 22430 47510
rect 21870 39410 22310 39420
rect 21930 39390 22310 39410
rect 22400 39360 22430 47500
rect 22520 45870 22550 61170
rect 22490 45860 22550 45870
rect 22490 45790 22550 45800
rect 22520 44160 22550 45790
rect 22490 44150 22550 44160
rect 22490 44080 22550 44090
rect 21870 39340 21930 39350
rect 22050 39350 22430 39360
rect 19160 39290 19480 39300
rect 19160 39270 19420 39290
rect 19040 39230 19300 39240
rect 19040 39210 19240 39230
rect 22110 39330 22430 39350
rect 22520 39300 22550 44080
rect 22640 42450 22670 64600
rect 22610 42440 22670 42450
rect 22610 42370 22670 42380
rect 22640 40740 22670 42370
rect 22610 40730 22670 40740
rect 22610 40660 22670 40670
rect 22050 39280 22110 39290
rect 22230 39290 22550 39300
rect 19420 39220 19480 39230
rect 22290 39270 22550 39290
rect 22640 39240 22670 40660
rect 22700 66470 22770 67050
rect 22700 66210 22720 66470
rect 22760 66210 22770 66470
rect 23780 66470 23850 67050
rect 23230 66440 23310 66450
rect 22920 66402 23120 66408
rect 22810 66370 22890 66390
rect 22810 66310 22820 66370
rect 22880 66358 22890 66370
rect 22920 66368 22932 66402
rect 23108 66400 23120 66402
rect 23230 66400 23240 66440
rect 23108 66380 23240 66400
rect 23300 66400 23310 66440
rect 23418 66402 23618 66408
rect 23418 66400 23430 66402
rect 23300 66380 23430 66400
rect 23108 66370 23430 66380
rect 23108 66368 23120 66370
rect 22920 66362 23120 66368
rect 23418 66368 23430 66370
rect 23606 66368 23618 66402
rect 23418 66362 23618 66368
rect 23650 66370 23730 66390
rect 22882 66324 22890 66358
rect 22880 66310 22890 66324
rect 22810 66290 22890 66310
rect 22920 66314 23120 66320
rect 22920 66280 22932 66314
rect 23108 66310 23120 66314
rect 23418 66314 23618 66320
rect 23418 66310 23430 66314
rect 23108 66280 23430 66310
rect 23606 66280 23618 66314
rect 23650 66310 23660 66370
rect 23720 66310 23730 66370
rect 23650 66290 23730 66310
rect 22920 66274 23120 66280
rect 22700 66150 22770 66210
rect 22700 65910 22720 66150
rect 22760 65910 22770 66150
rect 23230 66270 23310 66280
rect 23418 66274 23618 66280
rect 23230 66210 23240 66270
rect 23300 66210 23310 66270
rect 23230 66160 23310 66210
rect 23230 66100 23240 66160
rect 23300 66100 23310 66160
rect 22920 66092 23120 66098
rect 22810 66060 22890 66080
rect 22810 66000 22820 66060
rect 22880 66048 22890 66060
rect 22920 66058 22932 66092
rect 23108 66090 23120 66092
rect 23230 66090 23310 66100
rect 23780 66230 23790 66470
rect 23830 66230 23850 66470
rect 23780 66150 23850 66230
rect 23418 66092 23618 66098
rect 23418 66090 23430 66092
rect 23108 66060 23430 66090
rect 23108 66058 23120 66060
rect 22920 66052 23120 66058
rect 23418 66058 23430 66060
rect 23606 66058 23618 66092
rect 23418 66052 23618 66058
rect 23650 66060 23730 66080
rect 22882 66014 22890 66048
rect 22880 66000 22890 66014
rect 22810 65980 22890 66000
rect 22920 66004 23120 66010
rect 22920 65970 22932 66004
rect 23108 66000 23120 66004
rect 23418 66004 23618 66010
rect 23418 66000 23430 66004
rect 23108 65990 23430 66000
rect 23108 65970 23240 65990
rect 22920 65964 23120 65970
rect 23230 65930 23240 65970
rect 23300 65970 23430 65990
rect 23606 65970 23618 66004
rect 23650 66000 23660 66060
rect 23720 66000 23730 66060
rect 23650 65980 23730 66000
rect 23300 65930 23310 65970
rect 23418 65964 23618 65970
rect 23230 65920 23310 65930
rect 22700 64760 22770 65910
rect 22700 64500 22720 64760
rect 22760 64500 22770 64760
rect 23780 65910 23790 66150
rect 23830 65910 23850 66150
rect 23780 64760 23850 65910
rect 23230 64730 23310 64740
rect 22920 64692 23120 64698
rect 22810 64660 22890 64680
rect 22810 64600 22820 64660
rect 22880 64648 22890 64660
rect 22920 64658 22932 64692
rect 23108 64690 23120 64692
rect 23230 64690 23240 64730
rect 23108 64670 23240 64690
rect 23300 64690 23310 64730
rect 23418 64692 23618 64698
rect 23418 64690 23430 64692
rect 23300 64670 23430 64690
rect 23108 64660 23430 64670
rect 23108 64658 23120 64660
rect 22920 64652 23120 64658
rect 23418 64658 23430 64660
rect 23606 64658 23618 64692
rect 23418 64652 23618 64658
rect 23650 64660 23730 64680
rect 22882 64614 22890 64648
rect 22880 64600 22890 64614
rect 22810 64580 22890 64600
rect 22920 64604 23120 64610
rect 22920 64570 22932 64604
rect 23108 64600 23120 64604
rect 23418 64604 23618 64610
rect 23418 64600 23430 64604
rect 23108 64570 23430 64600
rect 23606 64570 23618 64604
rect 23650 64600 23660 64660
rect 23720 64600 23730 64660
rect 23650 64580 23730 64600
rect 22920 64564 23120 64570
rect 22700 64440 22770 64500
rect 22700 64200 22720 64440
rect 22760 64200 22770 64440
rect 23230 64560 23310 64570
rect 23418 64564 23618 64570
rect 23230 64500 23240 64560
rect 23300 64500 23310 64560
rect 23230 64450 23310 64500
rect 23230 64390 23240 64450
rect 23300 64390 23310 64450
rect 22920 64382 23120 64388
rect 22810 64350 22890 64370
rect 22810 64290 22820 64350
rect 22880 64338 22890 64350
rect 22920 64348 22932 64382
rect 23108 64380 23120 64382
rect 23230 64380 23310 64390
rect 23780 64520 23790 64760
rect 23830 64520 23850 64760
rect 23780 64440 23850 64520
rect 23418 64382 23618 64388
rect 23418 64380 23430 64382
rect 23108 64350 23430 64380
rect 23108 64348 23120 64350
rect 22920 64342 23120 64348
rect 23418 64348 23430 64350
rect 23606 64348 23618 64382
rect 23418 64342 23618 64348
rect 23650 64350 23730 64370
rect 22882 64304 22890 64338
rect 22880 64290 22890 64304
rect 22810 64270 22890 64290
rect 22920 64294 23120 64300
rect 22920 64260 22932 64294
rect 23108 64290 23120 64294
rect 23418 64294 23618 64300
rect 23418 64290 23430 64294
rect 23108 64280 23430 64290
rect 23108 64260 23240 64280
rect 22920 64254 23120 64260
rect 23230 64220 23240 64260
rect 23300 64260 23430 64280
rect 23606 64260 23618 64294
rect 23650 64290 23660 64350
rect 23720 64290 23730 64350
rect 23650 64270 23730 64290
rect 23300 64220 23310 64260
rect 23418 64254 23618 64260
rect 23230 64210 23310 64220
rect 22700 63050 22770 64200
rect 22700 62790 22720 63050
rect 22760 62790 22770 63050
rect 23780 64200 23790 64440
rect 23830 64200 23850 64440
rect 23780 63050 23850 64200
rect 23230 63020 23310 63030
rect 22920 62982 23120 62988
rect 22810 62950 22890 62970
rect 22810 62890 22820 62950
rect 22880 62938 22890 62950
rect 22920 62948 22932 62982
rect 23108 62980 23120 62982
rect 23230 62980 23240 63020
rect 23108 62960 23240 62980
rect 23300 62980 23310 63020
rect 23418 62982 23618 62988
rect 23418 62980 23430 62982
rect 23300 62960 23430 62980
rect 23108 62950 23430 62960
rect 23108 62948 23120 62950
rect 22920 62942 23120 62948
rect 23418 62948 23430 62950
rect 23606 62948 23618 62982
rect 23418 62942 23618 62948
rect 23650 62950 23730 62970
rect 22882 62904 22890 62938
rect 22880 62890 22890 62904
rect 22810 62870 22890 62890
rect 22920 62894 23120 62900
rect 22920 62860 22932 62894
rect 23108 62890 23120 62894
rect 23418 62894 23618 62900
rect 23418 62890 23430 62894
rect 23108 62860 23430 62890
rect 23606 62860 23618 62894
rect 23650 62890 23660 62950
rect 23720 62890 23730 62950
rect 23650 62870 23730 62890
rect 22920 62854 23120 62860
rect 22700 62730 22770 62790
rect 22700 62490 22720 62730
rect 22760 62490 22770 62730
rect 23230 62850 23310 62860
rect 23418 62854 23618 62860
rect 23230 62790 23240 62850
rect 23300 62790 23310 62850
rect 23230 62740 23310 62790
rect 23230 62680 23240 62740
rect 23300 62680 23310 62740
rect 22920 62672 23120 62678
rect 22810 62640 22890 62660
rect 22810 62580 22820 62640
rect 22880 62628 22890 62640
rect 22920 62638 22932 62672
rect 23108 62670 23120 62672
rect 23230 62670 23310 62680
rect 23780 62810 23790 63050
rect 23830 62810 23850 63050
rect 23780 62730 23850 62810
rect 23418 62672 23618 62678
rect 23418 62670 23430 62672
rect 23108 62640 23430 62670
rect 23108 62638 23120 62640
rect 22920 62632 23120 62638
rect 23418 62638 23430 62640
rect 23606 62638 23618 62672
rect 23418 62632 23618 62638
rect 23650 62640 23730 62660
rect 22882 62594 22890 62628
rect 22880 62580 22890 62594
rect 22810 62560 22890 62580
rect 22920 62584 23120 62590
rect 22920 62550 22932 62584
rect 23108 62580 23120 62584
rect 23418 62584 23618 62590
rect 23418 62580 23430 62584
rect 23108 62570 23430 62580
rect 23108 62550 23240 62570
rect 22920 62544 23120 62550
rect 23230 62510 23240 62550
rect 23300 62550 23430 62570
rect 23606 62550 23618 62584
rect 23650 62580 23660 62640
rect 23720 62580 23730 62640
rect 23650 62560 23730 62580
rect 23300 62510 23310 62550
rect 23418 62544 23618 62550
rect 23230 62500 23310 62510
rect 22700 61340 22770 62490
rect 22700 61080 22720 61340
rect 22760 61080 22770 61340
rect 23780 62490 23790 62730
rect 23830 62490 23850 62730
rect 23780 61340 23850 62490
rect 23230 61310 23310 61320
rect 22920 61272 23120 61278
rect 22810 61240 22890 61260
rect 22810 61180 22820 61240
rect 22880 61228 22890 61240
rect 22920 61238 22932 61272
rect 23108 61270 23120 61272
rect 23230 61270 23240 61310
rect 23108 61250 23240 61270
rect 23300 61270 23310 61310
rect 23418 61272 23618 61278
rect 23418 61270 23430 61272
rect 23300 61250 23430 61270
rect 23108 61240 23430 61250
rect 23108 61238 23120 61240
rect 22920 61232 23120 61238
rect 23418 61238 23430 61240
rect 23606 61238 23618 61272
rect 23418 61232 23618 61238
rect 23650 61240 23730 61260
rect 22882 61194 22890 61228
rect 22880 61180 22890 61194
rect 22810 61160 22890 61180
rect 22920 61184 23120 61190
rect 22920 61150 22932 61184
rect 23108 61180 23120 61184
rect 23418 61184 23618 61190
rect 23418 61180 23430 61184
rect 23108 61150 23430 61180
rect 23606 61150 23618 61184
rect 23650 61180 23660 61240
rect 23720 61180 23730 61240
rect 23650 61160 23730 61180
rect 22920 61144 23120 61150
rect 22700 61020 22770 61080
rect 22700 60780 22720 61020
rect 22760 60780 22770 61020
rect 23230 61140 23310 61150
rect 23418 61144 23618 61150
rect 23230 61080 23240 61140
rect 23300 61080 23310 61140
rect 23230 61030 23310 61080
rect 23230 60970 23240 61030
rect 23300 60970 23310 61030
rect 22920 60962 23120 60968
rect 22810 60930 22890 60950
rect 22810 60870 22820 60930
rect 22880 60918 22890 60930
rect 22920 60928 22932 60962
rect 23108 60960 23120 60962
rect 23230 60960 23310 60970
rect 23780 61100 23790 61340
rect 23830 61100 23850 61340
rect 23780 61020 23850 61100
rect 23418 60962 23618 60968
rect 23418 60960 23430 60962
rect 23108 60930 23430 60960
rect 23108 60928 23120 60930
rect 22920 60922 23120 60928
rect 23418 60928 23430 60930
rect 23606 60928 23618 60962
rect 23418 60922 23618 60928
rect 23650 60930 23730 60950
rect 22882 60884 22890 60918
rect 22880 60870 22890 60884
rect 22810 60850 22890 60870
rect 22920 60874 23120 60880
rect 22920 60840 22932 60874
rect 23108 60870 23120 60874
rect 23418 60874 23618 60880
rect 23418 60870 23430 60874
rect 23108 60860 23430 60870
rect 23108 60840 23240 60860
rect 22920 60834 23120 60840
rect 23230 60800 23240 60840
rect 23300 60840 23430 60860
rect 23606 60840 23618 60874
rect 23650 60870 23660 60930
rect 23720 60870 23730 60930
rect 23650 60850 23730 60870
rect 23300 60800 23310 60840
rect 23418 60834 23618 60840
rect 23230 60790 23310 60800
rect 22700 59630 22770 60780
rect 22700 59370 22720 59630
rect 22760 59370 22770 59630
rect 23780 60780 23790 61020
rect 23830 60780 23850 61020
rect 23780 59630 23850 60780
rect 23230 59600 23310 59610
rect 22920 59562 23120 59568
rect 22810 59530 22890 59550
rect 22810 59470 22820 59530
rect 22880 59518 22890 59530
rect 22920 59528 22932 59562
rect 23108 59560 23120 59562
rect 23230 59560 23240 59600
rect 23108 59540 23240 59560
rect 23300 59560 23310 59600
rect 23418 59562 23618 59568
rect 23418 59560 23430 59562
rect 23300 59540 23430 59560
rect 23108 59530 23430 59540
rect 23108 59528 23120 59530
rect 22920 59522 23120 59528
rect 23418 59528 23430 59530
rect 23606 59528 23618 59562
rect 23418 59522 23618 59528
rect 23650 59530 23730 59550
rect 22882 59484 22890 59518
rect 22880 59470 22890 59484
rect 22810 59450 22890 59470
rect 22920 59474 23120 59480
rect 22920 59440 22932 59474
rect 23108 59470 23120 59474
rect 23418 59474 23618 59480
rect 23418 59470 23430 59474
rect 23108 59440 23430 59470
rect 23606 59440 23618 59474
rect 23650 59470 23660 59530
rect 23720 59470 23730 59530
rect 23650 59450 23730 59470
rect 22920 59434 23120 59440
rect 22700 59310 22770 59370
rect 22700 59070 22720 59310
rect 22760 59070 22770 59310
rect 23230 59430 23310 59440
rect 23418 59434 23618 59440
rect 23230 59370 23240 59430
rect 23300 59370 23310 59430
rect 23230 59320 23310 59370
rect 23230 59260 23240 59320
rect 23300 59260 23310 59320
rect 22920 59252 23120 59258
rect 22810 59220 22890 59240
rect 22810 59160 22820 59220
rect 22880 59208 22890 59220
rect 22920 59218 22932 59252
rect 23108 59250 23120 59252
rect 23230 59250 23310 59260
rect 23780 59390 23790 59630
rect 23830 59390 23850 59630
rect 23780 59310 23850 59390
rect 23418 59252 23618 59258
rect 23418 59250 23430 59252
rect 23108 59220 23430 59250
rect 23108 59218 23120 59220
rect 22920 59212 23120 59218
rect 23418 59218 23430 59220
rect 23606 59218 23618 59252
rect 23418 59212 23618 59218
rect 23650 59220 23730 59240
rect 22882 59174 22890 59208
rect 22880 59160 22890 59174
rect 22810 59140 22890 59160
rect 22920 59164 23120 59170
rect 22920 59130 22932 59164
rect 23108 59160 23120 59164
rect 23418 59164 23618 59170
rect 23418 59160 23430 59164
rect 23108 59150 23430 59160
rect 23108 59130 23240 59150
rect 22920 59124 23120 59130
rect 23230 59090 23240 59130
rect 23300 59130 23430 59150
rect 23606 59130 23618 59164
rect 23650 59160 23660 59220
rect 23720 59160 23730 59220
rect 23650 59140 23730 59160
rect 23300 59090 23310 59130
rect 23418 59124 23618 59130
rect 23230 59080 23310 59090
rect 22700 57920 22770 59070
rect 22700 57660 22720 57920
rect 22760 57660 22770 57920
rect 23780 59070 23790 59310
rect 23830 59070 23850 59310
rect 23780 57920 23850 59070
rect 23230 57890 23310 57900
rect 22920 57852 23120 57858
rect 22810 57820 22890 57840
rect 22810 57760 22820 57820
rect 22880 57808 22890 57820
rect 22920 57818 22932 57852
rect 23108 57850 23120 57852
rect 23230 57850 23240 57890
rect 23108 57830 23240 57850
rect 23300 57850 23310 57890
rect 23418 57852 23618 57858
rect 23418 57850 23430 57852
rect 23300 57830 23430 57850
rect 23108 57820 23430 57830
rect 23108 57818 23120 57820
rect 22920 57812 23120 57818
rect 23418 57818 23430 57820
rect 23606 57818 23618 57852
rect 23418 57812 23618 57818
rect 23650 57820 23730 57840
rect 22882 57774 22890 57808
rect 22880 57760 22890 57774
rect 22810 57740 22890 57760
rect 22920 57764 23120 57770
rect 22920 57730 22932 57764
rect 23108 57760 23120 57764
rect 23418 57764 23618 57770
rect 23418 57760 23430 57764
rect 23108 57730 23430 57760
rect 23606 57730 23618 57764
rect 23650 57760 23660 57820
rect 23720 57760 23730 57820
rect 23650 57740 23730 57760
rect 22920 57724 23120 57730
rect 22700 57600 22770 57660
rect 22700 57360 22720 57600
rect 22760 57360 22770 57600
rect 23230 57720 23310 57730
rect 23418 57724 23618 57730
rect 23230 57660 23240 57720
rect 23300 57660 23310 57720
rect 23230 57610 23310 57660
rect 23230 57550 23240 57610
rect 23300 57550 23310 57610
rect 22920 57542 23120 57548
rect 22810 57510 22890 57530
rect 22810 57450 22820 57510
rect 22880 57498 22890 57510
rect 22920 57508 22932 57542
rect 23108 57540 23120 57542
rect 23230 57540 23310 57550
rect 23780 57680 23790 57920
rect 23830 57680 23850 57920
rect 23780 57600 23850 57680
rect 23418 57542 23618 57548
rect 23418 57540 23430 57542
rect 23108 57510 23430 57540
rect 23108 57508 23120 57510
rect 22920 57502 23120 57508
rect 23418 57508 23430 57510
rect 23606 57508 23618 57542
rect 23418 57502 23618 57508
rect 23650 57510 23730 57530
rect 22882 57464 22890 57498
rect 22880 57450 22890 57464
rect 22810 57430 22890 57450
rect 22920 57454 23120 57460
rect 22920 57420 22932 57454
rect 23108 57450 23120 57454
rect 23418 57454 23618 57460
rect 23418 57450 23430 57454
rect 23108 57440 23430 57450
rect 23108 57420 23240 57440
rect 22920 57414 23120 57420
rect 23230 57380 23240 57420
rect 23300 57420 23430 57440
rect 23606 57420 23618 57454
rect 23650 57450 23660 57510
rect 23720 57450 23730 57510
rect 23650 57430 23730 57450
rect 23300 57380 23310 57420
rect 23418 57414 23618 57420
rect 23230 57370 23310 57380
rect 22700 56210 22770 57360
rect 22700 55950 22720 56210
rect 22760 55950 22770 56210
rect 23780 57360 23790 57600
rect 23830 57360 23850 57600
rect 23780 56210 23850 57360
rect 23230 56180 23310 56190
rect 22920 56142 23120 56148
rect 22810 56110 22890 56130
rect 22810 56050 22820 56110
rect 22880 56098 22890 56110
rect 22920 56108 22932 56142
rect 23108 56140 23120 56142
rect 23230 56140 23240 56180
rect 23108 56120 23240 56140
rect 23300 56140 23310 56180
rect 23418 56142 23618 56148
rect 23418 56140 23430 56142
rect 23300 56120 23430 56140
rect 23108 56110 23430 56120
rect 23108 56108 23120 56110
rect 22920 56102 23120 56108
rect 23418 56108 23430 56110
rect 23606 56108 23618 56142
rect 23418 56102 23618 56108
rect 23650 56110 23730 56130
rect 22882 56064 22890 56098
rect 22880 56050 22890 56064
rect 22810 56030 22890 56050
rect 22920 56054 23120 56060
rect 22920 56020 22932 56054
rect 23108 56050 23120 56054
rect 23418 56054 23618 56060
rect 23418 56050 23430 56054
rect 23108 56020 23430 56050
rect 23606 56020 23618 56054
rect 23650 56050 23660 56110
rect 23720 56050 23730 56110
rect 23650 56030 23730 56050
rect 22920 56014 23120 56020
rect 22700 55890 22770 55950
rect 22700 55650 22720 55890
rect 22760 55650 22770 55890
rect 23230 56010 23310 56020
rect 23418 56014 23618 56020
rect 23230 55950 23240 56010
rect 23300 55950 23310 56010
rect 23230 55900 23310 55950
rect 23230 55840 23240 55900
rect 23300 55840 23310 55900
rect 22920 55832 23120 55838
rect 22810 55800 22890 55820
rect 22810 55740 22820 55800
rect 22880 55788 22890 55800
rect 22920 55798 22932 55832
rect 23108 55830 23120 55832
rect 23230 55830 23310 55840
rect 23780 55970 23790 56210
rect 23830 55970 23850 56210
rect 23780 55890 23850 55970
rect 23418 55832 23618 55838
rect 23418 55830 23430 55832
rect 23108 55800 23430 55830
rect 23108 55798 23120 55800
rect 22920 55792 23120 55798
rect 23418 55798 23430 55800
rect 23606 55798 23618 55832
rect 23418 55792 23618 55798
rect 23650 55800 23730 55820
rect 22882 55754 22890 55788
rect 22880 55740 22890 55754
rect 22810 55720 22890 55740
rect 22920 55744 23120 55750
rect 22920 55710 22932 55744
rect 23108 55740 23120 55744
rect 23418 55744 23618 55750
rect 23418 55740 23430 55744
rect 23108 55730 23430 55740
rect 23108 55710 23240 55730
rect 22920 55704 23120 55710
rect 23230 55670 23240 55710
rect 23300 55710 23430 55730
rect 23606 55710 23618 55744
rect 23650 55740 23660 55800
rect 23720 55740 23730 55800
rect 23650 55720 23730 55740
rect 23300 55670 23310 55710
rect 23418 55704 23618 55710
rect 23230 55660 23310 55670
rect 22700 54500 22770 55650
rect 22700 54240 22720 54500
rect 22760 54240 22770 54500
rect 23780 55650 23790 55890
rect 23830 55650 23850 55890
rect 23780 54500 23850 55650
rect 23230 54470 23310 54480
rect 22920 54432 23120 54438
rect 22810 54400 22890 54420
rect 22810 54340 22820 54400
rect 22880 54388 22890 54400
rect 22920 54398 22932 54432
rect 23108 54430 23120 54432
rect 23230 54430 23240 54470
rect 23108 54410 23240 54430
rect 23300 54430 23310 54470
rect 23418 54432 23618 54438
rect 23418 54430 23430 54432
rect 23300 54410 23430 54430
rect 23108 54400 23430 54410
rect 23108 54398 23120 54400
rect 22920 54392 23120 54398
rect 23418 54398 23430 54400
rect 23606 54398 23618 54432
rect 23418 54392 23618 54398
rect 23650 54400 23730 54420
rect 22882 54354 22890 54388
rect 22880 54340 22890 54354
rect 22810 54320 22890 54340
rect 22920 54344 23120 54350
rect 22920 54310 22932 54344
rect 23108 54340 23120 54344
rect 23418 54344 23618 54350
rect 23418 54340 23430 54344
rect 23108 54310 23430 54340
rect 23606 54310 23618 54344
rect 23650 54340 23660 54400
rect 23720 54340 23730 54400
rect 23650 54320 23730 54340
rect 22920 54304 23120 54310
rect 22700 54180 22770 54240
rect 22700 53940 22720 54180
rect 22760 53940 22770 54180
rect 23230 54300 23310 54310
rect 23418 54304 23618 54310
rect 23230 54240 23240 54300
rect 23300 54240 23310 54300
rect 23230 54190 23310 54240
rect 23230 54130 23240 54190
rect 23300 54130 23310 54190
rect 22920 54122 23120 54128
rect 22810 54090 22890 54110
rect 22810 54030 22820 54090
rect 22880 54078 22890 54090
rect 22920 54088 22932 54122
rect 23108 54120 23120 54122
rect 23230 54120 23310 54130
rect 23780 54260 23790 54500
rect 23830 54260 23850 54500
rect 23780 54180 23850 54260
rect 23418 54122 23618 54128
rect 23418 54120 23430 54122
rect 23108 54090 23430 54120
rect 23108 54088 23120 54090
rect 22920 54082 23120 54088
rect 23418 54088 23430 54090
rect 23606 54088 23618 54122
rect 23418 54082 23618 54088
rect 23650 54090 23730 54110
rect 22882 54044 22890 54078
rect 22880 54030 22890 54044
rect 22810 54010 22890 54030
rect 22920 54034 23120 54040
rect 22920 54000 22932 54034
rect 23108 54030 23120 54034
rect 23418 54034 23618 54040
rect 23418 54030 23430 54034
rect 23108 54020 23430 54030
rect 23108 54000 23240 54020
rect 22920 53994 23120 54000
rect 23230 53960 23240 54000
rect 23300 54000 23430 54020
rect 23606 54000 23618 54034
rect 23650 54030 23660 54090
rect 23720 54030 23730 54090
rect 23650 54010 23730 54030
rect 23300 53960 23310 54000
rect 23418 53994 23618 54000
rect 23230 53950 23310 53960
rect 22700 52790 22770 53940
rect 22700 52530 22720 52790
rect 22760 52530 22770 52790
rect 23780 53940 23790 54180
rect 23830 53940 23850 54180
rect 23780 52790 23850 53940
rect 23230 52760 23310 52770
rect 22920 52722 23120 52728
rect 22810 52690 22890 52710
rect 22810 52630 22820 52690
rect 22880 52678 22890 52690
rect 22920 52688 22932 52722
rect 23108 52720 23120 52722
rect 23230 52720 23240 52760
rect 23108 52700 23240 52720
rect 23300 52720 23310 52760
rect 23418 52722 23618 52728
rect 23418 52720 23430 52722
rect 23300 52700 23430 52720
rect 23108 52690 23430 52700
rect 23108 52688 23120 52690
rect 22920 52682 23120 52688
rect 23418 52688 23430 52690
rect 23606 52688 23618 52722
rect 23418 52682 23618 52688
rect 23650 52690 23730 52710
rect 22882 52644 22890 52678
rect 22880 52630 22890 52644
rect 22810 52610 22890 52630
rect 22920 52634 23120 52640
rect 22920 52600 22932 52634
rect 23108 52630 23120 52634
rect 23418 52634 23618 52640
rect 23418 52630 23430 52634
rect 23108 52600 23430 52630
rect 23606 52600 23618 52634
rect 23650 52630 23660 52690
rect 23720 52630 23730 52690
rect 23650 52610 23730 52630
rect 22920 52594 23120 52600
rect 22700 52470 22770 52530
rect 22700 52230 22720 52470
rect 22760 52230 22770 52470
rect 23230 52590 23310 52600
rect 23418 52594 23618 52600
rect 23230 52530 23240 52590
rect 23300 52530 23310 52590
rect 23230 52480 23310 52530
rect 23230 52420 23240 52480
rect 23300 52420 23310 52480
rect 22920 52412 23120 52418
rect 22810 52380 22890 52400
rect 22810 52320 22820 52380
rect 22880 52368 22890 52380
rect 22920 52378 22932 52412
rect 23108 52410 23120 52412
rect 23230 52410 23310 52420
rect 23780 52550 23790 52790
rect 23830 52550 23850 52790
rect 23780 52470 23850 52550
rect 23418 52412 23618 52418
rect 23418 52410 23430 52412
rect 23108 52380 23430 52410
rect 23108 52378 23120 52380
rect 22920 52372 23120 52378
rect 23418 52378 23430 52380
rect 23606 52378 23618 52412
rect 23418 52372 23618 52378
rect 23650 52380 23730 52400
rect 22882 52334 22890 52368
rect 22880 52320 22890 52334
rect 22810 52300 22890 52320
rect 22920 52324 23120 52330
rect 22920 52290 22932 52324
rect 23108 52320 23120 52324
rect 23418 52324 23618 52330
rect 23418 52320 23430 52324
rect 23108 52310 23430 52320
rect 23108 52290 23240 52310
rect 22920 52284 23120 52290
rect 23230 52250 23240 52290
rect 23300 52290 23430 52310
rect 23606 52290 23618 52324
rect 23650 52320 23660 52380
rect 23720 52320 23730 52380
rect 23650 52300 23730 52320
rect 23300 52250 23310 52290
rect 23418 52284 23618 52290
rect 23230 52240 23310 52250
rect 22700 51080 22770 52230
rect 22700 50820 22720 51080
rect 22760 50820 22770 51080
rect 23780 52230 23790 52470
rect 23830 52230 23850 52470
rect 23780 51080 23850 52230
rect 23230 51050 23310 51060
rect 22920 51012 23120 51018
rect 22810 50980 22890 51000
rect 22810 50920 22820 50980
rect 22880 50968 22890 50980
rect 22920 50978 22932 51012
rect 23108 51010 23120 51012
rect 23230 51010 23240 51050
rect 23108 50990 23240 51010
rect 23300 51010 23310 51050
rect 23418 51012 23618 51018
rect 23418 51010 23430 51012
rect 23300 50990 23430 51010
rect 23108 50980 23430 50990
rect 23108 50978 23120 50980
rect 22920 50972 23120 50978
rect 23418 50978 23430 50980
rect 23606 50978 23618 51012
rect 23418 50972 23618 50978
rect 23650 50980 23730 51000
rect 22882 50934 22890 50968
rect 22880 50920 22890 50934
rect 22810 50900 22890 50920
rect 22920 50924 23120 50930
rect 22920 50890 22932 50924
rect 23108 50920 23120 50924
rect 23418 50924 23618 50930
rect 23418 50920 23430 50924
rect 23108 50890 23430 50920
rect 23606 50890 23618 50924
rect 23650 50920 23660 50980
rect 23720 50920 23730 50980
rect 23650 50900 23730 50920
rect 22920 50884 23120 50890
rect 22700 50760 22770 50820
rect 22700 50520 22720 50760
rect 22760 50520 22770 50760
rect 23230 50880 23310 50890
rect 23418 50884 23618 50890
rect 23230 50820 23240 50880
rect 23300 50820 23310 50880
rect 23230 50770 23310 50820
rect 23230 50710 23240 50770
rect 23300 50710 23310 50770
rect 22920 50702 23120 50708
rect 22810 50670 22890 50690
rect 22810 50610 22820 50670
rect 22880 50658 22890 50670
rect 22920 50668 22932 50702
rect 23108 50700 23120 50702
rect 23230 50700 23310 50710
rect 23780 50840 23790 51080
rect 23830 50840 23850 51080
rect 23780 50760 23850 50840
rect 23418 50702 23618 50708
rect 23418 50700 23430 50702
rect 23108 50670 23430 50700
rect 23108 50668 23120 50670
rect 22920 50662 23120 50668
rect 23418 50668 23430 50670
rect 23606 50668 23618 50702
rect 23418 50662 23618 50668
rect 23650 50670 23730 50690
rect 22882 50624 22890 50658
rect 22880 50610 22890 50624
rect 22810 50590 22890 50610
rect 22920 50614 23120 50620
rect 22920 50580 22932 50614
rect 23108 50610 23120 50614
rect 23418 50614 23618 50620
rect 23418 50610 23430 50614
rect 23108 50600 23430 50610
rect 23108 50580 23240 50600
rect 22920 50574 23120 50580
rect 23230 50540 23240 50580
rect 23300 50580 23430 50600
rect 23606 50580 23618 50614
rect 23650 50610 23660 50670
rect 23720 50610 23730 50670
rect 23650 50590 23730 50610
rect 23300 50540 23310 50580
rect 23418 50574 23618 50580
rect 23230 50530 23310 50540
rect 22700 49370 22770 50520
rect 22700 49110 22720 49370
rect 22760 49110 22770 49370
rect 23780 50520 23790 50760
rect 23830 50520 23850 50760
rect 23780 49370 23850 50520
rect 23230 49340 23310 49350
rect 22920 49302 23120 49308
rect 22810 49270 22890 49290
rect 22810 49210 22820 49270
rect 22880 49258 22890 49270
rect 22920 49268 22932 49302
rect 23108 49300 23120 49302
rect 23230 49300 23240 49340
rect 23108 49280 23240 49300
rect 23300 49300 23310 49340
rect 23418 49302 23618 49308
rect 23418 49300 23430 49302
rect 23300 49280 23430 49300
rect 23108 49270 23430 49280
rect 23108 49268 23120 49270
rect 22920 49262 23120 49268
rect 23418 49268 23430 49270
rect 23606 49268 23618 49302
rect 23418 49262 23618 49268
rect 23650 49270 23730 49290
rect 22882 49224 22890 49258
rect 22880 49210 22890 49224
rect 22810 49190 22890 49210
rect 22920 49214 23120 49220
rect 22920 49180 22932 49214
rect 23108 49210 23120 49214
rect 23418 49214 23618 49220
rect 23418 49210 23430 49214
rect 23108 49180 23430 49210
rect 23606 49180 23618 49214
rect 23650 49210 23660 49270
rect 23720 49210 23730 49270
rect 23650 49190 23730 49210
rect 22920 49174 23120 49180
rect 22700 49050 22770 49110
rect 22700 48810 22720 49050
rect 22760 48810 22770 49050
rect 23230 49170 23310 49180
rect 23418 49174 23618 49180
rect 23230 49110 23240 49170
rect 23300 49110 23310 49170
rect 23230 49060 23310 49110
rect 23230 49000 23240 49060
rect 23300 49000 23310 49060
rect 22920 48992 23120 48998
rect 22810 48960 22890 48980
rect 22810 48900 22820 48960
rect 22880 48948 22890 48960
rect 22920 48958 22932 48992
rect 23108 48990 23120 48992
rect 23230 48990 23310 49000
rect 23780 49130 23790 49370
rect 23830 49130 23850 49370
rect 23780 49050 23850 49130
rect 23418 48992 23618 48998
rect 23418 48990 23430 48992
rect 23108 48960 23430 48990
rect 23108 48958 23120 48960
rect 22920 48952 23120 48958
rect 23418 48958 23430 48960
rect 23606 48958 23618 48992
rect 23418 48952 23618 48958
rect 23650 48960 23730 48980
rect 22882 48914 22890 48948
rect 22880 48900 22890 48914
rect 22810 48880 22890 48900
rect 22920 48904 23120 48910
rect 22920 48870 22932 48904
rect 23108 48900 23120 48904
rect 23418 48904 23618 48910
rect 23418 48900 23430 48904
rect 23108 48890 23430 48900
rect 23108 48870 23240 48890
rect 22920 48864 23120 48870
rect 23230 48830 23240 48870
rect 23300 48870 23430 48890
rect 23606 48870 23618 48904
rect 23650 48900 23660 48960
rect 23720 48900 23730 48960
rect 23650 48880 23730 48900
rect 23300 48830 23310 48870
rect 23418 48864 23618 48870
rect 23230 48820 23310 48830
rect 22700 47660 22770 48810
rect 22700 47400 22720 47660
rect 22760 47400 22770 47660
rect 23780 48810 23790 49050
rect 23830 48810 23850 49050
rect 23780 47660 23850 48810
rect 23230 47630 23310 47640
rect 22920 47592 23120 47598
rect 22810 47560 22890 47580
rect 22810 47500 22820 47560
rect 22880 47548 22890 47560
rect 22920 47558 22932 47592
rect 23108 47590 23120 47592
rect 23230 47590 23240 47630
rect 23108 47570 23240 47590
rect 23300 47590 23310 47630
rect 23418 47592 23618 47598
rect 23418 47590 23430 47592
rect 23300 47570 23430 47590
rect 23108 47560 23430 47570
rect 23108 47558 23120 47560
rect 22920 47552 23120 47558
rect 23418 47558 23430 47560
rect 23606 47558 23618 47592
rect 23418 47552 23618 47558
rect 23650 47560 23730 47580
rect 22882 47514 22890 47548
rect 22880 47500 22890 47514
rect 22810 47480 22890 47500
rect 22920 47504 23120 47510
rect 22920 47470 22932 47504
rect 23108 47500 23120 47504
rect 23418 47504 23618 47510
rect 23418 47500 23430 47504
rect 23108 47470 23430 47500
rect 23606 47470 23618 47504
rect 23650 47500 23660 47560
rect 23720 47500 23730 47560
rect 23650 47480 23730 47500
rect 22920 47464 23120 47470
rect 22700 47340 22770 47400
rect 22700 47100 22720 47340
rect 22760 47100 22770 47340
rect 23230 47460 23310 47470
rect 23418 47464 23618 47470
rect 23230 47400 23240 47460
rect 23300 47400 23310 47460
rect 23230 47350 23310 47400
rect 23230 47290 23240 47350
rect 23300 47290 23310 47350
rect 22920 47282 23120 47288
rect 22810 47250 22890 47270
rect 22810 47190 22820 47250
rect 22880 47238 22890 47250
rect 22920 47248 22932 47282
rect 23108 47280 23120 47282
rect 23230 47280 23310 47290
rect 23780 47420 23790 47660
rect 23830 47420 23850 47660
rect 23780 47340 23850 47420
rect 23418 47282 23618 47288
rect 23418 47280 23430 47282
rect 23108 47250 23430 47280
rect 23108 47248 23120 47250
rect 22920 47242 23120 47248
rect 23418 47248 23430 47250
rect 23606 47248 23618 47282
rect 23418 47242 23618 47248
rect 23650 47250 23730 47270
rect 22882 47204 22890 47238
rect 22880 47190 22890 47204
rect 22810 47170 22890 47190
rect 22920 47194 23120 47200
rect 22920 47160 22932 47194
rect 23108 47190 23120 47194
rect 23418 47194 23618 47200
rect 23418 47190 23430 47194
rect 23108 47180 23430 47190
rect 23108 47160 23240 47180
rect 22920 47154 23120 47160
rect 23230 47120 23240 47160
rect 23300 47160 23430 47180
rect 23606 47160 23618 47194
rect 23650 47190 23660 47250
rect 23720 47190 23730 47250
rect 23650 47170 23730 47190
rect 23300 47120 23310 47160
rect 23418 47154 23618 47160
rect 23230 47110 23310 47120
rect 22700 45950 22770 47100
rect 22700 45690 22720 45950
rect 22760 45690 22770 45950
rect 23780 47100 23790 47340
rect 23830 47100 23850 47340
rect 23780 45950 23850 47100
rect 23230 45920 23310 45930
rect 22920 45882 23120 45888
rect 22810 45850 22890 45870
rect 22810 45790 22820 45850
rect 22880 45838 22890 45850
rect 22920 45848 22932 45882
rect 23108 45880 23120 45882
rect 23230 45880 23240 45920
rect 23108 45860 23240 45880
rect 23300 45880 23310 45920
rect 23418 45882 23618 45888
rect 23418 45880 23430 45882
rect 23300 45860 23430 45880
rect 23108 45850 23430 45860
rect 23108 45848 23120 45850
rect 22920 45842 23120 45848
rect 23418 45848 23430 45850
rect 23606 45848 23618 45882
rect 23418 45842 23618 45848
rect 23650 45850 23730 45870
rect 22882 45804 22890 45838
rect 22880 45790 22890 45804
rect 22810 45770 22890 45790
rect 22920 45794 23120 45800
rect 22920 45760 22932 45794
rect 23108 45790 23120 45794
rect 23418 45794 23618 45800
rect 23418 45790 23430 45794
rect 23108 45760 23430 45790
rect 23606 45760 23618 45794
rect 23650 45790 23660 45850
rect 23720 45790 23730 45850
rect 23650 45770 23730 45790
rect 22920 45754 23120 45760
rect 22700 45630 22770 45690
rect 22700 45390 22720 45630
rect 22760 45390 22770 45630
rect 23230 45750 23310 45760
rect 23418 45754 23618 45760
rect 23230 45690 23240 45750
rect 23300 45690 23310 45750
rect 23230 45640 23310 45690
rect 23230 45580 23240 45640
rect 23300 45580 23310 45640
rect 22920 45572 23120 45578
rect 22810 45540 22890 45560
rect 22810 45480 22820 45540
rect 22880 45528 22890 45540
rect 22920 45538 22932 45572
rect 23108 45570 23120 45572
rect 23230 45570 23310 45580
rect 23780 45710 23790 45950
rect 23830 45710 23850 45950
rect 23780 45630 23850 45710
rect 23418 45572 23618 45578
rect 23418 45570 23430 45572
rect 23108 45540 23430 45570
rect 23108 45538 23120 45540
rect 22920 45532 23120 45538
rect 23418 45538 23430 45540
rect 23606 45538 23618 45572
rect 23418 45532 23618 45538
rect 23650 45540 23730 45560
rect 22882 45494 22890 45528
rect 22880 45480 22890 45494
rect 22810 45460 22890 45480
rect 22920 45484 23120 45490
rect 22920 45450 22932 45484
rect 23108 45480 23120 45484
rect 23418 45484 23618 45490
rect 23418 45480 23430 45484
rect 23108 45470 23430 45480
rect 23108 45450 23240 45470
rect 22920 45444 23120 45450
rect 23230 45410 23240 45450
rect 23300 45450 23430 45470
rect 23606 45450 23618 45484
rect 23650 45480 23660 45540
rect 23720 45480 23730 45540
rect 23650 45460 23730 45480
rect 23300 45410 23310 45450
rect 23418 45444 23618 45450
rect 23230 45400 23310 45410
rect 22700 44240 22770 45390
rect 22700 43980 22720 44240
rect 22760 43980 22770 44240
rect 23780 45390 23790 45630
rect 23830 45390 23850 45630
rect 23780 44240 23850 45390
rect 23230 44210 23310 44220
rect 22920 44172 23120 44178
rect 22810 44140 22890 44160
rect 22810 44080 22820 44140
rect 22880 44128 22890 44140
rect 22920 44138 22932 44172
rect 23108 44170 23120 44172
rect 23230 44170 23240 44210
rect 23108 44150 23240 44170
rect 23300 44170 23310 44210
rect 23418 44172 23618 44178
rect 23418 44170 23430 44172
rect 23300 44150 23430 44170
rect 23108 44140 23430 44150
rect 23108 44138 23120 44140
rect 22920 44132 23120 44138
rect 23418 44138 23430 44140
rect 23606 44138 23618 44172
rect 23418 44132 23618 44138
rect 23650 44140 23730 44160
rect 22882 44094 22890 44128
rect 22880 44080 22890 44094
rect 22810 44060 22890 44080
rect 22920 44084 23120 44090
rect 22920 44050 22932 44084
rect 23108 44080 23120 44084
rect 23418 44084 23618 44090
rect 23418 44080 23430 44084
rect 23108 44050 23430 44080
rect 23606 44050 23618 44084
rect 23650 44080 23660 44140
rect 23720 44080 23730 44140
rect 23650 44060 23730 44080
rect 22920 44044 23120 44050
rect 22700 43920 22770 43980
rect 22700 43680 22720 43920
rect 22760 43680 22770 43920
rect 23230 44040 23310 44050
rect 23418 44044 23618 44050
rect 23230 43980 23240 44040
rect 23300 43980 23310 44040
rect 23230 43930 23310 43980
rect 23230 43870 23240 43930
rect 23300 43870 23310 43930
rect 22920 43862 23120 43868
rect 22810 43830 22890 43850
rect 22810 43770 22820 43830
rect 22880 43818 22890 43830
rect 22920 43828 22932 43862
rect 23108 43860 23120 43862
rect 23230 43860 23310 43870
rect 23780 44000 23790 44240
rect 23830 44000 23850 44240
rect 23780 43920 23850 44000
rect 23418 43862 23618 43868
rect 23418 43860 23430 43862
rect 23108 43830 23430 43860
rect 23108 43828 23120 43830
rect 22920 43822 23120 43828
rect 23418 43828 23430 43830
rect 23606 43828 23618 43862
rect 23418 43822 23618 43828
rect 23650 43830 23730 43850
rect 22882 43784 22890 43818
rect 22880 43770 22890 43784
rect 22810 43750 22890 43770
rect 22920 43774 23120 43780
rect 22920 43740 22932 43774
rect 23108 43770 23120 43774
rect 23418 43774 23618 43780
rect 23418 43770 23430 43774
rect 23108 43760 23430 43770
rect 23108 43740 23240 43760
rect 22920 43734 23120 43740
rect 23230 43700 23240 43740
rect 23300 43740 23430 43760
rect 23606 43740 23618 43774
rect 23650 43770 23660 43830
rect 23720 43770 23730 43830
rect 23650 43750 23730 43770
rect 23300 43700 23310 43740
rect 23418 43734 23618 43740
rect 23230 43690 23310 43700
rect 22700 42530 22770 43680
rect 22700 42270 22720 42530
rect 22760 42270 22770 42530
rect 23780 43680 23790 43920
rect 23830 43680 23850 43920
rect 23780 42530 23850 43680
rect 23230 42500 23310 42510
rect 22920 42462 23120 42468
rect 22810 42430 22890 42450
rect 22810 42370 22820 42430
rect 22880 42418 22890 42430
rect 22920 42428 22932 42462
rect 23108 42460 23120 42462
rect 23230 42460 23240 42500
rect 23108 42440 23240 42460
rect 23300 42460 23310 42500
rect 23418 42462 23618 42468
rect 23418 42460 23430 42462
rect 23300 42440 23430 42460
rect 23108 42430 23430 42440
rect 23108 42428 23120 42430
rect 22920 42422 23120 42428
rect 23418 42428 23430 42430
rect 23606 42428 23618 42462
rect 23418 42422 23618 42428
rect 23650 42430 23730 42450
rect 22882 42384 22890 42418
rect 22880 42370 22890 42384
rect 22810 42350 22890 42370
rect 22920 42374 23120 42380
rect 22920 42340 22932 42374
rect 23108 42370 23120 42374
rect 23418 42374 23618 42380
rect 23418 42370 23430 42374
rect 23108 42340 23430 42370
rect 23606 42340 23618 42374
rect 23650 42370 23660 42430
rect 23720 42370 23730 42430
rect 23650 42350 23730 42370
rect 22920 42334 23120 42340
rect 22700 42210 22770 42270
rect 22700 41970 22720 42210
rect 22760 41970 22770 42210
rect 23230 42330 23310 42340
rect 23418 42334 23618 42340
rect 23230 42270 23240 42330
rect 23300 42270 23310 42330
rect 23230 42220 23310 42270
rect 23230 42160 23240 42220
rect 23300 42160 23310 42220
rect 22920 42152 23120 42158
rect 22810 42120 22890 42140
rect 22810 42060 22820 42120
rect 22880 42108 22890 42120
rect 22920 42118 22932 42152
rect 23108 42150 23120 42152
rect 23230 42150 23310 42160
rect 23780 42290 23790 42530
rect 23830 42290 23850 42530
rect 23780 42210 23850 42290
rect 23418 42152 23618 42158
rect 23418 42150 23430 42152
rect 23108 42120 23430 42150
rect 23108 42118 23120 42120
rect 22920 42112 23120 42118
rect 23418 42118 23430 42120
rect 23606 42118 23618 42152
rect 23418 42112 23618 42118
rect 23650 42120 23730 42140
rect 22882 42074 22890 42108
rect 22880 42060 22890 42074
rect 22810 42040 22890 42060
rect 22920 42064 23120 42070
rect 22920 42030 22932 42064
rect 23108 42060 23120 42064
rect 23418 42064 23618 42070
rect 23418 42060 23430 42064
rect 23108 42050 23430 42060
rect 23108 42030 23240 42050
rect 22920 42024 23120 42030
rect 23230 41990 23240 42030
rect 23300 42030 23430 42050
rect 23606 42030 23618 42064
rect 23650 42060 23660 42120
rect 23720 42060 23730 42120
rect 23650 42040 23730 42060
rect 23300 41990 23310 42030
rect 23418 42024 23618 42030
rect 23230 41980 23310 41990
rect 22700 40820 22770 41970
rect 22700 40560 22720 40820
rect 22760 40560 22770 40820
rect 23780 41970 23790 42210
rect 23830 41970 23850 42210
rect 23780 40820 23850 41970
rect 23230 40790 23310 40800
rect 22920 40752 23120 40758
rect 22810 40720 22890 40740
rect 22810 40660 22820 40720
rect 22880 40708 22890 40720
rect 22920 40718 22932 40752
rect 23108 40750 23120 40752
rect 23230 40750 23240 40790
rect 23108 40730 23240 40750
rect 23300 40750 23310 40790
rect 23418 40752 23618 40758
rect 23418 40750 23430 40752
rect 23300 40730 23430 40750
rect 23108 40720 23430 40730
rect 23108 40718 23120 40720
rect 22920 40712 23120 40718
rect 23418 40718 23430 40720
rect 23606 40718 23618 40752
rect 23418 40712 23618 40718
rect 23650 40720 23730 40740
rect 22882 40674 22890 40708
rect 22880 40660 22890 40674
rect 22810 40640 22890 40660
rect 22920 40664 23120 40670
rect 22920 40630 22932 40664
rect 23108 40660 23120 40664
rect 23418 40664 23618 40670
rect 23418 40660 23430 40664
rect 23108 40630 23430 40660
rect 23606 40630 23618 40664
rect 23650 40660 23660 40720
rect 23720 40660 23730 40720
rect 23650 40640 23730 40660
rect 22920 40624 23120 40630
rect 22700 40500 22770 40560
rect 22700 40260 22720 40500
rect 22760 40260 22770 40500
rect 23230 40620 23310 40630
rect 23418 40624 23618 40630
rect 23230 40560 23240 40620
rect 23300 40560 23310 40620
rect 23230 40510 23310 40560
rect 23230 40450 23240 40510
rect 23300 40450 23310 40510
rect 22920 40442 23120 40448
rect 22810 40410 22890 40430
rect 22810 40350 22820 40410
rect 22880 40398 22890 40410
rect 22920 40408 22932 40442
rect 23108 40440 23120 40442
rect 23230 40440 23310 40450
rect 23780 40580 23790 40820
rect 23830 40580 23850 40820
rect 23780 40500 23850 40580
rect 23418 40442 23618 40448
rect 23418 40440 23430 40442
rect 23108 40410 23430 40440
rect 23108 40408 23120 40410
rect 22920 40402 23120 40408
rect 23418 40408 23430 40410
rect 23606 40408 23618 40442
rect 23418 40402 23618 40408
rect 23650 40410 23730 40430
rect 22882 40364 22890 40398
rect 22880 40350 22890 40364
rect 22810 40330 22890 40350
rect 22920 40354 23120 40360
rect 22920 40320 22932 40354
rect 23108 40350 23120 40354
rect 23418 40354 23618 40360
rect 23418 40350 23430 40354
rect 23108 40340 23430 40350
rect 23108 40320 23240 40340
rect 22920 40314 23120 40320
rect 23230 40280 23240 40320
rect 23300 40320 23430 40340
rect 23606 40320 23618 40354
rect 23650 40350 23660 40410
rect 23720 40350 23730 40410
rect 23650 40330 23730 40350
rect 23300 40280 23310 40320
rect 23418 40314 23618 40320
rect 23230 40270 23310 40280
rect 22700 39690 22770 40260
rect 23780 40260 23790 40500
rect 23830 40260 23850 40500
rect 23780 39690 23850 40260
rect 22700 39680 22780 39690
rect 22700 39620 22710 39680
rect 22770 39620 22780 39680
rect 23770 39680 23850 39690
rect 23770 39620 23780 39680
rect 23840 39620 23850 39680
rect 23770 39610 23850 39620
rect 23880 66480 23910 67050
rect 23880 66470 23940 66480
rect 23880 66400 23940 66410
rect 23880 64770 23910 66400
rect 23970 65950 24000 67050
rect 23940 65940 24000 65950
rect 23940 65870 24000 65880
rect 23880 64760 23940 64770
rect 23880 64690 23940 64700
rect 23880 63060 23910 64690
rect 23970 64240 24000 65870
rect 23940 64230 24000 64240
rect 23940 64160 24000 64170
rect 23880 63050 23940 63060
rect 23880 62980 23940 62990
rect 23880 61350 23910 62980
rect 23970 62530 24000 64160
rect 23940 62520 24000 62530
rect 23940 62450 24000 62460
rect 23880 61340 23940 61350
rect 23880 61270 23940 61280
rect 23880 59640 23910 61270
rect 23970 60820 24000 62450
rect 23940 60810 24000 60820
rect 23940 60740 24000 60750
rect 23880 59630 23940 59640
rect 23880 59560 23940 59570
rect 23880 57930 23910 59560
rect 23970 59110 24000 60740
rect 23940 59100 24000 59110
rect 23940 59030 24000 59040
rect 23880 57920 23940 57930
rect 23880 57850 23940 57860
rect 23880 56220 23910 57850
rect 23970 57400 24000 59030
rect 23940 57390 24000 57400
rect 23940 57320 24000 57330
rect 23880 56210 23940 56220
rect 23880 56140 23940 56150
rect 23880 54510 23910 56140
rect 23970 55690 24000 57320
rect 23940 55680 24000 55690
rect 23940 55610 24000 55620
rect 23880 54500 23940 54510
rect 23880 54430 23940 54440
rect 23880 52800 23910 54430
rect 23970 53980 24000 55610
rect 23940 53970 24000 53980
rect 23940 53900 24000 53910
rect 23880 52790 23940 52800
rect 23880 52720 23940 52730
rect 23880 51090 23910 52720
rect 23970 52270 24000 53900
rect 23940 52260 24000 52270
rect 23940 52190 24000 52200
rect 23880 51080 23940 51090
rect 23880 51010 23940 51020
rect 23880 49380 23910 51010
rect 23970 50560 24000 52190
rect 23940 50550 24000 50560
rect 23940 50480 24000 50490
rect 23880 49370 23940 49380
rect 23880 49300 23940 49310
rect 23880 47670 23910 49300
rect 23970 48850 24000 50480
rect 23940 48840 24000 48850
rect 23940 48770 24000 48780
rect 23880 47660 23940 47670
rect 23880 47590 23940 47600
rect 23880 45960 23910 47590
rect 23970 47140 24000 48770
rect 23940 47130 24000 47140
rect 23940 47060 24000 47070
rect 23880 45950 23940 45960
rect 23880 45880 23940 45890
rect 23880 44250 23910 45880
rect 23970 45430 24000 47060
rect 23940 45420 24000 45430
rect 23940 45350 24000 45360
rect 23880 44240 23940 44250
rect 23880 44170 23940 44180
rect 23880 42540 23910 44170
rect 23970 43720 24000 45350
rect 23940 43710 24000 43720
rect 23940 43640 24000 43650
rect 23880 42530 23940 42540
rect 23880 42460 23940 42470
rect 23880 40830 23910 42460
rect 23970 42010 24000 43640
rect 23940 42000 24000 42010
rect 23940 41930 24000 41940
rect 23880 40820 23940 40830
rect 23880 40750 23940 40760
rect 22230 39220 22290 39230
rect 22410 39230 22670 39240
rect 19240 39160 19300 39170
rect 22470 39210 22670 39230
rect 22410 39160 22470 39170
rect 23880 38840 23910 40750
rect 23970 40300 24000 41930
rect 23940 40290 24000 40300
rect 23940 40220 24000 40230
rect 23970 39690 24000 40220
rect 23940 39680 24000 39690
rect 23940 39610 24000 39620
rect 24030 66390 24060 67050
rect 24030 66380 24090 66390
rect 24030 66310 24090 66320
rect 24030 64680 24060 66310
rect 24030 64670 24090 64680
rect 24030 64600 24090 64610
rect 24030 42450 24060 64600
rect 24150 62970 24180 67050
rect 24150 62960 24210 62970
rect 24150 62890 24210 62900
rect 24150 61250 24180 62890
rect 24150 61240 24210 61250
rect 24150 61170 24210 61180
rect 24150 45870 24180 61170
rect 24270 59550 24300 67050
rect 24270 59540 24330 59550
rect 24270 59470 24330 59480
rect 24270 47580 24300 59470
rect 24390 57840 24420 67050
rect 24390 57830 24450 57840
rect 24390 57760 24450 57770
rect 24390 56130 24420 57760
rect 24390 56120 24450 56130
rect 24390 56050 24450 56060
rect 24390 54420 24420 56050
rect 24390 54410 24450 54420
rect 24390 54340 24450 54350
rect 24390 52710 24420 54340
rect 24390 52700 24450 52710
rect 24390 52630 24450 52640
rect 24390 51000 24420 52630
rect 24390 50990 24450 51000
rect 24390 50920 24450 50930
rect 24390 49290 24420 50920
rect 24390 49280 24450 49290
rect 24390 49210 24450 49220
rect 24270 47570 24330 47580
rect 24270 47500 24330 47510
rect 24150 45860 24210 45870
rect 24150 45790 24210 45800
rect 24150 44160 24180 45790
rect 24150 44150 24210 44160
rect 24150 44080 24210 44090
rect 24030 42440 24090 42450
rect 24030 42370 24090 42380
rect 24030 40740 24060 42370
rect 24030 40730 24090 40740
rect 24030 40660 24090 40670
rect 24030 39240 24060 40660
rect 24150 39300 24180 44080
rect 24270 39360 24300 47500
rect 24390 39420 24420 49210
rect 24510 39690 24540 67050
rect 24630 39690 24660 67050
rect 24750 39690 24780 67050
rect 26910 39690 26940 67050
rect 27030 39690 27060 67050
rect 27150 39690 27180 67050
rect 27270 57840 27300 67050
rect 27390 59550 27420 67050
rect 27510 62970 27540 67050
rect 27630 66390 27660 67050
rect 27600 66380 27660 66390
rect 27600 66310 27660 66320
rect 27630 64680 27660 66310
rect 27600 64670 27660 64680
rect 27600 64600 27660 64610
rect 27480 62960 27540 62970
rect 27480 62890 27540 62900
rect 27510 61250 27540 62890
rect 27480 61240 27540 61250
rect 27480 61170 27540 61180
rect 27360 59540 27420 59550
rect 27360 59470 27420 59480
rect 27240 57830 27300 57840
rect 27240 57760 27300 57770
rect 27270 56130 27300 57760
rect 27240 56120 27300 56130
rect 27240 56050 27300 56060
rect 27270 54420 27300 56050
rect 27240 54410 27300 54420
rect 27240 54340 27300 54350
rect 27270 52710 27300 54340
rect 27240 52700 27300 52710
rect 27240 52630 27300 52640
rect 27270 51000 27300 52630
rect 27240 50990 27300 51000
rect 27240 50920 27300 50930
rect 27270 49290 27300 50920
rect 27240 49280 27300 49290
rect 27240 49210 27300 49220
rect 27270 39420 27300 49210
rect 27390 47580 27420 59470
rect 27360 47570 27420 47580
rect 27360 47500 27420 47510
rect 24390 39410 24830 39420
rect 24390 39390 24770 39410
rect 24270 39350 24650 39360
rect 24270 39330 24590 39350
rect 24150 39290 24470 39300
rect 24150 39270 24410 39290
rect 24030 39230 24290 39240
rect 24030 39210 24230 39230
rect 24770 39340 24830 39350
rect 26860 39410 27300 39420
rect 26920 39390 27300 39410
rect 27390 39360 27420 47500
rect 27510 45870 27540 61170
rect 27480 45860 27540 45870
rect 27480 45790 27540 45800
rect 27510 44160 27540 45790
rect 27480 44150 27540 44160
rect 27480 44080 27540 44090
rect 26860 39340 26920 39350
rect 27040 39350 27420 39360
rect 24590 39280 24650 39290
rect 27100 39330 27420 39350
rect 27510 39300 27540 44080
rect 27630 42450 27660 64600
rect 27600 42440 27660 42450
rect 27600 42370 27660 42380
rect 27630 40740 27660 42370
rect 27600 40730 27660 40740
rect 27600 40660 27660 40670
rect 27040 39280 27100 39290
rect 27220 39290 27540 39300
rect 24410 39220 24470 39230
rect 27280 39270 27540 39290
rect 27630 39240 27660 40660
rect 27690 66470 27760 67050
rect 27690 66210 27710 66470
rect 27750 66210 27760 66470
rect 28770 66470 28840 67050
rect 28220 66440 28300 66450
rect 27910 66402 28110 66408
rect 27800 66370 27880 66390
rect 27800 66310 27810 66370
rect 27870 66358 27880 66370
rect 27910 66368 27922 66402
rect 28098 66400 28110 66402
rect 28220 66400 28230 66440
rect 28098 66380 28230 66400
rect 28290 66400 28300 66440
rect 28408 66402 28608 66408
rect 28408 66400 28420 66402
rect 28290 66380 28420 66400
rect 28098 66370 28420 66380
rect 28098 66368 28110 66370
rect 27910 66362 28110 66368
rect 28408 66368 28420 66370
rect 28596 66368 28608 66402
rect 28408 66362 28608 66368
rect 28640 66370 28720 66390
rect 27872 66324 27880 66358
rect 27870 66310 27880 66324
rect 27800 66290 27880 66310
rect 27910 66314 28110 66320
rect 27910 66280 27922 66314
rect 28098 66310 28110 66314
rect 28408 66314 28608 66320
rect 28408 66310 28420 66314
rect 28098 66280 28420 66310
rect 28596 66280 28608 66314
rect 28640 66310 28650 66370
rect 28710 66310 28720 66370
rect 28640 66290 28720 66310
rect 27910 66274 28110 66280
rect 27690 66150 27760 66210
rect 27690 65910 27710 66150
rect 27750 65910 27760 66150
rect 28220 66270 28300 66280
rect 28408 66274 28608 66280
rect 28220 66210 28230 66270
rect 28290 66210 28300 66270
rect 28220 66160 28300 66210
rect 28220 66100 28230 66160
rect 28290 66100 28300 66160
rect 27910 66092 28110 66098
rect 27800 66060 27880 66080
rect 27800 66000 27810 66060
rect 27870 66048 27880 66060
rect 27910 66058 27922 66092
rect 28098 66090 28110 66092
rect 28220 66090 28300 66100
rect 28770 66230 28780 66470
rect 28820 66230 28840 66470
rect 28770 66150 28840 66230
rect 28408 66092 28608 66098
rect 28408 66090 28420 66092
rect 28098 66060 28420 66090
rect 28098 66058 28110 66060
rect 27910 66052 28110 66058
rect 28408 66058 28420 66060
rect 28596 66058 28608 66092
rect 28408 66052 28608 66058
rect 28640 66060 28720 66080
rect 27872 66014 27880 66048
rect 27870 66000 27880 66014
rect 27800 65980 27880 66000
rect 27910 66004 28110 66010
rect 27910 65970 27922 66004
rect 28098 66000 28110 66004
rect 28408 66004 28608 66010
rect 28408 66000 28420 66004
rect 28098 65990 28420 66000
rect 28098 65970 28230 65990
rect 27910 65964 28110 65970
rect 28220 65930 28230 65970
rect 28290 65970 28420 65990
rect 28596 65970 28608 66004
rect 28640 66000 28650 66060
rect 28710 66000 28720 66060
rect 28640 65980 28720 66000
rect 28290 65930 28300 65970
rect 28408 65964 28608 65970
rect 28220 65920 28300 65930
rect 27690 64760 27760 65910
rect 27690 64500 27710 64760
rect 27750 64500 27760 64760
rect 28770 65910 28780 66150
rect 28820 65910 28840 66150
rect 28770 64760 28840 65910
rect 28220 64730 28300 64740
rect 27910 64692 28110 64698
rect 27800 64660 27880 64680
rect 27800 64600 27810 64660
rect 27870 64648 27880 64660
rect 27910 64658 27922 64692
rect 28098 64690 28110 64692
rect 28220 64690 28230 64730
rect 28098 64670 28230 64690
rect 28290 64690 28300 64730
rect 28408 64692 28608 64698
rect 28408 64690 28420 64692
rect 28290 64670 28420 64690
rect 28098 64660 28420 64670
rect 28098 64658 28110 64660
rect 27910 64652 28110 64658
rect 28408 64658 28420 64660
rect 28596 64658 28608 64692
rect 28408 64652 28608 64658
rect 28640 64660 28720 64680
rect 27872 64614 27880 64648
rect 27870 64600 27880 64614
rect 27800 64580 27880 64600
rect 27910 64604 28110 64610
rect 27910 64570 27922 64604
rect 28098 64600 28110 64604
rect 28408 64604 28608 64610
rect 28408 64600 28420 64604
rect 28098 64570 28420 64600
rect 28596 64570 28608 64604
rect 28640 64600 28650 64660
rect 28710 64600 28720 64660
rect 28640 64580 28720 64600
rect 27910 64564 28110 64570
rect 27690 64440 27760 64500
rect 27690 64200 27710 64440
rect 27750 64200 27760 64440
rect 28220 64560 28300 64570
rect 28408 64564 28608 64570
rect 28220 64500 28230 64560
rect 28290 64500 28300 64560
rect 28220 64450 28300 64500
rect 28220 64390 28230 64450
rect 28290 64390 28300 64450
rect 27910 64382 28110 64388
rect 27800 64350 27880 64370
rect 27800 64290 27810 64350
rect 27870 64338 27880 64350
rect 27910 64348 27922 64382
rect 28098 64380 28110 64382
rect 28220 64380 28300 64390
rect 28770 64520 28780 64760
rect 28820 64520 28840 64760
rect 28770 64440 28840 64520
rect 28408 64382 28608 64388
rect 28408 64380 28420 64382
rect 28098 64350 28420 64380
rect 28098 64348 28110 64350
rect 27910 64342 28110 64348
rect 28408 64348 28420 64350
rect 28596 64348 28608 64382
rect 28408 64342 28608 64348
rect 28640 64350 28720 64370
rect 27872 64304 27880 64338
rect 27870 64290 27880 64304
rect 27800 64270 27880 64290
rect 27910 64294 28110 64300
rect 27910 64260 27922 64294
rect 28098 64290 28110 64294
rect 28408 64294 28608 64300
rect 28408 64290 28420 64294
rect 28098 64280 28420 64290
rect 28098 64260 28230 64280
rect 27910 64254 28110 64260
rect 28220 64220 28230 64260
rect 28290 64260 28420 64280
rect 28596 64260 28608 64294
rect 28640 64290 28650 64350
rect 28710 64290 28720 64350
rect 28640 64270 28720 64290
rect 28290 64220 28300 64260
rect 28408 64254 28608 64260
rect 28220 64210 28300 64220
rect 27690 63050 27760 64200
rect 27690 62790 27710 63050
rect 27750 62790 27760 63050
rect 28770 64200 28780 64440
rect 28820 64200 28840 64440
rect 28770 63050 28840 64200
rect 28220 63020 28300 63030
rect 27910 62982 28110 62988
rect 27800 62950 27880 62970
rect 27800 62890 27810 62950
rect 27870 62938 27880 62950
rect 27910 62948 27922 62982
rect 28098 62980 28110 62982
rect 28220 62980 28230 63020
rect 28098 62960 28230 62980
rect 28290 62980 28300 63020
rect 28408 62982 28608 62988
rect 28408 62980 28420 62982
rect 28290 62960 28420 62980
rect 28098 62950 28420 62960
rect 28098 62948 28110 62950
rect 27910 62942 28110 62948
rect 28408 62948 28420 62950
rect 28596 62948 28608 62982
rect 28408 62942 28608 62948
rect 28640 62950 28720 62970
rect 27872 62904 27880 62938
rect 27870 62890 27880 62904
rect 27800 62870 27880 62890
rect 27910 62894 28110 62900
rect 27910 62860 27922 62894
rect 28098 62890 28110 62894
rect 28408 62894 28608 62900
rect 28408 62890 28420 62894
rect 28098 62860 28420 62890
rect 28596 62860 28608 62894
rect 28640 62890 28650 62950
rect 28710 62890 28720 62950
rect 28640 62870 28720 62890
rect 27910 62854 28110 62860
rect 27690 62730 27760 62790
rect 27690 62490 27710 62730
rect 27750 62490 27760 62730
rect 28220 62850 28300 62860
rect 28408 62854 28608 62860
rect 28220 62790 28230 62850
rect 28290 62790 28300 62850
rect 28220 62740 28300 62790
rect 28220 62680 28230 62740
rect 28290 62680 28300 62740
rect 27910 62672 28110 62678
rect 27800 62640 27880 62660
rect 27800 62580 27810 62640
rect 27870 62628 27880 62640
rect 27910 62638 27922 62672
rect 28098 62670 28110 62672
rect 28220 62670 28300 62680
rect 28770 62810 28780 63050
rect 28820 62810 28840 63050
rect 28770 62730 28840 62810
rect 28408 62672 28608 62678
rect 28408 62670 28420 62672
rect 28098 62640 28420 62670
rect 28098 62638 28110 62640
rect 27910 62632 28110 62638
rect 28408 62638 28420 62640
rect 28596 62638 28608 62672
rect 28408 62632 28608 62638
rect 28640 62640 28720 62660
rect 27872 62594 27880 62628
rect 27870 62580 27880 62594
rect 27800 62560 27880 62580
rect 27910 62584 28110 62590
rect 27910 62550 27922 62584
rect 28098 62580 28110 62584
rect 28408 62584 28608 62590
rect 28408 62580 28420 62584
rect 28098 62570 28420 62580
rect 28098 62550 28230 62570
rect 27910 62544 28110 62550
rect 28220 62510 28230 62550
rect 28290 62550 28420 62570
rect 28596 62550 28608 62584
rect 28640 62580 28650 62640
rect 28710 62580 28720 62640
rect 28640 62560 28720 62580
rect 28290 62510 28300 62550
rect 28408 62544 28608 62550
rect 28220 62500 28300 62510
rect 27690 61340 27760 62490
rect 27690 61080 27710 61340
rect 27750 61080 27760 61340
rect 28770 62490 28780 62730
rect 28820 62490 28840 62730
rect 28770 61340 28840 62490
rect 28220 61310 28300 61320
rect 27910 61272 28110 61278
rect 27800 61240 27880 61260
rect 27800 61180 27810 61240
rect 27870 61228 27880 61240
rect 27910 61238 27922 61272
rect 28098 61270 28110 61272
rect 28220 61270 28230 61310
rect 28098 61250 28230 61270
rect 28290 61270 28300 61310
rect 28408 61272 28608 61278
rect 28408 61270 28420 61272
rect 28290 61250 28420 61270
rect 28098 61240 28420 61250
rect 28098 61238 28110 61240
rect 27910 61232 28110 61238
rect 28408 61238 28420 61240
rect 28596 61238 28608 61272
rect 28408 61232 28608 61238
rect 28640 61240 28720 61260
rect 27872 61194 27880 61228
rect 27870 61180 27880 61194
rect 27800 61160 27880 61180
rect 27910 61184 28110 61190
rect 27910 61150 27922 61184
rect 28098 61180 28110 61184
rect 28408 61184 28608 61190
rect 28408 61180 28420 61184
rect 28098 61150 28420 61180
rect 28596 61150 28608 61184
rect 28640 61180 28650 61240
rect 28710 61180 28720 61240
rect 28640 61160 28720 61180
rect 27910 61144 28110 61150
rect 27690 61020 27760 61080
rect 27690 60780 27710 61020
rect 27750 60780 27760 61020
rect 28220 61140 28300 61150
rect 28408 61144 28608 61150
rect 28220 61080 28230 61140
rect 28290 61080 28300 61140
rect 28220 61030 28300 61080
rect 28220 60970 28230 61030
rect 28290 60970 28300 61030
rect 27910 60962 28110 60968
rect 27800 60930 27880 60950
rect 27800 60870 27810 60930
rect 27870 60918 27880 60930
rect 27910 60928 27922 60962
rect 28098 60960 28110 60962
rect 28220 60960 28300 60970
rect 28770 61100 28780 61340
rect 28820 61100 28840 61340
rect 28770 61020 28840 61100
rect 28408 60962 28608 60968
rect 28408 60960 28420 60962
rect 28098 60930 28420 60960
rect 28098 60928 28110 60930
rect 27910 60922 28110 60928
rect 28408 60928 28420 60930
rect 28596 60928 28608 60962
rect 28408 60922 28608 60928
rect 28640 60930 28720 60950
rect 27872 60884 27880 60918
rect 27870 60870 27880 60884
rect 27800 60850 27880 60870
rect 27910 60874 28110 60880
rect 27910 60840 27922 60874
rect 28098 60870 28110 60874
rect 28408 60874 28608 60880
rect 28408 60870 28420 60874
rect 28098 60860 28420 60870
rect 28098 60840 28230 60860
rect 27910 60834 28110 60840
rect 28220 60800 28230 60840
rect 28290 60840 28420 60860
rect 28596 60840 28608 60874
rect 28640 60870 28650 60930
rect 28710 60870 28720 60930
rect 28640 60850 28720 60870
rect 28290 60800 28300 60840
rect 28408 60834 28608 60840
rect 28220 60790 28300 60800
rect 27690 59630 27760 60780
rect 27690 59370 27710 59630
rect 27750 59370 27760 59630
rect 28770 60780 28780 61020
rect 28820 60780 28840 61020
rect 28770 59630 28840 60780
rect 28220 59600 28300 59610
rect 27910 59562 28110 59568
rect 27800 59530 27880 59550
rect 27800 59470 27810 59530
rect 27870 59518 27880 59530
rect 27910 59528 27922 59562
rect 28098 59560 28110 59562
rect 28220 59560 28230 59600
rect 28098 59540 28230 59560
rect 28290 59560 28300 59600
rect 28408 59562 28608 59568
rect 28408 59560 28420 59562
rect 28290 59540 28420 59560
rect 28098 59530 28420 59540
rect 28098 59528 28110 59530
rect 27910 59522 28110 59528
rect 28408 59528 28420 59530
rect 28596 59528 28608 59562
rect 28408 59522 28608 59528
rect 28640 59530 28720 59550
rect 27872 59484 27880 59518
rect 27870 59470 27880 59484
rect 27800 59450 27880 59470
rect 27910 59474 28110 59480
rect 27910 59440 27922 59474
rect 28098 59470 28110 59474
rect 28408 59474 28608 59480
rect 28408 59470 28420 59474
rect 28098 59440 28420 59470
rect 28596 59440 28608 59474
rect 28640 59470 28650 59530
rect 28710 59470 28720 59530
rect 28640 59450 28720 59470
rect 27910 59434 28110 59440
rect 27690 59310 27760 59370
rect 27690 59070 27710 59310
rect 27750 59070 27760 59310
rect 28220 59430 28300 59440
rect 28408 59434 28608 59440
rect 28220 59370 28230 59430
rect 28290 59370 28300 59430
rect 28220 59320 28300 59370
rect 28220 59260 28230 59320
rect 28290 59260 28300 59320
rect 27910 59252 28110 59258
rect 27800 59220 27880 59240
rect 27800 59160 27810 59220
rect 27870 59208 27880 59220
rect 27910 59218 27922 59252
rect 28098 59250 28110 59252
rect 28220 59250 28300 59260
rect 28770 59390 28780 59630
rect 28820 59390 28840 59630
rect 28770 59310 28840 59390
rect 28408 59252 28608 59258
rect 28408 59250 28420 59252
rect 28098 59220 28420 59250
rect 28098 59218 28110 59220
rect 27910 59212 28110 59218
rect 28408 59218 28420 59220
rect 28596 59218 28608 59252
rect 28408 59212 28608 59218
rect 28640 59220 28720 59240
rect 27872 59174 27880 59208
rect 27870 59160 27880 59174
rect 27800 59140 27880 59160
rect 27910 59164 28110 59170
rect 27910 59130 27922 59164
rect 28098 59160 28110 59164
rect 28408 59164 28608 59170
rect 28408 59160 28420 59164
rect 28098 59150 28420 59160
rect 28098 59130 28230 59150
rect 27910 59124 28110 59130
rect 28220 59090 28230 59130
rect 28290 59130 28420 59150
rect 28596 59130 28608 59164
rect 28640 59160 28650 59220
rect 28710 59160 28720 59220
rect 28640 59140 28720 59160
rect 28290 59090 28300 59130
rect 28408 59124 28608 59130
rect 28220 59080 28300 59090
rect 27690 57920 27760 59070
rect 27690 57660 27710 57920
rect 27750 57660 27760 57920
rect 28770 59070 28780 59310
rect 28820 59070 28840 59310
rect 28770 57920 28840 59070
rect 28220 57890 28300 57900
rect 27910 57852 28110 57858
rect 27800 57820 27880 57840
rect 27800 57760 27810 57820
rect 27870 57808 27880 57820
rect 27910 57818 27922 57852
rect 28098 57850 28110 57852
rect 28220 57850 28230 57890
rect 28098 57830 28230 57850
rect 28290 57850 28300 57890
rect 28408 57852 28608 57858
rect 28408 57850 28420 57852
rect 28290 57830 28420 57850
rect 28098 57820 28420 57830
rect 28098 57818 28110 57820
rect 27910 57812 28110 57818
rect 28408 57818 28420 57820
rect 28596 57818 28608 57852
rect 28408 57812 28608 57818
rect 28640 57820 28720 57840
rect 27872 57774 27880 57808
rect 27870 57760 27880 57774
rect 27800 57740 27880 57760
rect 27910 57764 28110 57770
rect 27910 57730 27922 57764
rect 28098 57760 28110 57764
rect 28408 57764 28608 57770
rect 28408 57760 28420 57764
rect 28098 57730 28420 57760
rect 28596 57730 28608 57764
rect 28640 57760 28650 57820
rect 28710 57760 28720 57820
rect 28640 57740 28720 57760
rect 27910 57724 28110 57730
rect 27690 57600 27760 57660
rect 27690 57360 27710 57600
rect 27750 57360 27760 57600
rect 28220 57720 28300 57730
rect 28408 57724 28608 57730
rect 28220 57660 28230 57720
rect 28290 57660 28300 57720
rect 28220 57610 28300 57660
rect 28220 57550 28230 57610
rect 28290 57550 28300 57610
rect 27910 57542 28110 57548
rect 27800 57510 27880 57530
rect 27800 57450 27810 57510
rect 27870 57498 27880 57510
rect 27910 57508 27922 57542
rect 28098 57540 28110 57542
rect 28220 57540 28300 57550
rect 28770 57680 28780 57920
rect 28820 57680 28840 57920
rect 28770 57600 28840 57680
rect 28408 57542 28608 57548
rect 28408 57540 28420 57542
rect 28098 57510 28420 57540
rect 28098 57508 28110 57510
rect 27910 57502 28110 57508
rect 28408 57508 28420 57510
rect 28596 57508 28608 57542
rect 28408 57502 28608 57508
rect 28640 57510 28720 57530
rect 27872 57464 27880 57498
rect 27870 57450 27880 57464
rect 27800 57430 27880 57450
rect 27910 57454 28110 57460
rect 27910 57420 27922 57454
rect 28098 57450 28110 57454
rect 28408 57454 28608 57460
rect 28408 57450 28420 57454
rect 28098 57440 28420 57450
rect 28098 57420 28230 57440
rect 27910 57414 28110 57420
rect 28220 57380 28230 57420
rect 28290 57420 28420 57440
rect 28596 57420 28608 57454
rect 28640 57450 28650 57510
rect 28710 57450 28720 57510
rect 28640 57430 28720 57450
rect 28290 57380 28300 57420
rect 28408 57414 28608 57420
rect 28220 57370 28300 57380
rect 27690 56210 27760 57360
rect 27690 55950 27710 56210
rect 27750 55950 27760 56210
rect 28770 57360 28780 57600
rect 28820 57360 28840 57600
rect 28770 56210 28840 57360
rect 28220 56180 28300 56190
rect 27910 56142 28110 56148
rect 27800 56110 27880 56130
rect 27800 56050 27810 56110
rect 27870 56098 27880 56110
rect 27910 56108 27922 56142
rect 28098 56140 28110 56142
rect 28220 56140 28230 56180
rect 28098 56120 28230 56140
rect 28290 56140 28300 56180
rect 28408 56142 28608 56148
rect 28408 56140 28420 56142
rect 28290 56120 28420 56140
rect 28098 56110 28420 56120
rect 28098 56108 28110 56110
rect 27910 56102 28110 56108
rect 28408 56108 28420 56110
rect 28596 56108 28608 56142
rect 28408 56102 28608 56108
rect 28640 56110 28720 56130
rect 27872 56064 27880 56098
rect 27870 56050 27880 56064
rect 27800 56030 27880 56050
rect 27910 56054 28110 56060
rect 27910 56020 27922 56054
rect 28098 56050 28110 56054
rect 28408 56054 28608 56060
rect 28408 56050 28420 56054
rect 28098 56020 28420 56050
rect 28596 56020 28608 56054
rect 28640 56050 28650 56110
rect 28710 56050 28720 56110
rect 28640 56030 28720 56050
rect 27910 56014 28110 56020
rect 27690 55890 27760 55950
rect 27690 55650 27710 55890
rect 27750 55650 27760 55890
rect 28220 56010 28300 56020
rect 28408 56014 28608 56020
rect 28220 55950 28230 56010
rect 28290 55950 28300 56010
rect 28220 55900 28300 55950
rect 28220 55840 28230 55900
rect 28290 55840 28300 55900
rect 27910 55832 28110 55838
rect 27800 55800 27880 55820
rect 27800 55740 27810 55800
rect 27870 55788 27880 55800
rect 27910 55798 27922 55832
rect 28098 55830 28110 55832
rect 28220 55830 28300 55840
rect 28770 55970 28780 56210
rect 28820 55970 28840 56210
rect 28770 55890 28840 55970
rect 28408 55832 28608 55838
rect 28408 55830 28420 55832
rect 28098 55800 28420 55830
rect 28098 55798 28110 55800
rect 27910 55792 28110 55798
rect 28408 55798 28420 55800
rect 28596 55798 28608 55832
rect 28408 55792 28608 55798
rect 28640 55800 28720 55820
rect 27872 55754 27880 55788
rect 27870 55740 27880 55754
rect 27800 55720 27880 55740
rect 27910 55744 28110 55750
rect 27910 55710 27922 55744
rect 28098 55740 28110 55744
rect 28408 55744 28608 55750
rect 28408 55740 28420 55744
rect 28098 55730 28420 55740
rect 28098 55710 28230 55730
rect 27910 55704 28110 55710
rect 28220 55670 28230 55710
rect 28290 55710 28420 55730
rect 28596 55710 28608 55744
rect 28640 55740 28650 55800
rect 28710 55740 28720 55800
rect 28640 55720 28720 55740
rect 28290 55670 28300 55710
rect 28408 55704 28608 55710
rect 28220 55660 28300 55670
rect 27690 54500 27760 55650
rect 27690 54240 27710 54500
rect 27750 54240 27760 54500
rect 28770 55650 28780 55890
rect 28820 55650 28840 55890
rect 28770 54500 28840 55650
rect 28220 54470 28300 54480
rect 27910 54432 28110 54438
rect 27800 54400 27880 54420
rect 27800 54340 27810 54400
rect 27870 54388 27880 54400
rect 27910 54398 27922 54432
rect 28098 54430 28110 54432
rect 28220 54430 28230 54470
rect 28098 54410 28230 54430
rect 28290 54430 28300 54470
rect 28408 54432 28608 54438
rect 28408 54430 28420 54432
rect 28290 54410 28420 54430
rect 28098 54400 28420 54410
rect 28098 54398 28110 54400
rect 27910 54392 28110 54398
rect 28408 54398 28420 54400
rect 28596 54398 28608 54432
rect 28408 54392 28608 54398
rect 28640 54400 28720 54420
rect 27872 54354 27880 54388
rect 27870 54340 27880 54354
rect 27800 54320 27880 54340
rect 27910 54344 28110 54350
rect 27910 54310 27922 54344
rect 28098 54340 28110 54344
rect 28408 54344 28608 54350
rect 28408 54340 28420 54344
rect 28098 54310 28420 54340
rect 28596 54310 28608 54344
rect 28640 54340 28650 54400
rect 28710 54340 28720 54400
rect 28640 54320 28720 54340
rect 27910 54304 28110 54310
rect 27690 54180 27760 54240
rect 27690 53940 27710 54180
rect 27750 53940 27760 54180
rect 28220 54300 28300 54310
rect 28408 54304 28608 54310
rect 28220 54240 28230 54300
rect 28290 54240 28300 54300
rect 28220 54190 28300 54240
rect 28220 54130 28230 54190
rect 28290 54130 28300 54190
rect 27910 54122 28110 54128
rect 27800 54090 27880 54110
rect 27800 54030 27810 54090
rect 27870 54078 27880 54090
rect 27910 54088 27922 54122
rect 28098 54120 28110 54122
rect 28220 54120 28300 54130
rect 28770 54260 28780 54500
rect 28820 54260 28840 54500
rect 28770 54180 28840 54260
rect 28408 54122 28608 54128
rect 28408 54120 28420 54122
rect 28098 54090 28420 54120
rect 28098 54088 28110 54090
rect 27910 54082 28110 54088
rect 28408 54088 28420 54090
rect 28596 54088 28608 54122
rect 28408 54082 28608 54088
rect 28640 54090 28720 54110
rect 27872 54044 27880 54078
rect 27870 54030 27880 54044
rect 27800 54010 27880 54030
rect 27910 54034 28110 54040
rect 27910 54000 27922 54034
rect 28098 54030 28110 54034
rect 28408 54034 28608 54040
rect 28408 54030 28420 54034
rect 28098 54020 28420 54030
rect 28098 54000 28230 54020
rect 27910 53994 28110 54000
rect 28220 53960 28230 54000
rect 28290 54000 28420 54020
rect 28596 54000 28608 54034
rect 28640 54030 28650 54090
rect 28710 54030 28720 54090
rect 28640 54010 28720 54030
rect 28290 53960 28300 54000
rect 28408 53994 28608 54000
rect 28220 53950 28300 53960
rect 27690 52790 27760 53940
rect 27690 52530 27710 52790
rect 27750 52530 27760 52790
rect 28770 53940 28780 54180
rect 28820 53940 28840 54180
rect 28770 52790 28840 53940
rect 28220 52760 28300 52770
rect 27910 52722 28110 52728
rect 27800 52690 27880 52710
rect 27800 52630 27810 52690
rect 27870 52678 27880 52690
rect 27910 52688 27922 52722
rect 28098 52720 28110 52722
rect 28220 52720 28230 52760
rect 28098 52700 28230 52720
rect 28290 52720 28300 52760
rect 28408 52722 28608 52728
rect 28408 52720 28420 52722
rect 28290 52700 28420 52720
rect 28098 52690 28420 52700
rect 28098 52688 28110 52690
rect 27910 52682 28110 52688
rect 28408 52688 28420 52690
rect 28596 52688 28608 52722
rect 28408 52682 28608 52688
rect 28640 52690 28720 52710
rect 27872 52644 27880 52678
rect 27870 52630 27880 52644
rect 27800 52610 27880 52630
rect 27910 52634 28110 52640
rect 27910 52600 27922 52634
rect 28098 52630 28110 52634
rect 28408 52634 28608 52640
rect 28408 52630 28420 52634
rect 28098 52600 28420 52630
rect 28596 52600 28608 52634
rect 28640 52630 28650 52690
rect 28710 52630 28720 52690
rect 28640 52610 28720 52630
rect 27910 52594 28110 52600
rect 27690 52470 27760 52530
rect 27690 52230 27710 52470
rect 27750 52230 27760 52470
rect 28220 52590 28300 52600
rect 28408 52594 28608 52600
rect 28220 52530 28230 52590
rect 28290 52530 28300 52590
rect 28220 52480 28300 52530
rect 28220 52420 28230 52480
rect 28290 52420 28300 52480
rect 27910 52412 28110 52418
rect 27800 52380 27880 52400
rect 27800 52320 27810 52380
rect 27870 52368 27880 52380
rect 27910 52378 27922 52412
rect 28098 52410 28110 52412
rect 28220 52410 28300 52420
rect 28770 52550 28780 52790
rect 28820 52550 28840 52790
rect 28770 52470 28840 52550
rect 28408 52412 28608 52418
rect 28408 52410 28420 52412
rect 28098 52380 28420 52410
rect 28098 52378 28110 52380
rect 27910 52372 28110 52378
rect 28408 52378 28420 52380
rect 28596 52378 28608 52412
rect 28408 52372 28608 52378
rect 28640 52380 28720 52400
rect 27872 52334 27880 52368
rect 27870 52320 27880 52334
rect 27800 52300 27880 52320
rect 27910 52324 28110 52330
rect 27910 52290 27922 52324
rect 28098 52320 28110 52324
rect 28408 52324 28608 52330
rect 28408 52320 28420 52324
rect 28098 52310 28420 52320
rect 28098 52290 28230 52310
rect 27910 52284 28110 52290
rect 28220 52250 28230 52290
rect 28290 52290 28420 52310
rect 28596 52290 28608 52324
rect 28640 52320 28650 52380
rect 28710 52320 28720 52380
rect 28640 52300 28720 52320
rect 28290 52250 28300 52290
rect 28408 52284 28608 52290
rect 28220 52240 28300 52250
rect 27690 51080 27760 52230
rect 27690 50820 27710 51080
rect 27750 50820 27760 51080
rect 28770 52230 28780 52470
rect 28820 52230 28840 52470
rect 28770 51080 28840 52230
rect 28220 51050 28300 51060
rect 27910 51012 28110 51018
rect 27800 50980 27880 51000
rect 27800 50920 27810 50980
rect 27870 50968 27880 50980
rect 27910 50978 27922 51012
rect 28098 51010 28110 51012
rect 28220 51010 28230 51050
rect 28098 50990 28230 51010
rect 28290 51010 28300 51050
rect 28408 51012 28608 51018
rect 28408 51010 28420 51012
rect 28290 50990 28420 51010
rect 28098 50980 28420 50990
rect 28098 50978 28110 50980
rect 27910 50972 28110 50978
rect 28408 50978 28420 50980
rect 28596 50978 28608 51012
rect 28408 50972 28608 50978
rect 28640 50980 28720 51000
rect 27872 50934 27880 50968
rect 27870 50920 27880 50934
rect 27800 50900 27880 50920
rect 27910 50924 28110 50930
rect 27910 50890 27922 50924
rect 28098 50920 28110 50924
rect 28408 50924 28608 50930
rect 28408 50920 28420 50924
rect 28098 50890 28420 50920
rect 28596 50890 28608 50924
rect 28640 50920 28650 50980
rect 28710 50920 28720 50980
rect 28640 50900 28720 50920
rect 27910 50884 28110 50890
rect 27690 50760 27760 50820
rect 27690 50520 27710 50760
rect 27750 50520 27760 50760
rect 28220 50880 28300 50890
rect 28408 50884 28608 50890
rect 28220 50820 28230 50880
rect 28290 50820 28300 50880
rect 28220 50770 28300 50820
rect 28220 50710 28230 50770
rect 28290 50710 28300 50770
rect 27910 50702 28110 50708
rect 27800 50670 27880 50690
rect 27800 50610 27810 50670
rect 27870 50658 27880 50670
rect 27910 50668 27922 50702
rect 28098 50700 28110 50702
rect 28220 50700 28300 50710
rect 28770 50840 28780 51080
rect 28820 50840 28840 51080
rect 28770 50760 28840 50840
rect 28408 50702 28608 50708
rect 28408 50700 28420 50702
rect 28098 50670 28420 50700
rect 28098 50668 28110 50670
rect 27910 50662 28110 50668
rect 28408 50668 28420 50670
rect 28596 50668 28608 50702
rect 28408 50662 28608 50668
rect 28640 50670 28720 50690
rect 27872 50624 27880 50658
rect 27870 50610 27880 50624
rect 27800 50590 27880 50610
rect 27910 50614 28110 50620
rect 27910 50580 27922 50614
rect 28098 50610 28110 50614
rect 28408 50614 28608 50620
rect 28408 50610 28420 50614
rect 28098 50600 28420 50610
rect 28098 50580 28230 50600
rect 27910 50574 28110 50580
rect 28220 50540 28230 50580
rect 28290 50580 28420 50600
rect 28596 50580 28608 50614
rect 28640 50610 28650 50670
rect 28710 50610 28720 50670
rect 28640 50590 28720 50610
rect 28290 50540 28300 50580
rect 28408 50574 28608 50580
rect 28220 50530 28300 50540
rect 27690 49370 27760 50520
rect 27690 49110 27710 49370
rect 27750 49110 27760 49370
rect 28770 50520 28780 50760
rect 28820 50520 28840 50760
rect 28770 49370 28840 50520
rect 28220 49340 28300 49350
rect 27910 49302 28110 49308
rect 27800 49270 27880 49290
rect 27800 49210 27810 49270
rect 27870 49258 27880 49270
rect 27910 49268 27922 49302
rect 28098 49300 28110 49302
rect 28220 49300 28230 49340
rect 28098 49280 28230 49300
rect 28290 49300 28300 49340
rect 28408 49302 28608 49308
rect 28408 49300 28420 49302
rect 28290 49280 28420 49300
rect 28098 49270 28420 49280
rect 28098 49268 28110 49270
rect 27910 49262 28110 49268
rect 28408 49268 28420 49270
rect 28596 49268 28608 49302
rect 28408 49262 28608 49268
rect 28640 49270 28720 49290
rect 27872 49224 27880 49258
rect 27870 49210 27880 49224
rect 27800 49190 27880 49210
rect 27910 49214 28110 49220
rect 27910 49180 27922 49214
rect 28098 49210 28110 49214
rect 28408 49214 28608 49220
rect 28408 49210 28420 49214
rect 28098 49180 28420 49210
rect 28596 49180 28608 49214
rect 28640 49210 28650 49270
rect 28710 49210 28720 49270
rect 28640 49190 28720 49210
rect 27910 49174 28110 49180
rect 27690 49050 27760 49110
rect 27690 48810 27710 49050
rect 27750 48810 27760 49050
rect 28220 49170 28300 49180
rect 28408 49174 28608 49180
rect 28220 49110 28230 49170
rect 28290 49110 28300 49170
rect 28220 49060 28300 49110
rect 28220 49000 28230 49060
rect 28290 49000 28300 49060
rect 27910 48992 28110 48998
rect 27800 48960 27880 48980
rect 27800 48900 27810 48960
rect 27870 48948 27880 48960
rect 27910 48958 27922 48992
rect 28098 48990 28110 48992
rect 28220 48990 28300 49000
rect 28770 49130 28780 49370
rect 28820 49130 28840 49370
rect 28770 49050 28840 49130
rect 28408 48992 28608 48998
rect 28408 48990 28420 48992
rect 28098 48960 28420 48990
rect 28098 48958 28110 48960
rect 27910 48952 28110 48958
rect 28408 48958 28420 48960
rect 28596 48958 28608 48992
rect 28408 48952 28608 48958
rect 28640 48960 28720 48980
rect 27872 48914 27880 48948
rect 27870 48900 27880 48914
rect 27800 48880 27880 48900
rect 27910 48904 28110 48910
rect 27910 48870 27922 48904
rect 28098 48900 28110 48904
rect 28408 48904 28608 48910
rect 28408 48900 28420 48904
rect 28098 48890 28420 48900
rect 28098 48870 28230 48890
rect 27910 48864 28110 48870
rect 28220 48830 28230 48870
rect 28290 48870 28420 48890
rect 28596 48870 28608 48904
rect 28640 48900 28650 48960
rect 28710 48900 28720 48960
rect 28640 48880 28720 48900
rect 28290 48830 28300 48870
rect 28408 48864 28608 48870
rect 28220 48820 28300 48830
rect 27690 47660 27760 48810
rect 27690 47400 27710 47660
rect 27750 47400 27760 47660
rect 28770 48810 28780 49050
rect 28820 48810 28840 49050
rect 28770 47660 28840 48810
rect 28220 47630 28300 47640
rect 27910 47592 28110 47598
rect 27800 47560 27880 47580
rect 27800 47500 27810 47560
rect 27870 47548 27880 47560
rect 27910 47558 27922 47592
rect 28098 47590 28110 47592
rect 28220 47590 28230 47630
rect 28098 47570 28230 47590
rect 28290 47590 28300 47630
rect 28408 47592 28608 47598
rect 28408 47590 28420 47592
rect 28290 47570 28420 47590
rect 28098 47560 28420 47570
rect 28098 47558 28110 47560
rect 27910 47552 28110 47558
rect 28408 47558 28420 47560
rect 28596 47558 28608 47592
rect 28408 47552 28608 47558
rect 28640 47560 28720 47580
rect 27872 47514 27880 47548
rect 27870 47500 27880 47514
rect 27800 47480 27880 47500
rect 27910 47504 28110 47510
rect 27910 47470 27922 47504
rect 28098 47500 28110 47504
rect 28408 47504 28608 47510
rect 28408 47500 28420 47504
rect 28098 47470 28420 47500
rect 28596 47470 28608 47504
rect 28640 47500 28650 47560
rect 28710 47500 28720 47560
rect 28640 47480 28720 47500
rect 27910 47464 28110 47470
rect 27690 47340 27760 47400
rect 27690 47100 27710 47340
rect 27750 47100 27760 47340
rect 28220 47460 28300 47470
rect 28408 47464 28608 47470
rect 28220 47400 28230 47460
rect 28290 47400 28300 47460
rect 28220 47350 28300 47400
rect 28220 47290 28230 47350
rect 28290 47290 28300 47350
rect 27910 47282 28110 47288
rect 27800 47250 27880 47270
rect 27800 47190 27810 47250
rect 27870 47238 27880 47250
rect 27910 47248 27922 47282
rect 28098 47280 28110 47282
rect 28220 47280 28300 47290
rect 28770 47420 28780 47660
rect 28820 47420 28840 47660
rect 28770 47340 28840 47420
rect 28408 47282 28608 47288
rect 28408 47280 28420 47282
rect 28098 47250 28420 47280
rect 28098 47248 28110 47250
rect 27910 47242 28110 47248
rect 28408 47248 28420 47250
rect 28596 47248 28608 47282
rect 28408 47242 28608 47248
rect 28640 47250 28720 47270
rect 27872 47204 27880 47238
rect 27870 47190 27880 47204
rect 27800 47170 27880 47190
rect 27910 47194 28110 47200
rect 27910 47160 27922 47194
rect 28098 47190 28110 47194
rect 28408 47194 28608 47200
rect 28408 47190 28420 47194
rect 28098 47180 28420 47190
rect 28098 47160 28230 47180
rect 27910 47154 28110 47160
rect 28220 47120 28230 47160
rect 28290 47160 28420 47180
rect 28596 47160 28608 47194
rect 28640 47190 28650 47250
rect 28710 47190 28720 47250
rect 28640 47170 28720 47190
rect 28290 47120 28300 47160
rect 28408 47154 28608 47160
rect 28220 47110 28300 47120
rect 27690 45950 27760 47100
rect 27690 45690 27710 45950
rect 27750 45690 27760 45950
rect 28770 47100 28780 47340
rect 28820 47100 28840 47340
rect 28770 45950 28840 47100
rect 28220 45920 28300 45930
rect 27910 45882 28110 45888
rect 27800 45850 27880 45870
rect 27800 45790 27810 45850
rect 27870 45838 27880 45850
rect 27910 45848 27922 45882
rect 28098 45880 28110 45882
rect 28220 45880 28230 45920
rect 28098 45860 28230 45880
rect 28290 45880 28300 45920
rect 28408 45882 28608 45888
rect 28408 45880 28420 45882
rect 28290 45860 28420 45880
rect 28098 45850 28420 45860
rect 28098 45848 28110 45850
rect 27910 45842 28110 45848
rect 28408 45848 28420 45850
rect 28596 45848 28608 45882
rect 28408 45842 28608 45848
rect 28640 45850 28720 45870
rect 27872 45804 27880 45838
rect 27870 45790 27880 45804
rect 27800 45770 27880 45790
rect 27910 45794 28110 45800
rect 27910 45760 27922 45794
rect 28098 45790 28110 45794
rect 28408 45794 28608 45800
rect 28408 45790 28420 45794
rect 28098 45760 28420 45790
rect 28596 45760 28608 45794
rect 28640 45790 28650 45850
rect 28710 45790 28720 45850
rect 28640 45770 28720 45790
rect 27910 45754 28110 45760
rect 27690 45630 27760 45690
rect 27690 45390 27710 45630
rect 27750 45390 27760 45630
rect 28220 45750 28300 45760
rect 28408 45754 28608 45760
rect 28220 45690 28230 45750
rect 28290 45690 28300 45750
rect 28220 45640 28300 45690
rect 28220 45580 28230 45640
rect 28290 45580 28300 45640
rect 27910 45572 28110 45578
rect 27800 45540 27880 45560
rect 27800 45480 27810 45540
rect 27870 45528 27880 45540
rect 27910 45538 27922 45572
rect 28098 45570 28110 45572
rect 28220 45570 28300 45580
rect 28770 45710 28780 45950
rect 28820 45710 28840 45950
rect 28770 45630 28840 45710
rect 28408 45572 28608 45578
rect 28408 45570 28420 45572
rect 28098 45540 28420 45570
rect 28098 45538 28110 45540
rect 27910 45532 28110 45538
rect 28408 45538 28420 45540
rect 28596 45538 28608 45572
rect 28408 45532 28608 45538
rect 28640 45540 28720 45560
rect 27872 45494 27880 45528
rect 27870 45480 27880 45494
rect 27800 45460 27880 45480
rect 27910 45484 28110 45490
rect 27910 45450 27922 45484
rect 28098 45480 28110 45484
rect 28408 45484 28608 45490
rect 28408 45480 28420 45484
rect 28098 45470 28420 45480
rect 28098 45450 28230 45470
rect 27910 45444 28110 45450
rect 28220 45410 28230 45450
rect 28290 45450 28420 45470
rect 28596 45450 28608 45484
rect 28640 45480 28650 45540
rect 28710 45480 28720 45540
rect 28640 45460 28720 45480
rect 28290 45410 28300 45450
rect 28408 45444 28608 45450
rect 28220 45400 28300 45410
rect 27690 44240 27760 45390
rect 27690 43980 27710 44240
rect 27750 43980 27760 44240
rect 28770 45390 28780 45630
rect 28820 45390 28840 45630
rect 28770 44240 28840 45390
rect 28220 44210 28300 44220
rect 27910 44172 28110 44178
rect 27800 44140 27880 44160
rect 27800 44080 27810 44140
rect 27870 44128 27880 44140
rect 27910 44138 27922 44172
rect 28098 44170 28110 44172
rect 28220 44170 28230 44210
rect 28098 44150 28230 44170
rect 28290 44170 28300 44210
rect 28408 44172 28608 44178
rect 28408 44170 28420 44172
rect 28290 44150 28420 44170
rect 28098 44140 28420 44150
rect 28098 44138 28110 44140
rect 27910 44132 28110 44138
rect 28408 44138 28420 44140
rect 28596 44138 28608 44172
rect 28408 44132 28608 44138
rect 28640 44140 28720 44160
rect 27872 44094 27880 44128
rect 27870 44080 27880 44094
rect 27800 44060 27880 44080
rect 27910 44084 28110 44090
rect 27910 44050 27922 44084
rect 28098 44080 28110 44084
rect 28408 44084 28608 44090
rect 28408 44080 28420 44084
rect 28098 44050 28420 44080
rect 28596 44050 28608 44084
rect 28640 44080 28650 44140
rect 28710 44080 28720 44140
rect 28640 44060 28720 44080
rect 27910 44044 28110 44050
rect 27690 43920 27760 43980
rect 27690 43680 27710 43920
rect 27750 43680 27760 43920
rect 28220 44040 28300 44050
rect 28408 44044 28608 44050
rect 28220 43980 28230 44040
rect 28290 43980 28300 44040
rect 28220 43930 28300 43980
rect 28220 43870 28230 43930
rect 28290 43870 28300 43930
rect 27910 43862 28110 43868
rect 27800 43830 27880 43850
rect 27800 43770 27810 43830
rect 27870 43818 27880 43830
rect 27910 43828 27922 43862
rect 28098 43860 28110 43862
rect 28220 43860 28300 43870
rect 28770 44000 28780 44240
rect 28820 44000 28840 44240
rect 28770 43920 28840 44000
rect 28408 43862 28608 43868
rect 28408 43860 28420 43862
rect 28098 43830 28420 43860
rect 28098 43828 28110 43830
rect 27910 43822 28110 43828
rect 28408 43828 28420 43830
rect 28596 43828 28608 43862
rect 28408 43822 28608 43828
rect 28640 43830 28720 43850
rect 27872 43784 27880 43818
rect 27870 43770 27880 43784
rect 27800 43750 27880 43770
rect 27910 43774 28110 43780
rect 27910 43740 27922 43774
rect 28098 43770 28110 43774
rect 28408 43774 28608 43780
rect 28408 43770 28420 43774
rect 28098 43760 28420 43770
rect 28098 43740 28230 43760
rect 27910 43734 28110 43740
rect 28220 43700 28230 43740
rect 28290 43740 28420 43760
rect 28596 43740 28608 43774
rect 28640 43770 28650 43830
rect 28710 43770 28720 43830
rect 28640 43750 28720 43770
rect 28290 43700 28300 43740
rect 28408 43734 28608 43740
rect 28220 43690 28300 43700
rect 27690 42530 27760 43680
rect 27690 42270 27710 42530
rect 27750 42270 27760 42530
rect 28770 43680 28780 43920
rect 28820 43680 28840 43920
rect 28770 42530 28840 43680
rect 28220 42500 28300 42510
rect 27910 42462 28110 42468
rect 27800 42430 27880 42450
rect 27800 42370 27810 42430
rect 27870 42418 27880 42430
rect 27910 42428 27922 42462
rect 28098 42460 28110 42462
rect 28220 42460 28230 42500
rect 28098 42440 28230 42460
rect 28290 42460 28300 42500
rect 28408 42462 28608 42468
rect 28408 42460 28420 42462
rect 28290 42440 28420 42460
rect 28098 42430 28420 42440
rect 28098 42428 28110 42430
rect 27910 42422 28110 42428
rect 28408 42428 28420 42430
rect 28596 42428 28608 42462
rect 28408 42422 28608 42428
rect 28640 42430 28720 42450
rect 27872 42384 27880 42418
rect 27870 42370 27880 42384
rect 27800 42350 27880 42370
rect 27910 42374 28110 42380
rect 27910 42340 27922 42374
rect 28098 42370 28110 42374
rect 28408 42374 28608 42380
rect 28408 42370 28420 42374
rect 28098 42340 28420 42370
rect 28596 42340 28608 42374
rect 28640 42370 28650 42430
rect 28710 42370 28720 42430
rect 28640 42350 28720 42370
rect 27910 42334 28110 42340
rect 27690 42210 27760 42270
rect 27690 41970 27710 42210
rect 27750 41970 27760 42210
rect 28220 42330 28300 42340
rect 28408 42334 28608 42340
rect 28220 42270 28230 42330
rect 28290 42270 28300 42330
rect 28220 42220 28300 42270
rect 28220 42160 28230 42220
rect 28290 42160 28300 42220
rect 27910 42152 28110 42158
rect 27800 42120 27880 42140
rect 27800 42060 27810 42120
rect 27870 42108 27880 42120
rect 27910 42118 27922 42152
rect 28098 42150 28110 42152
rect 28220 42150 28300 42160
rect 28770 42290 28780 42530
rect 28820 42290 28840 42530
rect 28770 42210 28840 42290
rect 28408 42152 28608 42158
rect 28408 42150 28420 42152
rect 28098 42120 28420 42150
rect 28098 42118 28110 42120
rect 27910 42112 28110 42118
rect 28408 42118 28420 42120
rect 28596 42118 28608 42152
rect 28408 42112 28608 42118
rect 28640 42120 28720 42140
rect 27872 42074 27880 42108
rect 27870 42060 27880 42074
rect 27800 42040 27880 42060
rect 27910 42064 28110 42070
rect 27910 42030 27922 42064
rect 28098 42060 28110 42064
rect 28408 42064 28608 42070
rect 28408 42060 28420 42064
rect 28098 42050 28420 42060
rect 28098 42030 28230 42050
rect 27910 42024 28110 42030
rect 28220 41990 28230 42030
rect 28290 42030 28420 42050
rect 28596 42030 28608 42064
rect 28640 42060 28650 42120
rect 28710 42060 28720 42120
rect 28640 42040 28720 42060
rect 28290 41990 28300 42030
rect 28408 42024 28608 42030
rect 28220 41980 28300 41990
rect 27690 40820 27760 41970
rect 27690 40560 27710 40820
rect 27750 40560 27760 40820
rect 28770 41970 28780 42210
rect 28820 41970 28840 42210
rect 28770 40820 28840 41970
rect 28220 40790 28300 40800
rect 27910 40752 28110 40758
rect 27800 40720 27880 40740
rect 27800 40660 27810 40720
rect 27870 40708 27880 40720
rect 27910 40718 27922 40752
rect 28098 40750 28110 40752
rect 28220 40750 28230 40790
rect 28098 40730 28230 40750
rect 28290 40750 28300 40790
rect 28408 40752 28608 40758
rect 28408 40750 28420 40752
rect 28290 40730 28420 40750
rect 28098 40720 28420 40730
rect 28098 40718 28110 40720
rect 27910 40712 28110 40718
rect 28408 40718 28420 40720
rect 28596 40718 28608 40752
rect 28408 40712 28608 40718
rect 28640 40720 28720 40740
rect 27872 40674 27880 40708
rect 27870 40660 27880 40674
rect 27800 40640 27880 40660
rect 27910 40664 28110 40670
rect 27910 40630 27922 40664
rect 28098 40660 28110 40664
rect 28408 40664 28608 40670
rect 28408 40660 28420 40664
rect 28098 40630 28420 40660
rect 28596 40630 28608 40664
rect 28640 40660 28650 40720
rect 28710 40660 28720 40720
rect 28640 40640 28720 40660
rect 27910 40624 28110 40630
rect 27690 40500 27760 40560
rect 27690 40260 27710 40500
rect 27750 40260 27760 40500
rect 28220 40620 28300 40630
rect 28408 40624 28608 40630
rect 28220 40560 28230 40620
rect 28290 40560 28300 40620
rect 28220 40510 28300 40560
rect 28220 40450 28230 40510
rect 28290 40450 28300 40510
rect 27910 40442 28110 40448
rect 27800 40410 27880 40430
rect 27800 40350 27810 40410
rect 27870 40398 27880 40410
rect 27910 40408 27922 40442
rect 28098 40440 28110 40442
rect 28220 40440 28300 40450
rect 28770 40580 28780 40820
rect 28820 40580 28840 40820
rect 28770 40500 28840 40580
rect 28408 40442 28608 40448
rect 28408 40440 28420 40442
rect 28098 40410 28420 40440
rect 28098 40408 28110 40410
rect 27910 40402 28110 40408
rect 28408 40408 28420 40410
rect 28596 40408 28608 40442
rect 28408 40402 28608 40408
rect 28640 40410 28720 40430
rect 27872 40364 27880 40398
rect 27870 40350 27880 40364
rect 27800 40330 27880 40350
rect 27910 40354 28110 40360
rect 27910 40320 27922 40354
rect 28098 40350 28110 40354
rect 28408 40354 28608 40360
rect 28408 40350 28420 40354
rect 28098 40340 28420 40350
rect 28098 40320 28230 40340
rect 27910 40314 28110 40320
rect 28220 40280 28230 40320
rect 28290 40320 28420 40340
rect 28596 40320 28608 40354
rect 28640 40350 28650 40410
rect 28710 40350 28720 40410
rect 28640 40330 28720 40350
rect 28290 40280 28300 40320
rect 28408 40314 28608 40320
rect 28220 40270 28300 40280
rect 27690 39690 27760 40260
rect 28770 40260 28780 40500
rect 28820 40260 28840 40500
rect 28770 39690 28840 40260
rect 27690 39680 27770 39690
rect 27690 39620 27700 39680
rect 27760 39620 27770 39680
rect 28760 39680 28840 39690
rect 28760 39620 28770 39680
rect 28830 39620 28840 39680
rect 28760 39610 28840 39620
rect 28870 66480 28900 67050
rect 28870 66470 28930 66480
rect 28870 66400 28930 66410
rect 28870 64770 28900 66400
rect 28960 65950 28990 67050
rect 28930 65940 28990 65950
rect 28930 65870 28990 65880
rect 28870 64760 28930 64770
rect 28870 64690 28930 64700
rect 28870 63060 28900 64690
rect 28960 64240 28990 65870
rect 28930 64230 28990 64240
rect 28930 64160 28990 64170
rect 28870 63050 28930 63060
rect 28870 62980 28930 62990
rect 28870 61350 28900 62980
rect 28960 62530 28990 64160
rect 28930 62520 28990 62530
rect 28930 62450 28990 62460
rect 28870 61340 28930 61350
rect 28870 61270 28930 61280
rect 28870 59640 28900 61270
rect 28960 60820 28990 62450
rect 28930 60810 28990 60820
rect 28930 60740 28990 60750
rect 28870 59630 28930 59640
rect 28870 59560 28930 59570
rect 28870 57930 28900 59560
rect 28960 59110 28990 60740
rect 28930 59100 28990 59110
rect 28930 59030 28990 59040
rect 28870 57920 28930 57930
rect 28870 57850 28930 57860
rect 28870 56220 28900 57850
rect 28960 57400 28990 59030
rect 28930 57390 28990 57400
rect 28930 57320 28990 57330
rect 28870 56210 28930 56220
rect 28870 56140 28930 56150
rect 28870 54510 28900 56140
rect 28960 55690 28990 57320
rect 28930 55680 28990 55690
rect 28930 55610 28990 55620
rect 28870 54500 28930 54510
rect 28870 54430 28930 54440
rect 28870 52800 28900 54430
rect 28960 53980 28990 55610
rect 28930 53970 28990 53980
rect 28930 53900 28990 53910
rect 28870 52790 28930 52800
rect 28870 52720 28930 52730
rect 28870 51090 28900 52720
rect 28960 52270 28990 53900
rect 28930 52260 28990 52270
rect 28930 52190 28990 52200
rect 28870 51080 28930 51090
rect 28870 51010 28930 51020
rect 28870 49380 28900 51010
rect 28960 50560 28990 52190
rect 28930 50550 28990 50560
rect 28930 50480 28990 50490
rect 28870 49370 28930 49380
rect 28870 49300 28930 49310
rect 28870 47670 28900 49300
rect 28960 48850 28990 50480
rect 28930 48840 28990 48850
rect 28930 48770 28990 48780
rect 28870 47660 28930 47670
rect 28870 47590 28930 47600
rect 28870 45960 28900 47590
rect 28960 47140 28990 48770
rect 28930 47130 28990 47140
rect 28930 47060 28990 47070
rect 28870 45950 28930 45960
rect 28870 45880 28930 45890
rect 28870 44250 28900 45880
rect 28960 45430 28990 47060
rect 28930 45420 28990 45430
rect 28930 45350 28990 45360
rect 28870 44240 28930 44250
rect 28870 44170 28930 44180
rect 28870 42540 28900 44170
rect 28960 43720 28990 45350
rect 28930 43710 28990 43720
rect 28930 43640 28990 43650
rect 28870 42530 28930 42540
rect 28870 42460 28930 42470
rect 28870 40830 28900 42460
rect 28960 42010 28990 43640
rect 28930 42000 28990 42010
rect 28930 41930 28990 41940
rect 28870 40820 28930 40830
rect 28870 40750 28930 40760
rect 27220 39220 27280 39230
rect 27400 39230 27660 39240
rect 24230 39160 24290 39170
rect 27460 39210 27660 39230
rect 27400 39160 27460 39170
rect 28870 38840 28900 40750
rect 28960 40300 28990 41930
rect 28930 40290 28990 40300
rect 28930 40220 28990 40230
rect 28960 39690 28990 40220
rect 28930 39680 28990 39690
rect 28930 39610 28990 39620
rect 29020 66390 29050 67050
rect 29020 66380 29080 66390
rect 29020 66310 29080 66320
rect 29020 64680 29050 66310
rect 29020 64670 29080 64680
rect 29020 64600 29080 64610
rect 29020 42450 29050 64600
rect 29140 62970 29170 67050
rect 29140 62960 29200 62970
rect 29140 62890 29200 62900
rect 29140 61250 29170 62890
rect 29140 61240 29200 61250
rect 29140 61170 29200 61180
rect 29140 45870 29170 61170
rect 29260 59550 29290 67050
rect 29260 59540 29320 59550
rect 29260 59470 29320 59480
rect 29260 47580 29290 59470
rect 29380 57840 29410 67050
rect 29380 57830 29440 57840
rect 29380 57760 29440 57770
rect 29380 56130 29410 57760
rect 29380 56120 29440 56130
rect 29380 56050 29440 56060
rect 29380 54420 29410 56050
rect 29380 54410 29440 54420
rect 29380 54340 29440 54350
rect 29380 52710 29410 54340
rect 29380 52700 29440 52710
rect 29380 52630 29440 52640
rect 29380 51000 29410 52630
rect 29380 50990 29440 51000
rect 29380 50920 29440 50930
rect 29380 49290 29410 50920
rect 29380 49280 29440 49290
rect 29380 49210 29440 49220
rect 29260 47570 29320 47580
rect 29260 47500 29320 47510
rect 29140 45860 29200 45870
rect 29140 45790 29200 45800
rect 29140 44160 29170 45790
rect 29140 44150 29200 44160
rect 29140 44080 29200 44090
rect 29020 42440 29080 42450
rect 29020 42370 29080 42380
rect 29020 40740 29050 42370
rect 29020 40730 29080 40740
rect 29020 40660 29080 40670
rect 29020 39240 29050 40660
rect 29140 39300 29170 44080
rect 29260 39360 29290 47500
rect 29380 39420 29410 49210
rect 29500 39690 29530 67050
rect 29620 39690 29650 67050
rect 29740 39690 29770 67050
rect 31900 39690 31930 67050
rect 32020 54420 32050 67050
rect 32140 56130 32170 67050
rect 32260 57840 32290 67050
rect 32380 59550 32410 67050
rect 32500 62970 32530 67050
rect 32620 66390 32650 67050
rect 32590 66380 32650 66390
rect 32590 66310 32650 66320
rect 32620 64680 32650 66310
rect 32590 64670 32650 64680
rect 32590 64600 32650 64610
rect 32470 62960 32530 62970
rect 32470 62890 32530 62900
rect 32500 61260 32530 62890
rect 32470 61250 32530 61260
rect 32470 61180 32530 61190
rect 32350 59540 32410 59550
rect 32350 59470 32410 59480
rect 32230 57830 32290 57840
rect 32230 57760 32290 57770
rect 32110 56120 32170 56130
rect 32110 56050 32170 56060
rect 31990 54410 32050 54420
rect 31990 54340 32050 54350
rect 32020 52710 32050 54340
rect 31990 52700 32050 52710
rect 31990 52630 32050 52640
rect 32020 39540 32050 52630
rect 32140 51000 32170 56050
rect 32110 50990 32170 51000
rect 32110 50920 32170 50930
rect 31490 39530 32050 39540
rect 31550 39510 32050 39530
rect 32140 39480 32170 50920
rect 32260 49290 32290 57760
rect 32230 49280 32290 49290
rect 32230 49210 32290 49220
rect 31490 39460 31550 39470
rect 31670 39470 32170 39480
rect 29380 39410 29820 39420
rect 29380 39390 29760 39410
rect 29260 39350 29640 39360
rect 29260 39330 29580 39350
rect 29140 39290 29460 39300
rect 29140 39270 29400 39290
rect 29020 39230 29280 39240
rect 29020 39210 29220 39230
rect 31730 39450 32170 39470
rect 32260 39420 32290 49210
rect 32380 47580 32410 59470
rect 32350 47570 32410 47580
rect 32350 47500 32410 47510
rect 31670 39400 31730 39410
rect 31850 39410 32290 39420
rect 29760 39340 29820 39350
rect 31910 39390 32290 39410
rect 32380 39360 32410 47500
rect 32500 45870 32530 61180
rect 32470 45860 32530 45870
rect 32470 45790 32530 45800
rect 32500 44160 32530 45790
rect 32470 44150 32530 44160
rect 32470 44080 32530 44090
rect 31850 39340 31910 39350
rect 32030 39350 32410 39360
rect 29580 39280 29640 39290
rect 32090 39330 32410 39350
rect 32500 39300 32530 44080
rect 32620 42450 32650 64600
rect 32590 42440 32650 42450
rect 32590 42370 32650 42380
rect 32620 40740 32650 42370
rect 32590 40730 32650 40740
rect 32590 40660 32650 40670
rect 32030 39280 32090 39290
rect 32210 39290 32530 39300
rect 29400 39220 29460 39230
rect 32270 39270 32530 39290
rect 32620 39240 32650 40660
rect 32680 66470 32750 67050
rect 32680 66210 32700 66470
rect 32740 66210 32750 66470
rect 33760 66470 33830 67050
rect 33210 66440 33290 66450
rect 32900 66402 33100 66408
rect 32790 66370 32870 66390
rect 32790 66310 32800 66370
rect 32860 66358 32870 66370
rect 32900 66368 32912 66402
rect 33088 66400 33100 66402
rect 33210 66400 33220 66440
rect 33088 66380 33220 66400
rect 33280 66400 33290 66440
rect 33398 66402 33598 66408
rect 33398 66400 33410 66402
rect 33280 66380 33410 66400
rect 33088 66370 33410 66380
rect 33088 66368 33100 66370
rect 32900 66362 33100 66368
rect 33398 66368 33410 66370
rect 33586 66368 33598 66402
rect 33398 66362 33598 66368
rect 33630 66370 33710 66390
rect 32862 66324 32870 66358
rect 32860 66310 32870 66324
rect 32790 66290 32870 66310
rect 32900 66314 33100 66320
rect 32900 66280 32912 66314
rect 33088 66310 33100 66314
rect 33398 66314 33598 66320
rect 33398 66310 33410 66314
rect 33088 66280 33410 66310
rect 33586 66280 33598 66314
rect 33630 66310 33640 66370
rect 33700 66310 33710 66370
rect 33630 66290 33710 66310
rect 32900 66274 33100 66280
rect 32680 66150 32750 66210
rect 32680 65910 32700 66150
rect 32740 65910 32750 66150
rect 33210 66270 33290 66280
rect 33398 66274 33598 66280
rect 33210 66210 33220 66270
rect 33280 66210 33290 66270
rect 33210 66160 33290 66210
rect 33210 66100 33220 66160
rect 33280 66100 33290 66160
rect 32900 66092 33100 66098
rect 32790 66060 32870 66080
rect 32790 66000 32800 66060
rect 32860 66048 32870 66060
rect 32900 66058 32912 66092
rect 33088 66090 33100 66092
rect 33210 66090 33290 66100
rect 33760 66230 33770 66470
rect 33810 66230 33830 66470
rect 33760 66150 33830 66230
rect 33398 66092 33598 66098
rect 33398 66090 33410 66092
rect 33088 66060 33410 66090
rect 33088 66058 33100 66060
rect 32900 66052 33100 66058
rect 33398 66058 33410 66060
rect 33586 66058 33598 66092
rect 33398 66052 33598 66058
rect 33630 66060 33710 66080
rect 32862 66014 32870 66048
rect 32860 66000 32870 66014
rect 32790 65980 32870 66000
rect 32900 66004 33100 66010
rect 32900 65970 32912 66004
rect 33088 66000 33100 66004
rect 33398 66004 33598 66010
rect 33398 66000 33410 66004
rect 33088 65990 33410 66000
rect 33088 65970 33220 65990
rect 32900 65964 33100 65970
rect 33210 65930 33220 65970
rect 33280 65970 33410 65990
rect 33586 65970 33598 66004
rect 33630 66000 33640 66060
rect 33700 66000 33710 66060
rect 33630 65980 33710 66000
rect 33280 65930 33290 65970
rect 33398 65964 33598 65970
rect 33210 65920 33290 65930
rect 32680 64760 32750 65910
rect 32680 64500 32700 64760
rect 32740 64500 32750 64760
rect 33760 65910 33770 66150
rect 33810 65910 33830 66150
rect 33760 64760 33830 65910
rect 33210 64730 33290 64740
rect 32900 64692 33100 64698
rect 32790 64660 32870 64680
rect 32790 64600 32800 64660
rect 32860 64648 32870 64660
rect 32900 64658 32912 64692
rect 33088 64690 33100 64692
rect 33210 64690 33220 64730
rect 33088 64670 33220 64690
rect 33280 64690 33290 64730
rect 33398 64692 33598 64698
rect 33398 64690 33410 64692
rect 33280 64670 33410 64690
rect 33088 64660 33410 64670
rect 33088 64658 33100 64660
rect 32900 64652 33100 64658
rect 33398 64658 33410 64660
rect 33586 64658 33598 64692
rect 33398 64652 33598 64658
rect 33630 64660 33710 64680
rect 32862 64614 32870 64648
rect 32860 64600 32870 64614
rect 32790 64580 32870 64600
rect 32900 64604 33100 64610
rect 32900 64570 32912 64604
rect 33088 64600 33100 64604
rect 33398 64604 33598 64610
rect 33398 64600 33410 64604
rect 33088 64570 33410 64600
rect 33586 64570 33598 64604
rect 33630 64600 33640 64660
rect 33700 64600 33710 64660
rect 33630 64580 33710 64600
rect 32900 64564 33100 64570
rect 32680 64440 32750 64500
rect 32680 64200 32700 64440
rect 32740 64200 32750 64440
rect 33210 64560 33290 64570
rect 33398 64564 33598 64570
rect 33210 64500 33220 64560
rect 33280 64500 33290 64560
rect 33210 64450 33290 64500
rect 33210 64390 33220 64450
rect 33280 64390 33290 64450
rect 32900 64382 33100 64388
rect 32790 64350 32870 64370
rect 32790 64290 32800 64350
rect 32860 64338 32870 64350
rect 32900 64348 32912 64382
rect 33088 64380 33100 64382
rect 33210 64380 33290 64390
rect 33760 64520 33770 64760
rect 33810 64520 33830 64760
rect 33760 64440 33830 64520
rect 33398 64382 33598 64388
rect 33398 64380 33410 64382
rect 33088 64350 33410 64380
rect 33088 64348 33100 64350
rect 32900 64342 33100 64348
rect 33398 64348 33410 64350
rect 33586 64348 33598 64382
rect 33398 64342 33598 64348
rect 33630 64350 33710 64370
rect 32862 64304 32870 64338
rect 32860 64290 32870 64304
rect 32790 64270 32870 64290
rect 32900 64294 33100 64300
rect 32900 64260 32912 64294
rect 33088 64290 33100 64294
rect 33398 64294 33598 64300
rect 33398 64290 33410 64294
rect 33088 64280 33410 64290
rect 33088 64260 33220 64280
rect 32900 64254 33100 64260
rect 33210 64220 33220 64260
rect 33280 64260 33410 64280
rect 33586 64260 33598 64294
rect 33630 64290 33640 64350
rect 33700 64290 33710 64350
rect 33630 64270 33710 64290
rect 33280 64220 33290 64260
rect 33398 64254 33598 64260
rect 33210 64210 33290 64220
rect 32680 63050 32750 64200
rect 32680 62790 32700 63050
rect 32740 62790 32750 63050
rect 33760 64200 33770 64440
rect 33810 64200 33830 64440
rect 33760 63050 33830 64200
rect 33210 63020 33290 63030
rect 32900 62982 33100 62988
rect 32790 62950 32870 62970
rect 32790 62890 32800 62950
rect 32860 62938 32870 62950
rect 32900 62948 32912 62982
rect 33088 62980 33100 62982
rect 33210 62980 33220 63020
rect 33088 62960 33220 62980
rect 33280 62980 33290 63020
rect 33398 62982 33598 62988
rect 33398 62980 33410 62982
rect 33280 62960 33410 62980
rect 33088 62950 33410 62960
rect 33088 62948 33100 62950
rect 32900 62942 33100 62948
rect 33398 62948 33410 62950
rect 33586 62948 33598 62982
rect 33398 62942 33598 62948
rect 33630 62950 33710 62970
rect 32862 62904 32870 62938
rect 32860 62890 32870 62904
rect 32790 62870 32870 62890
rect 32900 62894 33100 62900
rect 32900 62860 32912 62894
rect 33088 62890 33100 62894
rect 33398 62894 33598 62900
rect 33398 62890 33410 62894
rect 33088 62860 33410 62890
rect 33586 62860 33598 62894
rect 33630 62890 33640 62950
rect 33700 62890 33710 62950
rect 33630 62870 33710 62890
rect 32900 62854 33100 62860
rect 32680 62730 32750 62790
rect 32680 62490 32700 62730
rect 32740 62490 32750 62730
rect 33210 62850 33290 62860
rect 33398 62854 33598 62860
rect 33210 62790 33220 62850
rect 33280 62790 33290 62850
rect 33210 62740 33290 62790
rect 33210 62680 33220 62740
rect 33280 62680 33290 62740
rect 32900 62672 33100 62678
rect 32790 62640 32870 62660
rect 32790 62580 32800 62640
rect 32860 62628 32870 62640
rect 32900 62638 32912 62672
rect 33088 62670 33100 62672
rect 33210 62670 33290 62680
rect 33760 62810 33770 63050
rect 33810 62810 33830 63050
rect 33760 62730 33830 62810
rect 33398 62672 33598 62678
rect 33398 62670 33410 62672
rect 33088 62640 33410 62670
rect 33088 62638 33100 62640
rect 32900 62632 33100 62638
rect 33398 62638 33410 62640
rect 33586 62638 33598 62672
rect 33398 62632 33598 62638
rect 33630 62640 33710 62660
rect 32862 62594 32870 62628
rect 32860 62580 32870 62594
rect 32790 62560 32870 62580
rect 32900 62584 33100 62590
rect 32900 62550 32912 62584
rect 33088 62580 33100 62584
rect 33398 62584 33598 62590
rect 33398 62580 33410 62584
rect 33088 62570 33410 62580
rect 33088 62550 33220 62570
rect 32900 62544 33100 62550
rect 33210 62510 33220 62550
rect 33280 62550 33410 62570
rect 33586 62550 33598 62584
rect 33630 62580 33640 62640
rect 33700 62580 33710 62640
rect 33630 62560 33710 62580
rect 33280 62510 33290 62550
rect 33398 62544 33598 62550
rect 33210 62500 33290 62510
rect 32680 61340 32750 62490
rect 32680 61080 32700 61340
rect 32740 61080 32750 61340
rect 33760 62490 33770 62730
rect 33810 62490 33830 62730
rect 33760 61340 33830 62490
rect 33210 61310 33290 61320
rect 32900 61272 33100 61278
rect 32790 61240 32870 61260
rect 32790 61180 32800 61240
rect 32860 61228 32870 61240
rect 32900 61238 32912 61272
rect 33088 61270 33100 61272
rect 33210 61270 33220 61310
rect 33088 61250 33220 61270
rect 33280 61270 33290 61310
rect 33398 61272 33598 61278
rect 33398 61270 33410 61272
rect 33280 61250 33410 61270
rect 33088 61240 33410 61250
rect 33088 61238 33100 61240
rect 32900 61232 33100 61238
rect 33398 61238 33410 61240
rect 33586 61238 33598 61272
rect 33398 61232 33598 61238
rect 33630 61240 33710 61260
rect 32862 61194 32870 61228
rect 32860 61180 32870 61194
rect 32790 61160 32870 61180
rect 32900 61184 33100 61190
rect 32900 61150 32912 61184
rect 33088 61180 33100 61184
rect 33398 61184 33598 61190
rect 33398 61180 33410 61184
rect 33088 61150 33410 61180
rect 33586 61150 33598 61184
rect 33630 61180 33640 61240
rect 33700 61180 33710 61240
rect 33630 61160 33710 61180
rect 32900 61144 33100 61150
rect 32680 61020 32750 61080
rect 32680 60780 32700 61020
rect 32740 60780 32750 61020
rect 33210 61140 33290 61150
rect 33398 61144 33598 61150
rect 33210 61080 33220 61140
rect 33280 61080 33290 61140
rect 33210 61030 33290 61080
rect 33210 60970 33220 61030
rect 33280 60970 33290 61030
rect 32900 60962 33100 60968
rect 32790 60930 32870 60950
rect 32790 60870 32800 60930
rect 32860 60918 32870 60930
rect 32900 60928 32912 60962
rect 33088 60960 33100 60962
rect 33210 60960 33290 60970
rect 33760 61100 33770 61340
rect 33810 61100 33830 61340
rect 33760 61020 33830 61100
rect 33398 60962 33598 60968
rect 33398 60960 33410 60962
rect 33088 60930 33410 60960
rect 33088 60928 33100 60930
rect 32900 60922 33100 60928
rect 33398 60928 33410 60930
rect 33586 60928 33598 60962
rect 33398 60922 33598 60928
rect 33630 60930 33710 60950
rect 32862 60884 32870 60918
rect 32860 60870 32870 60884
rect 32790 60850 32870 60870
rect 32900 60874 33100 60880
rect 32900 60840 32912 60874
rect 33088 60870 33100 60874
rect 33398 60874 33598 60880
rect 33398 60870 33410 60874
rect 33088 60860 33410 60870
rect 33088 60840 33220 60860
rect 32900 60834 33100 60840
rect 33210 60800 33220 60840
rect 33280 60840 33410 60860
rect 33586 60840 33598 60874
rect 33630 60870 33640 60930
rect 33700 60870 33710 60930
rect 33630 60850 33710 60870
rect 33280 60800 33290 60840
rect 33398 60834 33598 60840
rect 33210 60790 33290 60800
rect 32680 59630 32750 60780
rect 32680 59370 32700 59630
rect 32740 59370 32750 59630
rect 33760 60780 33770 61020
rect 33810 60780 33830 61020
rect 33760 59630 33830 60780
rect 33210 59600 33290 59610
rect 32900 59562 33100 59568
rect 32790 59530 32870 59550
rect 32790 59470 32800 59530
rect 32860 59518 32870 59530
rect 32900 59528 32912 59562
rect 33088 59560 33100 59562
rect 33210 59560 33220 59600
rect 33088 59540 33220 59560
rect 33280 59560 33290 59600
rect 33398 59562 33598 59568
rect 33398 59560 33410 59562
rect 33280 59540 33410 59560
rect 33088 59530 33410 59540
rect 33088 59528 33100 59530
rect 32900 59522 33100 59528
rect 33398 59528 33410 59530
rect 33586 59528 33598 59562
rect 33398 59522 33598 59528
rect 33630 59530 33710 59550
rect 32862 59484 32870 59518
rect 32860 59470 32870 59484
rect 32790 59450 32870 59470
rect 32900 59474 33100 59480
rect 32900 59440 32912 59474
rect 33088 59470 33100 59474
rect 33398 59474 33598 59480
rect 33398 59470 33410 59474
rect 33088 59440 33410 59470
rect 33586 59440 33598 59474
rect 33630 59470 33640 59530
rect 33700 59470 33710 59530
rect 33630 59450 33710 59470
rect 32900 59434 33100 59440
rect 32680 59310 32750 59370
rect 32680 59070 32700 59310
rect 32740 59070 32750 59310
rect 33210 59430 33290 59440
rect 33398 59434 33598 59440
rect 33210 59370 33220 59430
rect 33280 59370 33290 59430
rect 33210 59320 33290 59370
rect 33210 59260 33220 59320
rect 33280 59260 33290 59320
rect 32900 59252 33100 59258
rect 32790 59220 32870 59240
rect 32790 59160 32800 59220
rect 32860 59208 32870 59220
rect 32900 59218 32912 59252
rect 33088 59250 33100 59252
rect 33210 59250 33290 59260
rect 33760 59390 33770 59630
rect 33810 59390 33830 59630
rect 33760 59310 33830 59390
rect 33398 59252 33598 59258
rect 33398 59250 33410 59252
rect 33088 59220 33410 59250
rect 33088 59218 33100 59220
rect 32900 59212 33100 59218
rect 33398 59218 33410 59220
rect 33586 59218 33598 59252
rect 33398 59212 33598 59218
rect 33630 59220 33710 59240
rect 32862 59174 32870 59208
rect 32860 59160 32870 59174
rect 32790 59140 32870 59160
rect 32900 59164 33100 59170
rect 32900 59130 32912 59164
rect 33088 59160 33100 59164
rect 33398 59164 33598 59170
rect 33398 59160 33410 59164
rect 33088 59150 33410 59160
rect 33088 59130 33220 59150
rect 32900 59124 33100 59130
rect 33210 59090 33220 59130
rect 33280 59130 33410 59150
rect 33586 59130 33598 59164
rect 33630 59160 33640 59220
rect 33700 59160 33710 59220
rect 33630 59140 33710 59160
rect 33280 59090 33290 59130
rect 33398 59124 33598 59130
rect 33210 59080 33290 59090
rect 32680 57920 32750 59070
rect 32680 57660 32700 57920
rect 32740 57660 32750 57920
rect 33760 59070 33770 59310
rect 33810 59070 33830 59310
rect 33760 57920 33830 59070
rect 33210 57890 33290 57900
rect 32900 57852 33100 57858
rect 32790 57820 32870 57840
rect 32790 57760 32800 57820
rect 32860 57808 32870 57820
rect 32900 57818 32912 57852
rect 33088 57850 33100 57852
rect 33210 57850 33220 57890
rect 33088 57830 33220 57850
rect 33280 57850 33290 57890
rect 33398 57852 33598 57858
rect 33398 57850 33410 57852
rect 33280 57830 33410 57850
rect 33088 57820 33410 57830
rect 33088 57818 33100 57820
rect 32900 57812 33100 57818
rect 33398 57818 33410 57820
rect 33586 57818 33598 57852
rect 33398 57812 33598 57818
rect 33630 57820 33710 57840
rect 32862 57774 32870 57808
rect 32860 57760 32870 57774
rect 32790 57740 32870 57760
rect 32900 57764 33100 57770
rect 32900 57730 32912 57764
rect 33088 57760 33100 57764
rect 33398 57764 33598 57770
rect 33398 57760 33410 57764
rect 33088 57730 33410 57760
rect 33586 57730 33598 57764
rect 33630 57760 33640 57820
rect 33700 57760 33710 57820
rect 33630 57740 33710 57760
rect 32900 57724 33100 57730
rect 32680 57600 32750 57660
rect 32680 57360 32700 57600
rect 32740 57360 32750 57600
rect 33210 57720 33290 57730
rect 33398 57724 33598 57730
rect 33210 57660 33220 57720
rect 33280 57660 33290 57720
rect 33210 57610 33290 57660
rect 33210 57550 33220 57610
rect 33280 57550 33290 57610
rect 32900 57542 33100 57548
rect 32790 57510 32870 57530
rect 32790 57450 32800 57510
rect 32860 57498 32870 57510
rect 32900 57508 32912 57542
rect 33088 57540 33100 57542
rect 33210 57540 33290 57550
rect 33760 57680 33770 57920
rect 33810 57680 33830 57920
rect 33760 57600 33830 57680
rect 33398 57542 33598 57548
rect 33398 57540 33410 57542
rect 33088 57510 33410 57540
rect 33088 57508 33100 57510
rect 32900 57502 33100 57508
rect 33398 57508 33410 57510
rect 33586 57508 33598 57542
rect 33398 57502 33598 57508
rect 33630 57510 33710 57530
rect 32862 57464 32870 57498
rect 32860 57450 32870 57464
rect 32790 57430 32870 57450
rect 32900 57454 33100 57460
rect 32900 57420 32912 57454
rect 33088 57450 33100 57454
rect 33398 57454 33598 57460
rect 33398 57450 33410 57454
rect 33088 57440 33410 57450
rect 33088 57420 33220 57440
rect 32900 57414 33100 57420
rect 33210 57380 33220 57420
rect 33280 57420 33410 57440
rect 33586 57420 33598 57454
rect 33630 57450 33640 57510
rect 33700 57450 33710 57510
rect 33630 57430 33710 57450
rect 33280 57380 33290 57420
rect 33398 57414 33598 57420
rect 33210 57370 33290 57380
rect 32680 56210 32750 57360
rect 32680 55950 32700 56210
rect 32740 55950 32750 56210
rect 33760 57360 33770 57600
rect 33810 57360 33830 57600
rect 33760 56210 33830 57360
rect 33210 56180 33290 56190
rect 32900 56142 33100 56148
rect 32790 56110 32870 56130
rect 32790 56050 32800 56110
rect 32860 56098 32870 56110
rect 32900 56108 32912 56142
rect 33088 56140 33100 56142
rect 33210 56140 33220 56180
rect 33088 56120 33220 56140
rect 33280 56140 33290 56180
rect 33398 56142 33598 56148
rect 33398 56140 33410 56142
rect 33280 56120 33410 56140
rect 33088 56110 33410 56120
rect 33088 56108 33100 56110
rect 32900 56102 33100 56108
rect 33398 56108 33410 56110
rect 33586 56108 33598 56142
rect 33398 56102 33598 56108
rect 33630 56110 33710 56130
rect 32862 56064 32870 56098
rect 32860 56050 32870 56064
rect 32790 56030 32870 56050
rect 32900 56054 33100 56060
rect 32900 56020 32912 56054
rect 33088 56050 33100 56054
rect 33398 56054 33598 56060
rect 33398 56050 33410 56054
rect 33088 56020 33410 56050
rect 33586 56020 33598 56054
rect 33630 56050 33640 56110
rect 33700 56050 33710 56110
rect 33630 56030 33710 56050
rect 32900 56014 33100 56020
rect 32680 55890 32750 55950
rect 32680 55650 32700 55890
rect 32740 55650 32750 55890
rect 33210 56010 33290 56020
rect 33398 56014 33598 56020
rect 33210 55950 33220 56010
rect 33280 55950 33290 56010
rect 33210 55900 33290 55950
rect 33210 55840 33220 55900
rect 33280 55840 33290 55900
rect 32900 55832 33100 55838
rect 32790 55800 32870 55820
rect 32790 55740 32800 55800
rect 32860 55788 32870 55800
rect 32900 55798 32912 55832
rect 33088 55830 33100 55832
rect 33210 55830 33290 55840
rect 33760 55970 33770 56210
rect 33810 55970 33830 56210
rect 33760 55890 33830 55970
rect 33398 55832 33598 55838
rect 33398 55830 33410 55832
rect 33088 55800 33410 55830
rect 33088 55798 33100 55800
rect 32900 55792 33100 55798
rect 33398 55798 33410 55800
rect 33586 55798 33598 55832
rect 33398 55792 33598 55798
rect 33630 55800 33710 55820
rect 32862 55754 32870 55788
rect 32860 55740 32870 55754
rect 32790 55720 32870 55740
rect 32900 55744 33100 55750
rect 32900 55710 32912 55744
rect 33088 55740 33100 55744
rect 33398 55744 33598 55750
rect 33398 55740 33410 55744
rect 33088 55730 33410 55740
rect 33088 55710 33220 55730
rect 32900 55704 33100 55710
rect 33210 55670 33220 55710
rect 33280 55710 33410 55730
rect 33586 55710 33598 55744
rect 33630 55740 33640 55800
rect 33700 55740 33710 55800
rect 33630 55720 33710 55740
rect 33280 55670 33290 55710
rect 33398 55704 33598 55710
rect 33210 55660 33290 55670
rect 32680 54500 32750 55650
rect 32680 54240 32700 54500
rect 32740 54240 32750 54500
rect 33760 55650 33770 55890
rect 33810 55650 33830 55890
rect 33760 54500 33830 55650
rect 33210 54470 33290 54480
rect 32900 54432 33100 54438
rect 32790 54400 32870 54420
rect 32790 54340 32800 54400
rect 32860 54388 32870 54400
rect 32900 54398 32912 54432
rect 33088 54430 33100 54432
rect 33210 54430 33220 54470
rect 33088 54410 33220 54430
rect 33280 54430 33290 54470
rect 33398 54432 33598 54438
rect 33398 54430 33410 54432
rect 33280 54410 33410 54430
rect 33088 54400 33410 54410
rect 33088 54398 33100 54400
rect 32900 54392 33100 54398
rect 33398 54398 33410 54400
rect 33586 54398 33598 54432
rect 33398 54392 33598 54398
rect 33630 54400 33710 54420
rect 32862 54354 32870 54388
rect 32860 54340 32870 54354
rect 32790 54320 32870 54340
rect 32900 54344 33100 54350
rect 32900 54310 32912 54344
rect 33088 54340 33100 54344
rect 33398 54344 33598 54350
rect 33398 54340 33410 54344
rect 33088 54310 33410 54340
rect 33586 54310 33598 54344
rect 33630 54340 33640 54400
rect 33700 54340 33710 54400
rect 33630 54320 33710 54340
rect 32900 54304 33100 54310
rect 32680 54180 32750 54240
rect 32680 53940 32700 54180
rect 32740 53940 32750 54180
rect 33210 54300 33290 54310
rect 33398 54304 33598 54310
rect 33210 54240 33220 54300
rect 33280 54240 33290 54300
rect 33210 54190 33290 54240
rect 33210 54130 33220 54190
rect 33280 54130 33290 54190
rect 32900 54122 33100 54128
rect 32790 54090 32870 54110
rect 32790 54030 32800 54090
rect 32860 54078 32870 54090
rect 32900 54088 32912 54122
rect 33088 54120 33100 54122
rect 33210 54120 33290 54130
rect 33760 54260 33770 54500
rect 33810 54260 33830 54500
rect 33760 54180 33830 54260
rect 33398 54122 33598 54128
rect 33398 54120 33410 54122
rect 33088 54090 33410 54120
rect 33088 54088 33100 54090
rect 32900 54082 33100 54088
rect 33398 54088 33410 54090
rect 33586 54088 33598 54122
rect 33398 54082 33598 54088
rect 33630 54090 33710 54110
rect 32862 54044 32870 54078
rect 32860 54030 32870 54044
rect 32790 54010 32870 54030
rect 32900 54034 33100 54040
rect 32900 54000 32912 54034
rect 33088 54030 33100 54034
rect 33398 54034 33598 54040
rect 33398 54030 33410 54034
rect 33088 54020 33410 54030
rect 33088 54000 33220 54020
rect 32900 53994 33100 54000
rect 33210 53960 33220 54000
rect 33280 54000 33410 54020
rect 33586 54000 33598 54034
rect 33630 54030 33640 54090
rect 33700 54030 33710 54090
rect 33630 54010 33710 54030
rect 33280 53960 33290 54000
rect 33398 53994 33598 54000
rect 33210 53950 33290 53960
rect 32680 52790 32750 53940
rect 32680 52530 32700 52790
rect 32740 52530 32750 52790
rect 33760 53940 33770 54180
rect 33810 53940 33830 54180
rect 33760 52790 33830 53940
rect 33210 52760 33290 52770
rect 32900 52722 33100 52728
rect 32790 52690 32870 52710
rect 32790 52630 32800 52690
rect 32860 52678 32870 52690
rect 32900 52688 32912 52722
rect 33088 52720 33100 52722
rect 33210 52720 33220 52760
rect 33088 52700 33220 52720
rect 33280 52720 33290 52760
rect 33398 52722 33598 52728
rect 33398 52720 33410 52722
rect 33280 52700 33410 52720
rect 33088 52690 33410 52700
rect 33088 52688 33100 52690
rect 32900 52682 33100 52688
rect 33398 52688 33410 52690
rect 33586 52688 33598 52722
rect 33398 52682 33598 52688
rect 33630 52690 33710 52710
rect 32862 52644 32870 52678
rect 32860 52630 32870 52644
rect 32790 52610 32870 52630
rect 32900 52634 33100 52640
rect 32900 52600 32912 52634
rect 33088 52630 33100 52634
rect 33398 52634 33598 52640
rect 33398 52630 33410 52634
rect 33088 52600 33410 52630
rect 33586 52600 33598 52634
rect 33630 52630 33640 52690
rect 33700 52630 33710 52690
rect 33630 52610 33710 52630
rect 32900 52594 33100 52600
rect 32680 52470 32750 52530
rect 32680 52230 32700 52470
rect 32740 52230 32750 52470
rect 33210 52590 33290 52600
rect 33398 52594 33598 52600
rect 33210 52530 33220 52590
rect 33280 52530 33290 52590
rect 33210 52480 33290 52530
rect 33210 52420 33220 52480
rect 33280 52420 33290 52480
rect 32900 52412 33100 52418
rect 32790 52380 32870 52400
rect 32790 52320 32800 52380
rect 32860 52368 32870 52380
rect 32900 52378 32912 52412
rect 33088 52410 33100 52412
rect 33210 52410 33290 52420
rect 33760 52550 33770 52790
rect 33810 52550 33830 52790
rect 33760 52470 33830 52550
rect 33398 52412 33598 52418
rect 33398 52410 33410 52412
rect 33088 52380 33410 52410
rect 33088 52378 33100 52380
rect 32900 52372 33100 52378
rect 33398 52378 33410 52380
rect 33586 52378 33598 52412
rect 33398 52372 33598 52378
rect 33630 52380 33710 52400
rect 32862 52334 32870 52368
rect 32860 52320 32870 52334
rect 32790 52300 32870 52320
rect 32900 52324 33100 52330
rect 32900 52290 32912 52324
rect 33088 52320 33100 52324
rect 33398 52324 33598 52330
rect 33398 52320 33410 52324
rect 33088 52310 33410 52320
rect 33088 52290 33220 52310
rect 32900 52284 33100 52290
rect 33210 52250 33220 52290
rect 33280 52290 33410 52310
rect 33586 52290 33598 52324
rect 33630 52320 33640 52380
rect 33700 52320 33710 52380
rect 33630 52300 33710 52320
rect 33280 52250 33290 52290
rect 33398 52284 33598 52290
rect 33210 52240 33290 52250
rect 32680 51080 32750 52230
rect 32680 50820 32700 51080
rect 32740 50820 32750 51080
rect 33760 52230 33770 52470
rect 33810 52230 33830 52470
rect 33760 51080 33830 52230
rect 33210 51050 33290 51060
rect 32900 51012 33100 51018
rect 32790 50980 32870 51000
rect 32790 50920 32800 50980
rect 32860 50968 32870 50980
rect 32900 50978 32912 51012
rect 33088 51010 33100 51012
rect 33210 51010 33220 51050
rect 33088 50990 33220 51010
rect 33280 51010 33290 51050
rect 33398 51012 33598 51018
rect 33398 51010 33410 51012
rect 33280 50990 33410 51010
rect 33088 50980 33410 50990
rect 33088 50978 33100 50980
rect 32900 50972 33100 50978
rect 33398 50978 33410 50980
rect 33586 50978 33598 51012
rect 33398 50972 33598 50978
rect 33630 50980 33710 51000
rect 32862 50934 32870 50968
rect 32860 50920 32870 50934
rect 32790 50900 32870 50920
rect 32900 50924 33100 50930
rect 32900 50890 32912 50924
rect 33088 50920 33100 50924
rect 33398 50924 33598 50930
rect 33398 50920 33410 50924
rect 33088 50890 33410 50920
rect 33586 50890 33598 50924
rect 33630 50920 33640 50980
rect 33700 50920 33710 50980
rect 33630 50900 33710 50920
rect 32900 50884 33100 50890
rect 32680 50760 32750 50820
rect 32680 50520 32700 50760
rect 32740 50520 32750 50760
rect 33210 50880 33290 50890
rect 33398 50884 33598 50890
rect 33210 50820 33220 50880
rect 33280 50820 33290 50880
rect 33210 50770 33290 50820
rect 33210 50710 33220 50770
rect 33280 50710 33290 50770
rect 32900 50702 33100 50708
rect 32790 50670 32870 50690
rect 32790 50610 32800 50670
rect 32860 50658 32870 50670
rect 32900 50668 32912 50702
rect 33088 50700 33100 50702
rect 33210 50700 33290 50710
rect 33760 50840 33770 51080
rect 33810 50840 33830 51080
rect 33760 50760 33830 50840
rect 33398 50702 33598 50708
rect 33398 50700 33410 50702
rect 33088 50670 33410 50700
rect 33088 50668 33100 50670
rect 32900 50662 33100 50668
rect 33398 50668 33410 50670
rect 33586 50668 33598 50702
rect 33398 50662 33598 50668
rect 33630 50670 33710 50690
rect 32862 50624 32870 50658
rect 32860 50610 32870 50624
rect 32790 50590 32870 50610
rect 32900 50614 33100 50620
rect 32900 50580 32912 50614
rect 33088 50610 33100 50614
rect 33398 50614 33598 50620
rect 33398 50610 33410 50614
rect 33088 50600 33410 50610
rect 33088 50580 33220 50600
rect 32900 50574 33100 50580
rect 33210 50540 33220 50580
rect 33280 50580 33410 50600
rect 33586 50580 33598 50614
rect 33630 50610 33640 50670
rect 33700 50610 33710 50670
rect 33630 50590 33710 50610
rect 33280 50540 33290 50580
rect 33398 50574 33598 50580
rect 33210 50530 33290 50540
rect 32680 49370 32750 50520
rect 32680 49110 32700 49370
rect 32740 49110 32750 49370
rect 33760 50520 33770 50760
rect 33810 50520 33830 50760
rect 33760 49370 33830 50520
rect 33210 49340 33290 49350
rect 32900 49302 33100 49308
rect 32790 49270 32870 49290
rect 32790 49210 32800 49270
rect 32860 49258 32870 49270
rect 32900 49268 32912 49302
rect 33088 49300 33100 49302
rect 33210 49300 33220 49340
rect 33088 49280 33220 49300
rect 33280 49300 33290 49340
rect 33398 49302 33598 49308
rect 33398 49300 33410 49302
rect 33280 49280 33410 49300
rect 33088 49270 33410 49280
rect 33088 49268 33100 49270
rect 32900 49262 33100 49268
rect 33398 49268 33410 49270
rect 33586 49268 33598 49302
rect 33398 49262 33598 49268
rect 33630 49270 33710 49290
rect 32862 49224 32870 49258
rect 32860 49210 32870 49224
rect 32790 49190 32870 49210
rect 32900 49214 33100 49220
rect 32900 49180 32912 49214
rect 33088 49210 33100 49214
rect 33398 49214 33598 49220
rect 33398 49210 33410 49214
rect 33088 49180 33410 49210
rect 33586 49180 33598 49214
rect 33630 49210 33640 49270
rect 33700 49210 33710 49270
rect 33630 49190 33710 49210
rect 32900 49174 33100 49180
rect 32680 49050 32750 49110
rect 32680 48810 32700 49050
rect 32740 48810 32750 49050
rect 33210 49170 33290 49180
rect 33398 49174 33598 49180
rect 33210 49110 33220 49170
rect 33280 49110 33290 49170
rect 33210 49060 33290 49110
rect 33210 49000 33220 49060
rect 33280 49000 33290 49060
rect 32900 48992 33100 48998
rect 32790 48960 32870 48980
rect 32790 48900 32800 48960
rect 32860 48948 32870 48960
rect 32900 48958 32912 48992
rect 33088 48990 33100 48992
rect 33210 48990 33290 49000
rect 33760 49130 33770 49370
rect 33810 49130 33830 49370
rect 33760 49050 33830 49130
rect 33398 48992 33598 48998
rect 33398 48990 33410 48992
rect 33088 48960 33410 48990
rect 33088 48958 33100 48960
rect 32900 48952 33100 48958
rect 33398 48958 33410 48960
rect 33586 48958 33598 48992
rect 33398 48952 33598 48958
rect 33630 48960 33710 48980
rect 32862 48914 32870 48948
rect 32860 48900 32870 48914
rect 32790 48880 32870 48900
rect 32900 48904 33100 48910
rect 32900 48870 32912 48904
rect 33088 48900 33100 48904
rect 33398 48904 33598 48910
rect 33398 48900 33410 48904
rect 33088 48890 33410 48900
rect 33088 48870 33220 48890
rect 32900 48864 33100 48870
rect 33210 48830 33220 48870
rect 33280 48870 33410 48890
rect 33586 48870 33598 48904
rect 33630 48900 33640 48960
rect 33700 48900 33710 48960
rect 33630 48880 33710 48900
rect 33280 48830 33290 48870
rect 33398 48864 33598 48870
rect 33210 48820 33290 48830
rect 32680 47660 32750 48810
rect 32680 47400 32700 47660
rect 32740 47400 32750 47660
rect 33760 48810 33770 49050
rect 33810 48810 33830 49050
rect 33760 47660 33830 48810
rect 33210 47630 33290 47640
rect 32900 47592 33100 47598
rect 32790 47560 32870 47580
rect 32790 47500 32800 47560
rect 32860 47548 32870 47560
rect 32900 47558 32912 47592
rect 33088 47590 33100 47592
rect 33210 47590 33220 47630
rect 33088 47570 33220 47590
rect 33280 47590 33290 47630
rect 33398 47592 33598 47598
rect 33398 47590 33410 47592
rect 33280 47570 33410 47590
rect 33088 47560 33410 47570
rect 33088 47558 33100 47560
rect 32900 47552 33100 47558
rect 33398 47558 33410 47560
rect 33586 47558 33598 47592
rect 33398 47552 33598 47558
rect 33630 47560 33710 47580
rect 32862 47514 32870 47548
rect 32860 47500 32870 47514
rect 32790 47480 32870 47500
rect 32900 47504 33100 47510
rect 32900 47470 32912 47504
rect 33088 47500 33100 47504
rect 33398 47504 33598 47510
rect 33398 47500 33410 47504
rect 33088 47470 33410 47500
rect 33586 47470 33598 47504
rect 33630 47500 33640 47560
rect 33700 47500 33710 47560
rect 33630 47480 33710 47500
rect 32900 47464 33100 47470
rect 32680 47340 32750 47400
rect 32680 47100 32700 47340
rect 32740 47100 32750 47340
rect 33210 47460 33290 47470
rect 33398 47464 33598 47470
rect 33210 47400 33220 47460
rect 33280 47400 33290 47460
rect 33210 47350 33290 47400
rect 33210 47290 33220 47350
rect 33280 47290 33290 47350
rect 32900 47282 33100 47288
rect 32790 47250 32870 47270
rect 32790 47190 32800 47250
rect 32860 47238 32870 47250
rect 32900 47248 32912 47282
rect 33088 47280 33100 47282
rect 33210 47280 33290 47290
rect 33760 47420 33770 47660
rect 33810 47420 33830 47660
rect 33760 47340 33830 47420
rect 33398 47282 33598 47288
rect 33398 47280 33410 47282
rect 33088 47250 33410 47280
rect 33088 47248 33100 47250
rect 32900 47242 33100 47248
rect 33398 47248 33410 47250
rect 33586 47248 33598 47282
rect 33398 47242 33598 47248
rect 33630 47250 33710 47270
rect 32862 47204 32870 47238
rect 32860 47190 32870 47204
rect 32790 47170 32870 47190
rect 32900 47194 33100 47200
rect 32900 47160 32912 47194
rect 33088 47190 33100 47194
rect 33398 47194 33598 47200
rect 33398 47190 33410 47194
rect 33088 47180 33410 47190
rect 33088 47160 33220 47180
rect 32900 47154 33100 47160
rect 33210 47120 33220 47160
rect 33280 47160 33410 47180
rect 33586 47160 33598 47194
rect 33630 47190 33640 47250
rect 33700 47190 33710 47250
rect 33630 47170 33710 47190
rect 33280 47120 33290 47160
rect 33398 47154 33598 47160
rect 33210 47110 33290 47120
rect 32680 45950 32750 47100
rect 32680 45690 32700 45950
rect 32740 45690 32750 45950
rect 33760 47100 33770 47340
rect 33810 47100 33830 47340
rect 33760 45950 33830 47100
rect 33210 45920 33290 45930
rect 32900 45882 33100 45888
rect 32790 45850 32870 45870
rect 32790 45790 32800 45850
rect 32860 45838 32870 45850
rect 32900 45848 32912 45882
rect 33088 45880 33100 45882
rect 33210 45880 33220 45920
rect 33088 45860 33220 45880
rect 33280 45880 33290 45920
rect 33398 45882 33598 45888
rect 33398 45880 33410 45882
rect 33280 45860 33410 45880
rect 33088 45850 33410 45860
rect 33088 45848 33100 45850
rect 32900 45842 33100 45848
rect 33398 45848 33410 45850
rect 33586 45848 33598 45882
rect 33398 45842 33598 45848
rect 33630 45850 33710 45870
rect 32862 45804 32870 45838
rect 32860 45790 32870 45804
rect 32790 45770 32870 45790
rect 32900 45794 33100 45800
rect 32900 45760 32912 45794
rect 33088 45790 33100 45794
rect 33398 45794 33598 45800
rect 33398 45790 33410 45794
rect 33088 45760 33410 45790
rect 33586 45760 33598 45794
rect 33630 45790 33640 45850
rect 33700 45790 33710 45850
rect 33630 45770 33710 45790
rect 32900 45754 33100 45760
rect 32680 45630 32750 45690
rect 32680 45390 32700 45630
rect 32740 45390 32750 45630
rect 33210 45750 33290 45760
rect 33398 45754 33598 45760
rect 33210 45690 33220 45750
rect 33280 45690 33290 45750
rect 33210 45640 33290 45690
rect 33210 45580 33220 45640
rect 33280 45580 33290 45640
rect 32900 45572 33100 45578
rect 32790 45540 32870 45560
rect 32790 45480 32800 45540
rect 32860 45528 32870 45540
rect 32900 45538 32912 45572
rect 33088 45570 33100 45572
rect 33210 45570 33290 45580
rect 33760 45710 33770 45950
rect 33810 45710 33830 45950
rect 33760 45630 33830 45710
rect 33398 45572 33598 45578
rect 33398 45570 33410 45572
rect 33088 45540 33410 45570
rect 33088 45538 33100 45540
rect 32900 45532 33100 45538
rect 33398 45538 33410 45540
rect 33586 45538 33598 45572
rect 33398 45532 33598 45538
rect 33630 45540 33710 45560
rect 32862 45494 32870 45528
rect 32860 45480 32870 45494
rect 32790 45460 32870 45480
rect 32900 45484 33100 45490
rect 32900 45450 32912 45484
rect 33088 45480 33100 45484
rect 33398 45484 33598 45490
rect 33398 45480 33410 45484
rect 33088 45470 33410 45480
rect 33088 45450 33220 45470
rect 32900 45444 33100 45450
rect 33210 45410 33220 45450
rect 33280 45450 33410 45470
rect 33586 45450 33598 45484
rect 33630 45480 33640 45540
rect 33700 45480 33710 45540
rect 33630 45460 33710 45480
rect 33280 45410 33290 45450
rect 33398 45444 33598 45450
rect 33210 45400 33290 45410
rect 32680 44240 32750 45390
rect 32680 43980 32700 44240
rect 32740 43980 32750 44240
rect 33760 45390 33770 45630
rect 33810 45390 33830 45630
rect 33760 44240 33830 45390
rect 33210 44210 33290 44220
rect 32900 44172 33100 44178
rect 32790 44140 32870 44160
rect 32790 44080 32800 44140
rect 32860 44128 32870 44140
rect 32900 44138 32912 44172
rect 33088 44170 33100 44172
rect 33210 44170 33220 44210
rect 33088 44150 33220 44170
rect 33280 44170 33290 44210
rect 33398 44172 33598 44178
rect 33398 44170 33410 44172
rect 33280 44150 33410 44170
rect 33088 44140 33410 44150
rect 33088 44138 33100 44140
rect 32900 44132 33100 44138
rect 33398 44138 33410 44140
rect 33586 44138 33598 44172
rect 33398 44132 33598 44138
rect 33630 44140 33710 44160
rect 32862 44094 32870 44128
rect 32860 44080 32870 44094
rect 32790 44060 32870 44080
rect 32900 44084 33100 44090
rect 32900 44050 32912 44084
rect 33088 44080 33100 44084
rect 33398 44084 33598 44090
rect 33398 44080 33410 44084
rect 33088 44050 33410 44080
rect 33586 44050 33598 44084
rect 33630 44080 33640 44140
rect 33700 44080 33710 44140
rect 33630 44060 33710 44080
rect 32900 44044 33100 44050
rect 32680 43920 32750 43980
rect 32680 43680 32700 43920
rect 32740 43680 32750 43920
rect 33210 44040 33290 44050
rect 33398 44044 33598 44050
rect 33210 43980 33220 44040
rect 33280 43980 33290 44040
rect 33210 43930 33290 43980
rect 33210 43870 33220 43930
rect 33280 43870 33290 43930
rect 32900 43862 33100 43868
rect 32790 43830 32870 43850
rect 32790 43770 32800 43830
rect 32860 43818 32870 43830
rect 32900 43828 32912 43862
rect 33088 43860 33100 43862
rect 33210 43860 33290 43870
rect 33760 44000 33770 44240
rect 33810 44000 33830 44240
rect 33760 43920 33830 44000
rect 33398 43862 33598 43868
rect 33398 43860 33410 43862
rect 33088 43830 33410 43860
rect 33088 43828 33100 43830
rect 32900 43822 33100 43828
rect 33398 43828 33410 43830
rect 33586 43828 33598 43862
rect 33398 43822 33598 43828
rect 33630 43830 33710 43850
rect 32862 43784 32870 43818
rect 32860 43770 32870 43784
rect 32790 43750 32870 43770
rect 32900 43774 33100 43780
rect 32900 43740 32912 43774
rect 33088 43770 33100 43774
rect 33398 43774 33598 43780
rect 33398 43770 33410 43774
rect 33088 43760 33410 43770
rect 33088 43740 33220 43760
rect 32900 43734 33100 43740
rect 33210 43700 33220 43740
rect 33280 43740 33410 43760
rect 33586 43740 33598 43774
rect 33630 43770 33640 43830
rect 33700 43770 33710 43830
rect 33630 43750 33710 43770
rect 33280 43700 33290 43740
rect 33398 43734 33598 43740
rect 33210 43690 33290 43700
rect 32680 42530 32750 43680
rect 32680 42270 32700 42530
rect 32740 42270 32750 42530
rect 33760 43680 33770 43920
rect 33810 43680 33830 43920
rect 33760 42530 33830 43680
rect 33210 42500 33290 42510
rect 32900 42462 33100 42468
rect 32790 42430 32870 42450
rect 32790 42370 32800 42430
rect 32860 42418 32870 42430
rect 32900 42428 32912 42462
rect 33088 42460 33100 42462
rect 33210 42460 33220 42500
rect 33088 42440 33220 42460
rect 33280 42460 33290 42500
rect 33398 42462 33598 42468
rect 33398 42460 33410 42462
rect 33280 42440 33410 42460
rect 33088 42430 33410 42440
rect 33088 42428 33100 42430
rect 32900 42422 33100 42428
rect 33398 42428 33410 42430
rect 33586 42428 33598 42462
rect 33398 42422 33598 42428
rect 33630 42430 33710 42450
rect 32862 42384 32870 42418
rect 32860 42370 32870 42384
rect 32790 42350 32870 42370
rect 32900 42374 33100 42380
rect 32900 42340 32912 42374
rect 33088 42370 33100 42374
rect 33398 42374 33598 42380
rect 33398 42370 33410 42374
rect 33088 42340 33410 42370
rect 33586 42340 33598 42374
rect 33630 42370 33640 42430
rect 33700 42370 33710 42430
rect 33630 42350 33710 42370
rect 32900 42334 33100 42340
rect 32680 42210 32750 42270
rect 32680 41970 32700 42210
rect 32740 41970 32750 42210
rect 33210 42330 33290 42340
rect 33398 42334 33598 42340
rect 33210 42270 33220 42330
rect 33280 42270 33290 42330
rect 33210 42220 33290 42270
rect 33210 42160 33220 42220
rect 33280 42160 33290 42220
rect 32900 42152 33100 42158
rect 32790 42120 32870 42140
rect 32790 42060 32800 42120
rect 32860 42108 32870 42120
rect 32900 42118 32912 42152
rect 33088 42150 33100 42152
rect 33210 42150 33290 42160
rect 33760 42290 33770 42530
rect 33810 42290 33830 42530
rect 33760 42210 33830 42290
rect 33398 42152 33598 42158
rect 33398 42150 33410 42152
rect 33088 42120 33410 42150
rect 33088 42118 33100 42120
rect 32900 42112 33100 42118
rect 33398 42118 33410 42120
rect 33586 42118 33598 42152
rect 33398 42112 33598 42118
rect 33630 42120 33710 42140
rect 32862 42074 32870 42108
rect 32860 42060 32870 42074
rect 32790 42040 32870 42060
rect 32900 42064 33100 42070
rect 32900 42030 32912 42064
rect 33088 42060 33100 42064
rect 33398 42064 33598 42070
rect 33398 42060 33410 42064
rect 33088 42050 33410 42060
rect 33088 42030 33220 42050
rect 32900 42024 33100 42030
rect 33210 41990 33220 42030
rect 33280 42030 33410 42050
rect 33586 42030 33598 42064
rect 33630 42060 33640 42120
rect 33700 42060 33710 42120
rect 33630 42040 33710 42060
rect 33280 41990 33290 42030
rect 33398 42024 33598 42030
rect 33210 41980 33290 41990
rect 32680 40820 32750 41970
rect 32680 40560 32700 40820
rect 32740 40560 32750 40820
rect 33760 41970 33770 42210
rect 33810 41970 33830 42210
rect 33760 40820 33830 41970
rect 33210 40790 33290 40800
rect 32900 40752 33100 40758
rect 32790 40720 32870 40740
rect 32790 40660 32800 40720
rect 32860 40708 32870 40720
rect 32900 40718 32912 40752
rect 33088 40750 33100 40752
rect 33210 40750 33220 40790
rect 33088 40730 33220 40750
rect 33280 40750 33290 40790
rect 33398 40752 33598 40758
rect 33398 40750 33410 40752
rect 33280 40730 33410 40750
rect 33088 40720 33410 40730
rect 33088 40718 33100 40720
rect 32900 40712 33100 40718
rect 33398 40718 33410 40720
rect 33586 40718 33598 40752
rect 33398 40712 33598 40718
rect 33630 40720 33710 40740
rect 32862 40674 32870 40708
rect 32860 40660 32870 40674
rect 32790 40640 32870 40660
rect 32900 40664 33100 40670
rect 32900 40630 32912 40664
rect 33088 40660 33100 40664
rect 33398 40664 33598 40670
rect 33398 40660 33410 40664
rect 33088 40630 33410 40660
rect 33586 40630 33598 40664
rect 33630 40660 33640 40720
rect 33700 40660 33710 40720
rect 33630 40640 33710 40660
rect 32900 40624 33100 40630
rect 32680 40500 32750 40560
rect 32680 40260 32700 40500
rect 32740 40260 32750 40500
rect 33210 40620 33290 40630
rect 33398 40624 33598 40630
rect 33210 40560 33220 40620
rect 33280 40560 33290 40620
rect 33210 40510 33290 40560
rect 33210 40450 33220 40510
rect 33280 40450 33290 40510
rect 32900 40442 33100 40448
rect 32790 40410 32870 40430
rect 32790 40350 32800 40410
rect 32860 40398 32870 40410
rect 32900 40408 32912 40442
rect 33088 40440 33100 40442
rect 33210 40440 33290 40450
rect 33760 40580 33770 40820
rect 33810 40580 33830 40820
rect 33760 40500 33830 40580
rect 33398 40442 33598 40448
rect 33398 40440 33410 40442
rect 33088 40410 33410 40440
rect 33088 40408 33100 40410
rect 32900 40402 33100 40408
rect 33398 40408 33410 40410
rect 33586 40408 33598 40442
rect 33398 40402 33598 40408
rect 33630 40410 33710 40430
rect 32862 40364 32870 40398
rect 32860 40350 32870 40364
rect 32790 40330 32870 40350
rect 32900 40354 33100 40360
rect 32900 40320 32912 40354
rect 33088 40350 33100 40354
rect 33398 40354 33598 40360
rect 33398 40350 33410 40354
rect 33088 40340 33410 40350
rect 33088 40320 33220 40340
rect 32900 40314 33100 40320
rect 33210 40280 33220 40320
rect 33280 40320 33410 40340
rect 33586 40320 33598 40354
rect 33630 40350 33640 40410
rect 33700 40350 33710 40410
rect 33630 40330 33710 40350
rect 33280 40280 33290 40320
rect 33398 40314 33598 40320
rect 33210 40270 33290 40280
rect 32680 39690 32750 40260
rect 33760 40260 33770 40500
rect 33810 40260 33830 40500
rect 33760 39690 33830 40260
rect 32680 39680 32760 39690
rect 32680 39620 32690 39680
rect 32750 39620 32760 39680
rect 33750 39680 33830 39690
rect 33750 39620 33760 39680
rect 33820 39620 33830 39680
rect 33750 39610 33830 39620
rect 33860 66480 33890 67050
rect 33860 66470 33920 66480
rect 33860 66400 33920 66410
rect 33860 64770 33890 66400
rect 33950 65950 33980 67050
rect 33920 65940 33980 65950
rect 33920 65870 33980 65880
rect 33860 64760 33920 64770
rect 33860 64690 33920 64700
rect 33860 63060 33890 64690
rect 33950 64240 33980 65870
rect 33920 64230 33980 64240
rect 33920 64160 33980 64170
rect 33860 63050 33920 63060
rect 33860 62980 33920 62990
rect 33860 61350 33890 62980
rect 33950 62530 33980 64160
rect 33920 62520 33980 62530
rect 33920 62450 33980 62460
rect 33860 61340 33920 61350
rect 33860 61270 33920 61280
rect 33860 59640 33890 61270
rect 33950 60820 33980 62450
rect 33920 60810 33980 60820
rect 33920 60740 33980 60750
rect 33860 59630 33920 59640
rect 33860 59560 33920 59570
rect 33860 57930 33890 59560
rect 33950 59110 33980 60740
rect 33920 59100 33980 59110
rect 33920 59030 33980 59040
rect 33860 57920 33920 57930
rect 33860 57850 33920 57860
rect 33860 56220 33890 57850
rect 33950 57400 33980 59030
rect 33920 57390 33980 57400
rect 33920 57320 33980 57330
rect 33860 56210 33920 56220
rect 33860 56140 33920 56150
rect 33860 54510 33890 56140
rect 33950 55690 33980 57320
rect 33920 55680 33980 55690
rect 33920 55610 33980 55620
rect 33860 54500 33920 54510
rect 33860 54430 33920 54440
rect 33860 52800 33890 54430
rect 33950 53980 33980 55610
rect 33920 53970 33980 53980
rect 33920 53900 33980 53910
rect 33860 52790 33920 52800
rect 33860 52720 33920 52730
rect 33860 51090 33890 52720
rect 33950 52270 33980 53900
rect 33920 52260 33980 52270
rect 33920 52190 33980 52200
rect 33860 51080 33920 51090
rect 33860 51010 33920 51020
rect 33860 49380 33890 51010
rect 33950 50560 33980 52190
rect 33920 50550 33980 50560
rect 33920 50480 33980 50490
rect 33860 49370 33920 49380
rect 33860 49300 33920 49310
rect 33860 47670 33890 49300
rect 33950 48850 33980 50480
rect 33920 48840 33980 48850
rect 33920 48770 33980 48780
rect 33860 47660 33920 47670
rect 33860 47590 33920 47600
rect 33860 45960 33890 47590
rect 33950 47140 33980 48770
rect 33920 47130 33980 47140
rect 33920 47060 33980 47070
rect 33860 45950 33920 45960
rect 33860 45880 33920 45890
rect 33860 44250 33890 45880
rect 33950 45430 33980 47060
rect 33920 45420 33980 45430
rect 33920 45350 33980 45360
rect 33860 44240 33920 44250
rect 33860 44170 33920 44180
rect 33860 42540 33890 44170
rect 33950 43720 33980 45350
rect 33920 43710 33980 43720
rect 33920 43640 33980 43650
rect 33860 42530 33920 42540
rect 33860 42460 33920 42470
rect 33860 40830 33890 42460
rect 33950 42010 33980 43640
rect 33920 42000 33980 42010
rect 33920 41930 33980 41940
rect 33860 40820 33920 40830
rect 33860 40750 33920 40760
rect 32210 39220 32270 39230
rect 32390 39230 32650 39240
rect 29220 39160 29280 39170
rect 32450 39210 32650 39230
rect 32390 39160 32450 39170
rect 33860 38840 33890 40750
rect 33950 40300 33980 41930
rect 33920 40290 33980 40300
rect 33920 40220 33980 40230
rect 33950 39690 33980 40220
rect 33920 39680 33980 39690
rect 33920 39610 33980 39620
rect 34010 66390 34040 67050
rect 34010 66380 34070 66390
rect 34010 66310 34070 66320
rect 34010 64680 34040 66310
rect 34010 64670 34070 64680
rect 34010 64600 34070 64610
rect 34010 42450 34040 64600
rect 34130 62970 34160 67050
rect 34130 62960 34190 62970
rect 34130 62890 34190 62900
rect 34130 61260 34160 62890
rect 34130 61250 34190 61260
rect 34130 61180 34190 61190
rect 34130 45870 34160 61180
rect 34250 59550 34280 67050
rect 34250 59540 34310 59550
rect 34250 59470 34310 59480
rect 34250 47580 34280 59470
rect 34370 57840 34400 67050
rect 34370 57830 34430 57840
rect 34370 57760 34430 57770
rect 34370 49290 34400 57760
rect 34490 56130 34520 67050
rect 34490 56120 34550 56130
rect 34490 56050 34550 56060
rect 34490 51000 34520 56050
rect 34610 54420 34640 67050
rect 34610 54410 34670 54420
rect 34610 54340 34670 54350
rect 34610 52710 34640 54340
rect 34610 52700 34670 52710
rect 34610 52630 34670 52640
rect 34490 50990 34550 51000
rect 34490 50920 34550 50930
rect 34370 49280 34430 49290
rect 34370 49210 34430 49220
rect 34250 47570 34310 47580
rect 34250 47500 34310 47510
rect 34130 45860 34190 45870
rect 34130 45790 34190 45800
rect 34130 44160 34160 45790
rect 34130 44150 34190 44160
rect 34130 44080 34190 44090
rect 34010 42440 34070 42450
rect 34010 42370 34070 42380
rect 34010 40740 34040 42370
rect 34010 40730 34070 40740
rect 34010 40660 34070 40670
rect 34010 39240 34040 40660
rect 34130 39300 34160 44080
rect 34250 39360 34280 47500
rect 34370 39420 34400 49210
rect 34490 39480 34520 50920
rect 34610 39540 34640 52630
rect 34730 39690 34760 67050
rect 36890 54410 36920 67050
rect 36860 54400 36920 54410
rect 36860 54330 36920 54340
rect 36890 39600 36920 54330
rect 37010 52710 37040 67050
rect 37130 56130 37160 67050
rect 37250 57840 37280 67050
rect 37370 59550 37400 67050
rect 37490 62970 37520 67050
rect 37610 66390 37640 67050
rect 37580 66380 37640 66390
rect 37580 66310 37640 66320
rect 37610 64680 37640 66310
rect 37580 64670 37640 64680
rect 37580 64600 37640 64610
rect 37460 62960 37520 62970
rect 37460 62890 37520 62900
rect 37490 61260 37520 62890
rect 37460 61250 37520 61260
rect 37460 61180 37520 61190
rect 37340 59540 37400 59550
rect 37340 59470 37400 59480
rect 37220 57830 37280 57840
rect 37220 57760 37280 57770
rect 37100 56120 37160 56130
rect 37100 56050 37160 56060
rect 36980 52700 37040 52710
rect 36980 52630 37040 52640
rect 36300 39590 36920 39600
rect 34610 39530 35170 39540
rect 34610 39510 35110 39530
rect 34490 39470 34990 39480
rect 34490 39450 34930 39470
rect 34370 39410 34810 39420
rect 34370 39390 34750 39410
rect 34250 39350 34630 39360
rect 34250 39330 34570 39350
rect 34130 39290 34450 39300
rect 34130 39270 34390 39290
rect 34010 39230 34270 39240
rect 34010 39210 34210 39230
rect 36360 39570 36920 39590
rect 37010 39540 37040 52630
rect 37130 51000 37160 56050
rect 37100 50990 37160 51000
rect 37100 50920 37160 50930
rect 36300 39520 36360 39530
rect 36480 39530 37040 39540
rect 35110 39460 35170 39470
rect 36540 39510 37040 39530
rect 37130 39480 37160 50920
rect 37250 49290 37280 57760
rect 37220 49280 37280 49290
rect 37220 49210 37280 49220
rect 36480 39460 36540 39470
rect 36660 39470 37160 39480
rect 34930 39400 34990 39410
rect 36720 39450 37160 39470
rect 37250 39420 37280 49210
rect 37370 47580 37400 59470
rect 37340 47570 37400 47580
rect 37340 47500 37400 47510
rect 36660 39400 36720 39410
rect 36840 39410 37280 39420
rect 34750 39340 34810 39350
rect 36900 39390 37280 39410
rect 37370 39360 37400 47500
rect 37490 45870 37520 61180
rect 37460 45860 37520 45870
rect 37460 45790 37520 45800
rect 37490 44160 37520 45790
rect 37460 44150 37520 44160
rect 37460 44080 37520 44090
rect 36840 39340 36900 39350
rect 37020 39350 37400 39360
rect 34570 39280 34630 39290
rect 37080 39330 37400 39350
rect 37490 39300 37520 44080
rect 37610 42450 37640 64600
rect 37580 42440 37640 42450
rect 37580 42370 37640 42380
rect 37610 40740 37640 42370
rect 37580 40730 37640 40740
rect 37580 40660 37640 40670
rect 37020 39280 37080 39290
rect 37200 39290 37520 39300
rect 34390 39220 34450 39230
rect 37260 39270 37520 39290
rect 37610 39240 37640 40660
rect 37670 66470 37740 67050
rect 37670 66210 37690 66470
rect 37730 66210 37740 66470
rect 38750 66470 38820 67050
rect 38200 66440 38280 66450
rect 37890 66402 38090 66408
rect 37780 66370 37860 66390
rect 37780 66310 37790 66370
rect 37850 66358 37860 66370
rect 37890 66368 37902 66402
rect 38078 66400 38090 66402
rect 38200 66400 38210 66440
rect 38078 66380 38210 66400
rect 38270 66400 38280 66440
rect 38388 66402 38588 66408
rect 38388 66400 38400 66402
rect 38270 66380 38400 66400
rect 38078 66370 38400 66380
rect 38078 66368 38090 66370
rect 37890 66362 38090 66368
rect 38388 66368 38400 66370
rect 38576 66368 38588 66402
rect 38388 66362 38588 66368
rect 38620 66370 38700 66390
rect 37852 66324 37860 66358
rect 37850 66310 37860 66324
rect 37780 66290 37860 66310
rect 37890 66314 38090 66320
rect 37890 66280 37902 66314
rect 38078 66310 38090 66314
rect 38388 66314 38588 66320
rect 38388 66310 38400 66314
rect 38078 66280 38400 66310
rect 38576 66280 38588 66314
rect 38620 66310 38630 66370
rect 38690 66310 38700 66370
rect 38620 66290 38700 66310
rect 37890 66274 38090 66280
rect 37670 66150 37740 66210
rect 37670 65910 37690 66150
rect 37730 65910 37740 66150
rect 38200 66270 38280 66280
rect 38388 66274 38588 66280
rect 38200 66210 38210 66270
rect 38270 66210 38280 66270
rect 38200 66160 38280 66210
rect 38200 66100 38210 66160
rect 38270 66100 38280 66160
rect 37890 66092 38090 66098
rect 37780 66060 37860 66080
rect 37780 66000 37790 66060
rect 37850 66048 37860 66060
rect 37890 66058 37902 66092
rect 38078 66090 38090 66092
rect 38200 66090 38280 66100
rect 38750 66230 38760 66470
rect 38800 66230 38820 66470
rect 38750 66150 38820 66230
rect 38388 66092 38588 66098
rect 38388 66090 38400 66092
rect 38078 66060 38400 66090
rect 38078 66058 38090 66060
rect 37890 66052 38090 66058
rect 38388 66058 38400 66060
rect 38576 66058 38588 66092
rect 38388 66052 38588 66058
rect 38620 66060 38700 66080
rect 37852 66014 37860 66048
rect 37850 66000 37860 66014
rect 37780 65980 37860 66000
rect 37890 66004 38090 66010
rect 37890 65970 37902 66004
rect 38078 66000 38090 66004
rect 38388 66004 38588 66010
rect 38388 66000 38400 66004
rect 38078 65990 38400 66000
rect 38078 65970 38210 65990
rect 37890 65964 38090 65970
rect 38200 65930 38210 65970
rect 38270 65970 38400 65990
rect 38576 65970 38588 66004
rect 38620 66000 38630 66060
rect 38690 66000 38700 66060
rect 38620 65980 38700 66000
rect 38270 65930 38280 65970
rect 38388 65964 38588 65970
rect 38200 65920 38280 65930
rect 37670 64760 37740 65910
rect 37670 64500 37690 64760
rect 37730 64500 37740 64760
rect 38750 65910 38760 66150
rect 38800 65910 38820 66150
rect 38750 64760 38820 65910
rect 38200 64730 38280 64740
rect 37890 64692 38090 64698
rect 37780 64660 37860 64680
rect 37780 64600 37790 64660
rect 37850 64648 37860 64660
rect 37890 64658 37902 64692
rect 38078 64690 38090 64692
rect 38200 64690 38210 64730
rect 38078 64670 38210 64690
rect 38270 64690 38280 64730
rect 38388 64692 38588 64698
rect 38388 64690 38400 64692
rect 38270 64670 38400 64690
rect 38078 64660 38400 64670
rect 38078 64658 38090 64660
rect 37890 64652 38090 64658
rect 38388 64658 38400 64660
rect 38576 64658 38588 64692
rect 38388 64652 38588 64658
rect 38620 64660 38700 64680
rect 37852 64614 37860 64648
rect 37850 64600 37860 64614
rect 37780 64580 37860 64600
rect 37890 64604 38090 64610
rect 37890 64570 37902 64604
rect 38078 64600 38090 64604
rect 38388 64604 38588 64610
rect 38388 64600 38400 64604
rect 38078 64570 38400 64600
rect 38576 64570 38588 64604
rect 38620 64600 38630 64660
rect 38690 64600 38700 64660
rect 38620 64580 38700 64600
rect 37890 64564 38090 64570
rect 37670 64440 37740 64500
rect 37670 64200 37690 64440
rect 37730 64200 37740 64440
rect 38200 64560 38280 64570
rect 38388 64564 38588 64570
rect 38200 64500 38210 64560
rect 38270 64500 38280 64560
rect 38200 64450 38280 64500
rect 38200 64390 38210 64450
rect 38270 64390 38280 64450
rect 37890 64382 38090 64388
rect 37780 64350 37860 64370
rect 37780 64290 37790 64350
rect 37850 64338 37860 64350
rect 37890 64348 37902 64382
rect 38078 64380 38090 64382
rect 38200 64380 38280 64390
rect 38750 64520 38760 64760
rect 38800 64520 38820 64760
rect 38750 64440 38820 64520
rect 38388 64382 38588 64388
rect 38388 64380 38400 64382
rect 38078 64350 38400 64380
rect 38078 64348 38090 64350
rect 37890 64342 38090 64348
rect 38388 64348 38400 64350
rect 38576 64348 38588 64382
rect 38388 64342 38588 64348
rect 38620 64350 38700 64370
rect 37852 64304 37860 64338
rect 37850 64290 37860 64304
rect 37780 64270 37860 64290
rect 37890 64294 38090 64300
rect 37890 64260 37902 64294
rect 38078 64290 38090 64294
rect 38388 64294 38588 64300
rect 38388 64290 38400 64294
rect 38078 64280 38400 64290
rect 38078 64260 38210 64280
rect 37890 64254 38090 64260
rect 38200 64220 38210 64260
rect 38270 64260 38400 64280
rect 38576 64260 38588 64294
rect 38620 64290 38630 64350
rect 38690 64290 38700 64350
rect 38620 64270 38700 64290
rect 38270 64220 38280 64260
rect 38388 64254 38588 64260
rect 38200 64210 38280 64220
rect 37670 63050 37740 64200
rect 37670 62790 37690 63050
rect 37730 62790 37740 63050
rect 38750 64200 38760 64440
rect 38800 64200 38820 64440
rect 38750 63050 38820 64200
rect 38200 63020 38280 63030
rect 37890 62982 38090 62988
rect 37780 62950 37860 62970
rect 37780 62890 37790 62950
rect 37850 62938 37860 62950
rect 37890 62948 37902 62982
rect 38078 62980 38090 62982
rect 38200 62980 38210 63020
rect 38078 62960 38210 62980
rect 38270 62980 38280 63020
rect 38388 62982 38588 62988
rect 38388 62980 38400 62982
rect 38270 62960 38400 62980
rect 38078 62950 38400 62960
rect 38078 62948 38090 62950
rect 37890 62942 38090 62948
rect 38388 62948 38400 62950
rect 38576 62948 38588 62982
rect 38388 62942 38588 62948
rect 38620 62950 38700 62970
rect 37852 62904 37860 62938
rect 37850 62890 37860 62904
rect 37780 62870 37860 62890
rect 37890 62894 38090 62900
rect 37890 62860 37902 62894
rect 38078 62890 38090 62894
rect 38388 62894 38588 62900
rect 38388 62890 38400 62894
rect 38078 62860 38400 62890
rect 38576 62860 38588 62894
rect 38620 62890 38630 62950
rect 38690 62890 38700 62950
rect 38620 62870 38700 62890
rect 37890 62854 38090 62860
rect 37670 62730 37740 62790
rect 37670 62490 37690 62730
rect 37730 62490 37740 62730
rect 38200 62850 38280 62860
rect 38388 62854 38588 62860
rect 38200 62790 38210 62850
rect 38270 62790 38280 62850
rect 38200 62740 38280 62790
rect 38200 62680 38210 62740
rect 38270 62680 38280 62740
rect 37890 62672 38090 62678
rect 37780 62640 37860 62660
rect 37780 62580 37790 62640
rect 37850 62628 37860 62640
rect 37890 62638 37902 62672
rect 38078 62670 38090 62672
rect 38200 62670 38280 62680
rect 38750 62810 38760 63050
rect 38800 62810 38820 63050
rect 38750 62730 38820 62810
rect 38388 62672 38588 62678
rect 38388 62670 38400 62672
rect 38078 62640 38400 62670
rect 38078 62638 38090 62640
rect 37890 62632 38090 62638
rect 38388 62638 38400 62640
rect 38576 62638 38588 62672
rect 38388 62632 38588 62638
rect 38620 62640 38700 62660
rect 37852 62594 37860 62628
rect 37850 62580 37860 62594
rect 37780 62560 37860 62580
rect 37890 62584 38090 62590
rect 37890 62550 37902 62584
rect 38078 62580 38090 62584
rect 38388 62584 38588 62590
rect 38388 62580 38400 62584
rect 38078 62570 38400 62580
rect 38078 62550 38210 62570
rect 37890 62544 38090 62550
rect 38200 62510 38210 62550
rect 38270 62550 38400 62570
rect 38576 62550 38588 62584
rect 38620 62580 38630 62640
rect 38690 62580 38700 62640
rect 38620 62560 38700 62580
rect 38270 62510 38280 62550
rect 38388 62544 38588 62550
rect 38200 62500 38280 62510
rect 37670 61340 37740 62490
rect 37670 61080 37690 61340
rect 37730 61080 37740 61340
rect 38750 62490 38760 62730
rect 38800 62490 38820 62730
rect 38750 61340 38820 62490
rect 38200 61310 38280 61320
rect 37890 61272 38090 61278
rect 37780 61240 37860 61260
rect 37780 61180 37790 61240
rect 37850 61228 37860 61240
rect 37890 61238 37902 61272
rect 38078 61270 38090 61272
rect 38200 61270 38210 61310
rect 38078 61250 38210 61270
rect 38270 61270 38280 61310
rect 38388 61272 38588 61278
rect 38388 61270 38400 61272
rect 38270 61250 38400 61270
rect 38078 61240 38400 61250
rect 38078 61238 38090 61240
rect 37890 61232 38090 61238
rect 38388 61238 38400 61240
rect 38576 61238 38588 61272
rect 38388 61232 38588 61238
rect 38620 61240 38700 61260
rect 37852 61194 37860 61228
rect 37850 61180 37860 61194
rect 37780 61160 37860 61180
rect 37890 61184 38090 61190
rect 37890 61150 37902 61184
rect 38078 61180 38090 61184
rect 38388 61184 38588 61190
rect 38388 61180 38400 61184
rect 38078 61150 38400 61180
rect 38576 61150 38588 61184
rect 38620 61180 38630 61240
rect 38690 61180 38700 61240
rect 38620 61160 38700 61180
rect 37890 61144 38090 61150
rect 37670 61020 37740 61080
rect 37670 60780 37690 61020
rect 37730 60780 37740 61020
rect 38200 61140 38280 61150
rect 38388 61144 38588 61150
rect 38200 61080 38210 61140
rect 38270 61080 38280 61140
rect 38200 61030 38280 61080
rect 38200 60970 38210 61030
rect 38270 60970 38280 61030
rect 37890 60962 38090 60968
rect 37780 60930 37860 60950
rect 37780 60870 37790 60930
rect 37850 60918 37860 60930
rect 37890 60928 37902 60962
rect 38078 60960 38090 60962
rect 38200 60960 38280 60970
rect 38750 61100 38760 61340
rect 38800 61100 38820 61340
rect 38750 61020 38820 61100
rect 38388 60962 38588 60968
rect 38388 60960 38400 60962
rect 38078 60930 38400 60960
rect 38078 60928 38090 60930
rect 37890 60922 38090 60928
rect 38388 60928 38400 60930
rect 38576 60928 38588 60962
rect 38388 60922 38588 60928
rect 38620 60930 38700 60950
rect 37852 60884 37860 60918
rect 37850 60870 37860 60884
rect 37780 60850 37860 60870
rect 37890 60874 38090 60880
rect 37890 60840 37902 60874
rect 38078 60870 38090 60874
rect 38388 60874 38588 60880
rect 38388 60870 38400 60874
rect 38078 60860 38400 60870
rect 38078 60840 38210 60860
rect 37890 60834 38090 60840
rect 38200 60800 38210 60840
rect 38270 60840 38400 60860
rect 38576 60840 38588 60874
rect 38620 60870 38630 60930
rect 38690 60870 38700 60930
rect 38620 60850 38700 60870
rect 38270 60800 38280 60840
rect 38388 60834 38588 60840
rect 38200 60790 38280 60800
rect 37670 59630 37740 60780
rect 37670 59370 37690 59630
rect 37730 59370 37740 59630
rect 38750 60780 38760 61020
rect 38800 60780 38820 61020
rect 38750 59630 38820 60780
rect 38200 59600 38280 59610
rect 37890 59562 38090 59568
rect 37780 59530 37860 59550
rect 37780 59470 37790 59530
rect 37850 59518 37860 59530
rect 37890 59528 37902 59562
rect 38078 59560 38090 59562
rect 38200 59560 38210 59600
rect 38078 59540 38210 59560
rect 38270 59560 38280 59600
rect 38388 59562 38588 59568
rect 38388 59560 38400 59562
rect 38270 59540 38400 59560
rect 38078 59530 38400 59540
rect 38078 59528 38090 59530
rect 37890 59522 38090 59528
rect 38388 59528 38400 59530
rect 38576 59528 38588 59562
rect 38388 59522 38588 59528
rect 38620 59530 38700 59550
rect 37852 59484 37860 59518
rect 37850 59470 37860 59484
rect 37780 59450 37860 59470
rect 37890 59474 38090 59480
rect 37890 59440 37902 59474
rect 38078 59470 38090 59474
rect 38388 59474 38588 59480
rect 38388 59470 38400 59474
rect 38078 59440 38400 59470
rect 38576 59440 38588 59474
rect 38620 59470 38630 59530
rect 38690 59470 38700 59530
rect 38620 59450 38700 59470
rect 37890 59434 38090 59440
rect 37670 59310 37740 59370
rect 37670 59070 37690 59310
rect 37730 59070 37740 59310
rect 38200 59430 38280 59440
rect 38388 59434 38588 59440
rect 38200 59370 38210 59430
rect 38270 59370 38280 59430
rect 38200 59320 38280 59370
rect 38200 59260 38210 59320
rect 38270 59260 38280 59320
rect 37890 59252 38090 59258
rect 37780 59220 37860 59240
rect 37780 59160 37790 59220
rect 37850 59208 37860 59220
rect 37890 59218 37902 59252
rect 38078 59250 38090 59252
rect 38200 59250 38280 59260
rect 38750 59390 38760 59630
rect 38800 59390 38820 59630
rect 38750 59310 38820 59390
rect 38388 59252 38588 59258
rect 38388 59250 38400 59252
rect 38078 59220 38400 59250
rect 38078 59218 38090 59220
rect 37890 59212 38090 59218
rect 38388 59218 38400 59220
rect 38576 59218 38588 59252
rect 38388 59212 38588 59218
rect 38620 59220 38700 59240
rect 37852 59174 37860 59208
rect 37850 59160 37860 59174
rect 37780 59140 37860 59160
rect 37890 59164 38090 59170
rect 37890 59130 37902 59164
rect 38078 59160 38090 59164
rect 38388 59164 38588 59170
rect 38388 59160 38400 59164
rect 38078 59150 38400 59160
rect 38078 59130 38210 59150
rect 37890 59124 38090 59130
rect 38200 59090 38210 59130
rect 38270 59130 38400 59150
rect 38576 59130 38588 59164
rect 38620 59160 38630 59220
rect 38690 59160 38700 59220
rect 38620 59140 38700 59160
rect 38270 59090 38280 59130
rect 38388 59124 38588 59130
rect 38200 59080 38280 59090
rect 37670 57920 37740 59070
rect 37670 57660 37690 57920
rect 37730 57660 37740 57920
rect 38750 59070 38760 59310
rect 38800 59070 38820 59310
rect 38750 57920 38820 59070
rect 38200 57890 38280 57900
rect 37890 57852 38090 57858
rect 37780 57820 37860 57840
rect 37780 57760 37790 57820
rect 37850 57808 37860 57820
rect 37890 57818 37902 57852
rect 38078 57850 38090 57852
rect 38200 57850 38210 57890
rect 38078 57830 38210 57850
rect 38270 57850 38280 57890
rect 38388 57852 38588 57858
rect 38388 57850 38400 57852
rect 38270 57830 38400 57850
rect 38078 57820 38400 57830
rect 38078 57818 38090 57820
rect 37890 57812 38090 57818
rect 38388 57818 38400 57820
rect 38576 57818 38588 57852
rect 38388 57812 38588 57818
rect 38620 57820 38700 57840
rect 37852 57774 37860 57808
rect 37850 57760 37860 57774
rect 37780 57740 37860 57760
rect 37890 57764 38090 57770
rect 37890 57730 37902 57764
rect 38078 57760 38090 57764
rect 38388 57764 38588 57770
rect 38388 57760 38400 57764
rect 38078 57730 38400 57760
rect 38576 57730 38588 57764
rect 38620 57760 38630 57820
rect 38690 57760 38700 57820
rect 38620 57740 38700 57760
rect 37890 57724 38090 57730
rect 37670 57600 37740 57660
rect 37670 57360 37690 57600
rect 37730 57360 37740 57600
rect 38200 57720 38280 57730
rect 38388 57724 38588 57730
rect 38200 57660 38210 57720
rect 38270 57660 38280 57720
rect 38200 57610 38280 57660
rect 38200 57550 38210 57610
rect 38270 57550 38280 57610
rect 37890 57542 38090 57548
rect 37780 57510 37860 57530
rect 37780 57450 37790 57510
rect 37850 57498 37860 57510
rect 37890 57508 37902 57542
rect 38078 57540 38090 57542
rect 38200 57540 38280 57550
rect 38750 57680 38760 57920
rect 38800 57680 38820 57920
rect 38750 57600 38820 57680
rect 38388 57542 38588 57548
rect 38388 57540 38400 57542
rect 38078 57510 38400 57540
rect 38078 57508 38090 57510
rect 37890 57502 38090 57508
rect 38388 57508 38400 57510
rect 38576 57508 38588 57542
rect 38388 57502 38588 57508
rect 38620 57510 38700 57530
rect 37852 57464 37860 57498
rect 37850 57450 37860 57464
rect 37780 57430 37860 57450
rect 37890 57454 38090 57460
rect 37890 57420 37902 57454
rect 38078 57450 38090 57454
rect 38388 57454 38588 57460
rect 38388 57450 38400 57454
rect 38078 57440 38400 57450
rect 38078 57420 38210 57440
rect 37890 57414 38090 57420
rect 38200 57380 38210 57420
rect 38270 57420 38400 57440
rect 38576 57420 38588 57454
rect 38620 57450 38630 57510
rect 38690 57450 38700 57510
rect 38620 57430 38700 57450
rect 38270 57380 38280 57420
rect 38388 57414 38588 57420
rect 38200 57370 38280 57380
rect 37670 56210 37740 57360
rect 37670 55950 37690 56210
rect 37730 55950 37740 56210
rect 38750 57360 38760 57600
rect 38800 57360 38820 57600
rect 38750 56210 38820 57360
rect 38200 56180 38280 56190
rect 37890 56142 38090 56148
rect 37780 56110 37860 56130
rect 37780 56050 37790 56110
rect 37850 56098 37860 56110
rect 37890 56108 37902 56142
rect 38078 56140 38090 56142
rect 38200 56140 38210 56180
rect 38078 56120 38210 56140
rect 38270 56140 38280 56180
rect 38388 56142 38588 56148
rect 38388 56140 38400 56142
rect 38270 56120 38400 56140
rect 38078 56110 38400 56120
rect 38078 56108 38090 56110
rect 37890 56102 38090 56108
rect 38388 56108 38400 56110
rect 38576 56108 38588 56142
rect 38388 56102 38588 56108
rect 38620 56110 38700 56130
rect 37852 56064 37860 56098
rect 37850 56050 37860 56064
rect 37780 56030 37860 56050
rect 37890 56054 38090 56060
rect 37890 56020 37902 56054
rect 38078 56050 38090 56054
rect 38388 56054 38588 56060
rect 38388 56050 38400 56054
rect 38078 56020 38400 56050
rect 38576 56020 38588 56054
rect 38620 56050 38630 56110
rect 38690 56050 38700 56110
rect 38620 56030 38700 56050
rect 37890 56014 38090 56020
rect 37670 55890 37740 55950
rect 37670 55650 37690 55890
rect 37730 55650 37740 55890
rect 38200 56010 38280 56020
rect 38388 56014 38588 56020
rect 38200 55950 38210 56010
rect 38270 55950 38280 56010
rect 38200 55900 38280 55950
rect 38200 55840 38210 55900
rect 38270 55840 38280 55900
rect 37890 55832 38090 55838
rect 37780 55800 37860 55820
rect 37780 55740 37790 55800
rect 37850 55788 37860 55800
rect 37890 55798 37902 55832
rect 38078 55830 38090 55832
rect 38200 55830 38280 55840
rect 38750 55970 38760 56210
rect 38800 55970 38820 56210
rect 38750 55890 38820 55970
rect 38388 55832 38588 55838
rect 38388 55830 38400 55832
rect 38078 55800 38400 55830
rect 38078 55798 38090 55800
rect 37890 55792 38090 55798
rect 38388 55798 38400 55800
rect 38576 55798 38588 55832
rect 38388 55792 38588 55798
rect 38620 55800 38700 55820
rect 37852 55754 37860 55788
rect 37850 55740 37860 55754
rect 37780 55720 37860 55740
rect 37890 55744 38090 55750
rect 37890 55710 37902 55744
rect 38078 55740 38090 55744
rect 38388 55744 38588 55750
rect 38388 55740 38400 55744
rect 38078 55730 38400 55740
rect 38078 55710 38210 55730
rect 37890 55704 38090 55710
rect 38200 55670 38210 55710
rect 38270 55710 38400 55730
rect 38576 55710 38588 55744
rect 38620 55740 38630 55800
rect 38690 55740 38700 55800
rect 38620 55720 38700 55740
rect 38270 55670 38280 55710
rect 38388 55704 38588 55710
rect 38200 55660 38280 55670
rect 37670 54500 37740 55650
rect 37670 54240 37690 54500
rect 37730 54240 37740 54500
rect 38750 55650 38760 55890
rect 38800 55650 38820 55890
rect 38750 54500 38820 55650
rect 38200 54470 38280 54480
rect 37890 54432 38090 54438
rect 37780 54400 37860 54420
rect 37780 54340 37790 54400
rect 37850 54388 37860 54400
rect 37890 54398 37902 54432
rect 38078 54430 38090 54432
rect 38200 54430 38210 54470
rect 38078 54410 38210 54430
rect 38270 54430 38280 54470
rect 38388 54432 38588 54438
rect 38388 54430 38400 54432
rect 38270 54410 38400 54430
rect 38078 54400 38400 54410
rect 38078 54398 38090 54400
rect 37890 54392 38090 54398
rect 38388 54398 38400 54400
rect 38576 54398 38588 54432
rect 38388 54392 38588 54398
rect 38620 54400 38700 54420
rect 37852 54354 37860 54388
rect 37850 54340 37860 54354
rect 37780 54320 37860 54340
rect 37890 54344 38090 54350
rect 37890 54310 37902 54344
rect 38078 54340 38090 54344
rect 38388 54344 38588 54350
rect 38388 54340 38400 54344
rect 38078 54310 38400 54340
rect 38576 54310 38588 54344
rect 38620 54340 38630 54400
rect 38690 54340 38700 54400
rect 38620 54320 38700 54340
rect 37890 54304 38090 54310
rect 37670 54180 37740 54240
rect 37670 53940 37690 54180
rect 37730 53940 37740 54180
rect 38200 54300 38280 54310
rect 38388 54304 38588 54310
rect 38200 54240 38210 54300
rect 38270 54240 38280 54300
rect 38200 54190 38280 54240
rect 38200 54130 38210 54190
rect 38270 54130 38280 54190
rect 37890 54122 38090 54128
rect 37780 54090 37860 54110
rect 37780 54030 37790 54090
rect 37850 54078 37860 54090
rect 37890 54088 37902 54122
rect 38078 54120 38090 54122
rect 38200 54120 38280 54130
rect 38750 54260 38760 54500
rect 38800 54260 38820 54500
rect 38750 54180 38820 54260
rect 38388 54122 38588 54128
rect 38388 54120 38400 54122
rect 38078 54090 38400 54120
rect 38078 54088 38090 54090
rect 37890 54082 38090 54088
rect 38388 54088 38400 54090
rect 38576 54088 38588 54122
rect 38388 54082 38588 54088
rect 38620 54090 38700 54110
rect 37852 54044 37860 54078
rect 37850 54030 37860 54044
rect 37780 54010 37860 54030
rect 37890 54034 38090 54040
rect 37890 54000 37902 54034
rect 38078 54030 38090 54034
rect 38388 54034 38588 54040
rect 38388 54030 38400 54034
rect 38078 54020 38400 54030
rect 38078 54000 38210 54020
rect 37890 53994 38090 54000
rect 38200 53960 38210 54000
rect 38270 54000 38400 54020
rect 38576 54000 38588 54034
rect 38620 54030 38630 54090
rect 38690 54030 38700 54090
rect 38620 54010 38700 54030
rect 38270 53960 38280 54000
rect 38388 53994 38588 54000
rect 38200 53950 38280 53960
rect 37670 52790 37740 53940
rect 37670 52530 37690 52790
rect 37730 52530 37740 52790
rect 38750 53940 38760 54180
rect 38800 53940 38820 54180
rect 38750 52790 38820 53940
rect 38200 52760 38280 52770
rect 37890 52722 38090 52728
rect 37780 52690 37860 52710
rect 37780 52630 37790 52690
rect 37850 52678 37860 52690
rect 37890 52688 37902 52722
rect 38078 52720 38090 52722
rect 38200 52720 38210 52760
rect 38078 52700 38210 52720
rect 38270 52720 38280 52760
rect 38388 52722 38588 52728
rect 38388 52720 38400 52722
rect 38270 52700 38400 52720
rect 38078 52690 38400 52700
rect 38078 52688 38090 52690
rect 37890 52682 38090 52688
rect 38388 52688 38400 52690
rect 38576 52688 38588 52722
rect 38388 52682 38588 52688
rect 38620 52690 38700 52710
rect 37852 52644 37860 52678
rect 37850 52630 37860 52644
rect 37780 52610 37860 52630
rect 37890 52634 38090 52640
rect 37890 52600 37902 52634
rect 38078 52630 38090 52634
rect 38388 52634 38588 52640
rect 38388 52630 38400 52634
rect 38078 52600 38400 52630
rect 38576 52600 38588 52634
rect 38620 52630 38630 52690
rect 38690 52630 38700 52690
rect 38620 52610 38700 52630
rect 37890 52594 38090 52600
rect 37670 52470 37740 52530
rect 37670 52230 37690 52470
rect 37730 52230 37740 52470
rect 38200 52590 38280 52600
rect 38388 52594 38588 52600
rect 38200 52530 38210 52590
rect 38270 52530 38280 52590
rect 38200 52480 38280 52530
rect 38200 52420 38210 52480
rect 38270 52420 38280 52480
rect 37890 52412 38090 52418
rect 37780 52380 37860 52400
rect 37780 52320 37790 52380
rect 37850 52368 37860 52380
rect 37890 52378 37902 52412
rect 38078 52410 38090 52412
rect 38200 52410 38280 52420
rect 38750 52550 38760 52790
rect 38800 52550 38820 52790
rect 38750 52470 38820 52550
rect 38388 52412 38588 52418
rect 38388 52410 38400 52412
rect 38078 52380 38400 52410
rect 38078 52378 38090 52380
rect 37890 52372 38090 52378
rect 38388 52378 38400 52380
rect 38576 52378 38588 52412
rect 38388 52372 38588 52378
rect 38620 52380 38700 52400
rect 37852 52334 37860 52368
rect 37850 52320 37860 52334
rect 37780 52300 37860 52320
rect 37890 52324 38090 52330
rect 37890 52290 37902 52324
rect 38078 52320 38090 52324
rect 38388 52324 38588 52330
rect 38388 52320 38400 52324
rect 38078 52310 38400 52320
rect 38078 52290 38210 52310
rect 37890 52284 38090 52290
rect 38200 52250 38210 52290
rect 38270 52290 38400 52310
rect 38576 52290 38588 52324
rect 38620 52320 38630 52380
rect 38690 52320 38700 52380
rect 38620 52300 38700 52320
rect 38270 52250 38280 52290
rect 38388 52284 38588 52290
rect 38200 52240 38280 52250
rect 37670 51080 37740 52230
rect 37670 50820 37690 51080
rect 37730 50820 37740 51080
rect 38750 52230 38760 52470
rect 38800 52230 38820 52470
rect 38750 51080 38820 52230
rect 38200 51050 38280 51060
rect 37890 51012 38090 51018
rect 37780 50980 37860 51000
rect 37780 50920 37790 50980
rect 37850 50968 37860 50980
rect 37890 50978 37902 51012
rect 38078 51010 38090 51012
rect 38200 51010 38210 51050
rect 38078 50990 38210 51010
rect 38270 51010 38280 51050
rect 38388 51012 38588 51018
rect 38388 51010 38400 51012
rect 38270 50990 38400 51010
rect 38078 50980 38400 50990
rect 38078 50978 38090 50980
rect 37890 50972 38090 50978
rect 38388 50978 38400 50980
rect 38576 50978 38588 51012
rect 38388 50972 38588 50978
rect 38620 50980 38700 51000
rect 37852 50934 37860 50968
rect 37850 50920 37860 50934
rect 37780 50900 37860 50920
rect 37890 50924 38090 50930
rect 37890 50890 37902 50924
rect 38078 50920 38090 50924
rect 38388 50924 38588 50930
rect 38388 50920 38400 50924
rect 38078 50890 38400 50920
rect 38576 50890 38588 50924
rect 38620 50920 38630 50980
rect 38690 50920 38700 50980
rect 38620 50900 38700 50920
rect 37890 50884 38090 50890
rect 37670 50760 37740 50820
rect 37670 50520 37690 50760
rect 37730 50520 37740 50760
rect 38200 50880 38280 50890
rect 38388 50884 38588 50890
rect 38200 50820 38210 50880
rect 38270 50820 38280 50880
rect 38200 50770 38280 50820
rect 38200 50710 38210 50770
rect 38270 50710 38280 50770
rect 37890 50702 38090 50708
rect 37780 50670 37860 50690
rect 37780 50610 37790 50670
rect 37850 50658 37860 50670
rect 37890 50668 37902 50702
rect 38078 50700 38090 50702
rect 38200 50700 38280 50710
rect 38750 50840 38760 51080
rect 38800 50840 38820 51080
rect 38750 50760 38820 50840
rect 38388 50702 38588 50708
rect 38388 50700 38400 50702
rect 38078 50670 38400 50700
rect 38078 50668 38090 50670
rect 37890 50662 38090 50668
rect 38388 50668 38400 50670
rect 38576 50668 38588 50702
rect 38388 50662 38588 50668
rect 38620 50670 38700 50690
rect 37852 50624 37860 50658
rect 37850 50610 37860 50624
rect 37780 50590 37860 50610
rect 37890 50614 38090 50620
rect 37890 50580 37902 50614
rect 38078 50610 38090 50614
rect 38388 50614 38588 50620
rect 38388 50610 38400 50614
rect 38078 50600 38400 50610
rect 38078 50580 38210 50600
rect 37890 50574 38090 50580
rect 38200 50540 38210 50580
rect 38270 50580 38400 50600
rect 38576 50580 38588 50614
rect 38620 50610 38630 50670
rect 38690 50610 38700 50670
rect 38620 50590 38700 50610
rect 38270 50540 38280 50580
rect 38388 50574 38588 50580
rect 38200 50530 38280 50540
rect 37670 49370 37740 50520
rect 37670 49110 37690 49370
rect 37730 49110 37740 49370
rect 38750 50520 38760 50760
rect 38800 50520 38820 50760
rect 38750 49370 38820 50520
rect 38200 49340 38280 49350
rect 37890 49302 38090 49308
rect 37780 49270 37860 49290
rect 37780 49210 37790 49270
rect 37850 49258 37860 49270
rect 37890 49268 37902 49302
rect 38078 49300 38090 49302
rect 38200 49300 38210 49340
rect 38078 49280 38210 49300
rect 38270 49300 38280 49340
rect 38388 49302 38588 49308
rect 38388 49300 38400 49302
rect 38270 49280 38400 49300
rect 38078 49270 38400 49280
rect 38078 49268 38090 49270
rect 37890 49262 38090 49268
rect 38388 49268 38400 49270
rect 38576 49268 38588 49302
rect 38388 49262 38588 49268
rect 38620 49270 38700 49290
rect 37852 49224 37860 49258
rect 37850 49210 37860 49224
rect 37780 49190 37860 49210
rect 37890 49214 38090 49220
rect 37890 49180 37902 49214
rect 38078 49210 38090 49214
rect 38388 49214 38588 49220
rect 38388 49210 38400 49214
rect 38078 49180 38400 49210
rect 38576 49180 38588 49214
rect 38620 49210 38630 49270
rect 38690 49210 38700 49270
rect 38620 49190 38700 49210
rect 37890 49174 38090 49180
rect 37670 49050 37740 49110
rect 37670 48810 37690 49050
rect 37730 48810 37740 49050
rect 38200 49170 38280 49180
rect 38388 49174 38588 49180
rect 38200 49110 38210 49170
rect 38270 49110 38280 49170
rect 38200 49060 38280 49110
rect 38200 49000 38210 49060
rect 38270 49000 38280 49060
rect 37890 48992 38090 48998
rect 37780 48960 37860 48980
rect 37780 48900 37790 48960
rect 37850 48948 37860 48960
rect 37890 48958 37902 48992
rect 38078 48990 38090 48992
rect 38200 48990 38280 49000
rect 38750 49130 38760 49370
rect 38800 49130 38820 49370
rect 38750 49050 38820 49130
rect 38388 48992 38588 48998
rect 38388 48990 38400 48992
rect 38078 48960 38400 48990
rect 38078 48958 38090 48960
rect 37890 48952 38090 48958
rect 38388 48958 38400 48960
rect 38576 48958 38588 48992
rect 38388 48952 38588 48958
rect 38620 48960 38700 48980
rect 37852 48914 37860 48948
rect 37850 48900 37860 48914
rect 37780 48880 37860 48900
rect 37890 48904 38090 48910
rect 37890 48870 37902 48904
rect 38078 48900 38090 48904
rect 38388 48904 38588 48910
rect 38388 48900 38400 48904
rect 38078 48890 38400 48900
rect 38078 48870 38210 48890
rect 37890 48864 38090 48870
rect 38200 48830 38210 48870
rect 38270 48870 38400 48890
rect 38576 48870 38588 48904
rect 38620 48900 38630 48960
rect 38690 48900 38700 48960
rect 38620 48880 38700 48900
rect 38270 48830 38280 48870
rect 38388 48864 38588 48870
rect 38200 48820 38280 48830
rect 37670 47660 37740 48810
rect 37670 47400 37690 47660
rect 37730 47400 37740 47660
rect 38750 48810 38760 49050
rect 38800 48810 38820 49050
rect 38750 47660 38820 48810
rect 38200 47630 38280 47640
rect 37890 47592 38090 47598
rect 37780 47560 37860 47580
rect 37780 47500 37790 47560
rect 37850 47548 37860 47560
rect 37890 47558 37902 47592
rect 38078 47590 38090 47592
rect 38200 47590 38210 47630
rect 38078 47570 38210 47590
rect 38270 47590 38280 47630
rect 38388 47592 38588 47598
rect 38388 47590 38400 47592
rect 38270 47570 38400 47590
rect 38078 47560 38400 47570
rect 38078 47558 38090 47560
rect 37890 47552 38090 47558
rect 38388 47558 38400 47560
rect 38576 47558 38588 47592
rect 38388 47552 38588 47558
rect 38620 47560 38700 47580
rect 37852 47514 37860 47548
rect 37850 47500 37860 47514
rect 37780 47480 37860 47500
rect 37890 47504 38090 47510
rect 37890 47470 37902 47504
rect 38078 47500 38090 47504
rect 38388 47504 38588 47510
rect 38388 47500 38400 47504
rect 38078 47470 38400 47500
rect 38576 47470 38588 47504
rect 38620 47500 38630 47560
rect 38690 47500 38700 47560
rect 38620 47480 38700 47500
rect 37890 47464 38090 47470
rect 37670 47340 37740 47400
rect 37670 47100 37690 47340
rect 37730 47100 37740 47340
rect 38200 47460 38280 47470
rect 38388 47464 38588 47470
rect 38200 47400 38210 47460
rect 38270 47400 38280 47460
rect 38200 47350 38280 47400
rect 38200 47290 38210 47350
rect 38270 47290 38280 47350
rect 37890 47282 38090 47288
rect 37780 47250 37860 47270
rect 37780 47190 37790 47250
rect 37850 47238 37860 47250
rect 37890 47248 37902 47282
rect 38078 47280 38090 47282
rect 38200 47280 38280 47290
rect 38750 47420 38760 47660
rect 38800 47420 38820 47660
rect 38750 47340 38820 47420
rect 38388 47282 38588 47288
rect 38388 47280 38400 47282
rect 38078 47250 38400 47280
rect 38078 47248 38090 47250
rect 37890 47242 38090 47248
rect 38388 47248 38400 47250
rect 38576 47248 38588 47282
rect 38388 47242 38588 47248
rect 38620 47250 38700 47270
rect 37852 47204 37860 47238
rect 37850 47190 37860 47204
rect 37780 47170 37860 47190
rect 37890 47194 38090 47200
rect 37890 47160 37902 47194
rect 38078 47190 38090 47194
rect 38388 47194 38588 47200
rect 38388 47190 38400 47194
rect 38078 47180 38400 47190
rect 38078 47160 38210 47180
rect 37890 47154 38090 47160
rect 38200 47120 38210 47160
rect 38270 47160 38400 47180
rect 38576 47160 38588 47194
rect 38620 47190 38630 47250
rect 38690 47190 38700 47250
rect 38620 47170 38700 47190
rect 38270 47120 38280 47160
rect 38388 47154 38588 47160
rect 38200 47110 38280 47120
rect 37670 45950 37740 47100
rect 37670 45690 37690 45950
rect 37730 45690 37740 45950
rect 38750 47100 38760 47340
rect 38800 47100 38820 47340
rect 38750 45950 38820 47100
rect 38200 45920 38280 45930
rect 37890 45882 38090 45888
rect 37780 45850 37860 45870
rect 37780 45790 37790 45850
rect 37850 45838 37860 45850
rect 37890 45848 37902 45882
rect 38078 45880 38090 45882
rect 38200 45880 38210 45920
rect 38078 45860 38210 45880
rect 38270 45880 38280 45920
rect 38388 45882 38588 45888
rect 38388 45880 38400 45882
rect 38270 45860 38400 45880
rect 38078 45850 38400 45860
rect 38078 45848 38090 45850
rect 37890 45842 38090 45848
rect 38388 45848 38400 45850
rect 38576 45848 38588 45882
rect 38388 45842 38588 45848
rect 38620 45850 38700 45870
rect 37852 45804 37860 45838
rect 37850 45790 37860 45804
rect 37780 45770 37860 45790
rect 37890 45794 38090 45800
rect 37890 45760 37902 45794
rect 38078 45790 38090 45794
rect 38388 45794 38588 45800
rect 38388 45790 38400 45794
rect 38078 45760 38400 45790
rect 38576 45760 38588 45794
rect 38620 45790 38630 45850
rect 38690 45790 38700 45850
rect 38620 45770 38700 45790
rect 37890 45754 38090 45760
rect 37670 45630 37740 45690
rect 37670 45390 37690 45630
rect 37730 45390 37740 45630
rect 38200 45750 38280 45760
rect 38388 45754 38588 45760
rect 38200 45690 38210 45750
rect 38270 45690 38280 45750
rect 38200 45640 38280 45690
rect 38200 45580 38210 45640
rect 38270 45580 38280 45640
rect 37890 45572 38090 45578
rect 37780 45540 37860 45560
rect 37780 45480 37790 45540
rect 37850 45528 37860 45540
rect 37890 45538 37902 45572
rect 38078 45570 38090 45572
rect 38200 45570 38280 45580
rect 38750 45710 38760 45950
rect 38800 45710 38820 45950
rect 38750 45630 38820 45710
rect 38388 45572 38588 45578
rect 38388 45570 38400 45572
rect 38078 45540 38400 45570
rect 38078 45538 38090 45540
rect 37890 45532 38090 45538
rect 38388 45538 38400 45540
rect 38576 45538 38588 45572
rect 38388 45532 38588 45538
rect 38620 45540 38700 45560
rect 37852 45494 37860 45528
rect 37850 45480 37860 45494
rect 37780 45460 37860 45480
rect 37890 45484 38090 45490
rect 37890 45450 37902 45484
rect 38078 45480 38090 45484
rect 38388 45484 38588 45490
rect 38388 45480 38400 45484
rect 38078 45470 38400 45480
rect 38078 45450 38210 45470
rect 37890 45444 38090 45450
rect 38200 45410 38210 45450
rect 38270 45450 38400 45470
rect 38576 45450 38588 45484
rect 38620 45480 38630 45540
rect 38690 45480 38700 45540
rect 38620 45460 38700 45480
rect 38270 45410 38280 45450
rect 38388 45444 38588 45450
rect 38200 45400 38280 45410
rect 37670 44240 37740 45390
rect 37670 43980 37690 44240
rect 37730 43980 37740 44240
rect 38750 45390 38760 45630
rect 38800 45390 38820 45630
rect 38750 44240 38820 45390
rect 38200 44210 38280 44220
rect 37890 44172 38090 44178
rect 37780 44140 37860 44160
rect 37780 44080 37790 44140
rect 37850 44128 37860 44140
rect 37890 44138 37902 44172
rect 38078 44170 38090 44172
rect 38200 44170 38210 44210
rect 38078 44150 38210 44170
rect 38270 44170 38280 44210
rect 38388 44172 38588 44178
rect 38388 44170 38400 44172
rect 38270 44150 38400 44170
rect 38078 44140 38400 44150
rect 38078 44138 38090 44140
rect 37890 44132 38090 44138
rect 38388 44138 38400 44140
rect 38576 44138 38588 44172
rect 38388 44132 38588 44138
rect 38620 44140 38700 44160
rect 37852 44094 37860 44128
rect 37850 44080 37860 44094
rect 37780 44060 37860 44080
rect 37890 44084 38090 44090
rect 37890 44050 37902 44084
rect 38078 44080 38090 44084
rect 38388 44084 38588 44090
rect 38388 44080 38400 44084
rect 38078 44050 38400 44080
rect 38576 44050 38588 44084
rect 38620 44080 38630 44140
rect 38690 44080 38700 44140
rect 38620 44060 38700 44080
rect 37890 44044 38090 44050
rect 37670 43920 37740 43980
rect 37670 43680 37690 43920
rect 37730 43680 37740 43920
rect 38200 44040 38280 44050
rect 38388 44044 38588 44050
rect 38200 43980 38210 44040
rect 38270 43980 38280 44040
rect 38200 43930 38280 43980
rect 38200 43870 38210 43930
rect 38270 43870 38280 43930
rect 37890 43862 38090 43868
rect 37780 43830 37860 43850
rect 37780 43770 37790 43830
rect 37850 43818 37860 43830
rect 37890 43828 37902 43862
rect 38078 43860 38090 43862
rect 38200 43860 38280 43870
rect 38750 44000 38760 44240
rect 38800 44000 38820 44240
rect 38750 43920 38820 44000
rect 38388 43862 38588 43868
rect 38388 43860 38400 43862
rect 38078 43830 38400 43860
rect 38078 43828 38090 43830
rect 37890 43822 38090 43828
rect 38388 43828 38400 43830
rect 38576 43828 38588 43862
rect 38388 43822 38588 43828
rect 38620 43830 38700 43850
rect 37852 43784 37860 43818
rect 37850 43770 37860 43784
rect 37780 43750 37860 43770
rect 37890 43774 38090 43780
rect 37890 43740 37902 43774
rect 38078 43770 38090 43774
rect 38388 43774 38588 43780
rect 38388 43770 38400 43774
rect 38078 43760 38400 43770
rect 38078 43740 38210 43760
rect 37890 43734 38090 43740
rect 38200 43700 38210 43740
rect 38270 43740 38400 43760
rect 38576 43740 38588 43774
rect 38620 43770 38630 43830
rect 38690 43770 38700 43830
rect 38620 43750 38700 43770
rect 38270 43700 38280 43740
rect 38388 43734 38588 43740
rect 38200 43690 38280 43700
rect 37670 42530 37740 43680
rect 37670 42270 37690 42530
rect 37730 42270 37740 42530
rect 38750 43680 38760 43920
rect 38800 43680 38820 43920
rect 38750 42530 38820 43680
rect 38200 42500 38280 42510
rect 37890 42462 38090 42468
rect 37780 42430 37860 42450
rect 37780 42370 37790 42430
rect 37850 42418 37860 42430
rect 37890 42428 37902 42462
rect 38078 42460 38090 42462
rect 38200 42460 38210 42500
rect 38078 42440 38210 42460
rect 38270 42460 38280 42500
rect 38388 42462 38588 42468
rect 38388 42460 38400 42462
rect 38270 42440 38400 42460
rect 38078 42430 38400 42440
rect 38078 42428 38090 42430
rect 37890 42422 38090 42428
rect 38388 42428 38400 42430
rect 38576 42428 38588 42462
rect 38388 42422 38588 42428
rect 38620 42430 38700 42450
rect 37852 42384 37860 42418
rect 37850 42370 37860 42384
rect 37780 42350 37860 42370
rect 37890 42374 38090 42380
rect 37890 42340 37902 42374
rect 38078 42370 38090 42374
rect 38388 42374 38588 42380
rect 38388 42370 38400 42374
rect 38078 42340 38400 42370
rect 38576 42340 38588 42374
rect 38620 42370 38630 42430
rect 38690 42370 38700 42430
rect 38620 42350 38700 42370
rect 37890 42334 38090 42340
rect 37670 42210 37740 42270
rect 37670 41970 37690 42210
rect 37730 41970 37740 42210
rect 38200 42330 38280 42340
rect 38388 42334 38588 42340
rect 38200 42270 38210 42330
rect 38270 42270 38280 42330
rect 38200 42220 38280 42270
rect 38200 42160 38210 42220
rect 38270 42160 38280 42220
rect 37890 42152 38090 42158
rect 37780 42120 37860 42140
rect 37780 42060 37790 42120
rect 37850 42108 37860 42120
rect 37890 42118 37902 42152
rect 38078 42150 38090 42152
rect 38200 42150 38280 42160
rect 38750 42290 38760 42530
rect 38800 42290 38820 42530
rect 38750 42210 38820 42290
rect 38388 42152 38588 42158
rect 38388 42150 38400 42152
rect 38078 42120 38400 42150
rect 38078 42118 38090 42120
rect 37890 42112 38090 42118
rect 38388 42118 38400 42120
rect 38576 42118 38588 42152
rect 38388 42112 38588 42118
rect 38620 42120 38700 42140
rect 37852 42074 37860 42108
rect 37850 42060 37860 42074
rect 37780 42040 37860 42060
rect 37890 42064 38090 42070
rect 37890 42030 37902 42064
rect 38078 42060 38090 42064
rect 38388 42064 38588 42070
rect 38388 42060 38400 42064
rect 38078 42050 38400 42060
rect 38078 42030 38210 42050
rect 37890 42024 38090 42030
rect 38200 41990 38210 42030
rect 38270 42030 38400 42050
rect 38576 42030 38588 42064
rect 38620 42060 38630 42120
rect 38690 42060 38700 42120
rect 38620 42040 38700 42060
rect 38270 41990 38280 42030
rect 38388 42024 38588 42030
rect 38200 41980 38280 41990
rect 37670 40820 37740 41970
rect 37670 40560 37690 40820
rect 37730 40560 37740 40820
rect 38750 41970 38760 42210
rect 38800 41970 38820 42210
rect 38750 40820 38820 41970
rect 38200 40790 38280 40800
rect 37890 40752 38090 40758
rect 37780 40720 37860 40740
rect 37780 40660 37790 40720
rect 37850 40708 37860 40720
rect 37890 40718 37902 40752
rect 38078 40750 38090 40752
rect 38200 40750 38210 40790
rect 38078 40730 38210 40750
rect 38270 40750 38280 40790
rect 38388 40752 38588 40758
rect 38388 40750 38400 40752
rect 38270 40730 38400 40750
rect 38078 40720 38400 40730
rect 38078 40718 38090 40720
rect 37890 40712 38090 40718
rect 38388 40718 38400 40720
rect 38576 40718 38588 40752
rect 38388 40712 38588 40718
rect 38620 40720 38700 40740
rect 37852 40674 37860 40708
rect 37850 40660 37860 40674
rect 37780 40640 37860 40660
rect 37890 40664 38090 40670
rect 37890 40630 37902 40664
rect 38078 40660 38090 40664
rect 38388 40664 38588 40670
rect 38388 40660 38400 40664
rect 38078 40630 38400 40660
rect 38576 40630 38588 40664
rect 38620 40660 38630 40720
rect 38690 40660 38700 40720
rect 38620 40640 38700 40660
rect 37890 40624 38090 40630
rect 37670 40500 37740 40560
rect 37670 40260 37690 40500
rect 37730 40260 37740 40500
rect 38200 40620 38280 40630
rect 38388 40624 38588 40630
rect 38200 40560 38210 40620
rect 38270 40560 38280 40620
rect 38200 40510 38280 40560
rect 38200 40450 38210 40510
rect 38270 40450 38280 40510
rect 37890 40442 38090 40448
rect 37780 40410 37860 40430
rect 37780 40350 37790 40410
rect 37850 40398 37860 40410
rect 37890 40408 37902 40442
rect 38078 40440 38090 40442
rect 38200 40440 38280 40450
rect 38750 40580 38760 40820
rect 38800 40580 38820 40820
rect 38750 40500 38820 40580
rect 38388 40442 38588 40448
rect 38388 40440 38400 40442
rect 38078 40410 38400 40440
rect 38078 40408 38090 40410
rect 37890 40402 38090 40408
rect 38388 40408 38400 40410
rect 38576 40408 38588 40442
rect 38388 40402 38588 40408
rect 38620 40410 38700 40430
rect 37852 40364 37860 40398
rect 37850 40350 37860 40364
rect 37780 40330 37860 40350
rect 37890 40354 38090 40360
rect 37890 40320 37902 40354
rect 38078 40350 38090 40354
rect 38388 40354 38588 40360
rect 38388 40350 38400 40354
rect 38078 40340 38400 40350
rect 38078 40320 38210 40340
rect 37890 40314 38090 40320
rect 38200 40280 38210 40320
rect 38270 40320 38400 40340
rect 38576 40320 38588 40354
rect 38620 40350 38630 40410
rect 38690 40350 38700 40410
rect 38620 40330 38700 40350
rect 38270 40280 38280 40320
rect 38388 40314 38588 40320
rect 38200 40270 38280 40280
rect 37670 39690 37740 40260
rect 38750 40260 38760 40500
rect 38800 40260 38820 40500
rect 38750 39690 38820 40260
rect 37670 39680 37750 39690
rect 37670 39620 37680 39680
rect 37740 39620 37750 39680
rect 38740 39680 38820 39690
rect 38740 39620 38750 39680
rect 38810 39620 38820 39680
rect 38740 39610 38820 39620
rect 38850 66480 38880 67050
rect 38850 66470 38910 66480
rect 38850 66400 38910 66410
rect 38850 64770 38880 66400
rect 38940 65950 38970 67050
rect 38910 65940 38970 65950
rect 38910 65870 38970 65880
rect 38850 64760 38910 64770
rect 38850 64690 38910 64700
rect 38850 63060 38880 64690
rect 38940 64240 38970 65870
rect 38910 64230 38970 64240
rect 38910 64160 38970 64170
rect 38850 63050 38910 63060
rect 38850 62980 38910 62990
rect 38850 61350 38880 62980
rect 38940 62530 38970 64160
rect 38910 62520 38970 62530
rect 38910 62450 38970 62460
rect 38850 61340 38910 61350
rect 38850 61270 38910 61280
rect 38850 59640 38880 61270
rect 38940 60820 38970 62450
rect 38910 60810 38970 60820
rect 38910 60740 38970 60750
rect 38850 59630 38910 59640
rect 38850 59560 38910 59570
rect 38850 57930 38880 59560
rect 38940 59110 38970 60740
rect 38910 59100 38970 59110
rect 38910 59030 38970 59040
rect 38850 57920 38910 57930
rect 38850 57850 38910 57860
rect 38850 56220 38880 57850
rect 38940 57400 38970 59030
rect 38910 57390 38970 57400
rect 38910 57320 38970 57330
rect 38850 56210 38910 56220
rect 38850 56140 38910 56150
rect 38850 54510 38880 56140
rect 38940 55690 38970 57320
rect 38910 55680 38970 55690
rect 38910 55610 38970 55620
rect 38850 54500 38910 54510
rect 38850 54430 38910 54440
rect 38850 52800 38880 54430
rect 38940 53980 38970 55610
rect 38910 53970 38970 53980
rect 38910 53900 38970 53910
rect 38850 52790 38910 52800
rect 38850 52720 38910 52730
rect 38850 51090 38880 52720
rect 38940 52270 38970 53900
rect 38910 52260 38970 52270
rect 38910 52190 38970 52200
rect 38850 51080 38910 51090
rect 38850 51010 38910 51020
rect 38850 49380 38880 51010
rect 38940 50560 38970 52190
rect 38910 50550 38970 50560
rect 38910 50480 38970 50490
rect 38850 49370 38910 49380
rect 38850 49300 38910 49310
rect 38850 47670 38880 49300
rect 38940 48850 38970 50480
rect 38910 48840 38970 48850
rect 38910 48770 38970 48780
rect 38850 47660 38910 47670
rect 38850 47590 38910 47600
rect 38850 45960 38880 47590
rect 38940 47140 38970 48770
rect 38910 47130 38970 47140
rect 38910 47060 38970 47070
rect 38850 45950 38910 45960
rect 38850 45880 38910 45890
rect 38850 44250 38880 45880
rect 38940 45430 38970 47060
rect 38910 45420 38970 45430
rect 38910 45350 38970 45360
rect 38850 44240 38910 44250
rect 38850 44170 38910 44180
rect 38850 42540 38880 44170
rect 38940 43720 38970 45350
rect 38910 43710 38970 43720
rect 38910 43640 38970 43650
rect 38850 42530 38910 42540
rect 38850 42460 38910 42470
rect 38850 40830 38880 42460
rect 38940 42010 38970 43640
rect 38910 42000 38970 42010
rect 38910 41930 38970 41940
rect 38850 40820 38910 40830
rect 38850 40750 38910 40760
rect 37200 39220 37260 39230
rect 37380 39230 37640 39240
rect 34210 39160 34270 39170
rect 37440 39210 37640 39230
rect 37380 39160 37440 39170
rect 38850 38840 38880 40750
rect 38940 40300 38970 41930
rect 38910 40290 38970 40300
rect 38910 40220 38970 40230
rect 38940 39690 38970 40220
rect 38910 39680 38970 39690
rect 38910 39610 38970 39620
rect 39000 66390 39030 67050
rect 39000 66380 39060 66390
rect 39000 66310 39060 66320
rect 39000 64680 39030 66310
rect 39000 64670 39060 64680
rect 39000 64600 39060 64610
rect 39000 42440 39030 64600
rect 39120 62970 39150 67050
rect 39120 62960 39180 62970
rect 39120 62890 39180 62900
rect 39120 61260 39150 62890
rect 39120 61250 39180 61260
rect 39120 61180 39180 61190
rect 39120 45870 39150 61180
rect 39240 59550 39270 67050
rect 39240 59540 39300 59550
rect 39240 59470 39300 59480
rect 39240 47580 39270 59470
rect 39360 57840 39390 67050
rect 39360 57830 39420 57840
rect 39360 57760 39420 57770
rect 39360 49290 39390 57760
rect 39480 56130 39510 67050
rect 39480 56120 39540 56130
rect 39480 56050 39540 56060
rect 39480 51000 39510 56050
rect 39600 52710 39630 67050
rect 39720 54410 39750 67050
rect 41880 54410 41910 67050
rect 39720 54400 39780 54410
rect 39720 54330 39780 54340
rect 41850 54400 41910 54410
rect 41850 54330 41910 54340
rect 39600 52700 39660 52710
rect 39600 52630 39660 52640
rect 39480 50990 39540 51000
rect 39480 50920 39540 50930
rect 39360 49280 39420 49290
rect 39360 49210 39420 49220
rect 39240 47570 39300 47580
rect 39240 47500 39300 47510
rect 39120 45860 39180 45870
rect 39120 45790 39180 45800
rect 39120 44150 39150 45790
rect 39120 44140 39180 44150
rect 39120 44070 39180 44080
rect 39000 42430 39060 42440
rect 39000 42360 39060 42370
rect 39000 40740 39030 42360
rect 39000 40730 39060 40740
rect 39000 40660 39060 40670
rect 39000 39240 39030 40660
rect 39120 39300 39150 44070
rect 39240 39360 39270 47500
rect 39360 39420 39390 49210
rect 39480 39480 39510 50920
rect 39600 39540 39630 52630
rect 39720 39600 39750 54330
rect 41880 39600 41910 54330
rect 42000 52710 42030 67050
rect 42120 56130 42150 67050
rect 42240 57840 42270 67050
rect 42360 59550 42390 67050
rect 42480 62970 42510 67050
rect 42600 66390 42630 67050
rect 42570 66380 42630 66390
rect 42570 66310 42630 66320
rect 42600 64680 42630 66310
rect 42570 64670 42630 64680
rect 42570 64600 42630 64610
rect 42450 62960 42510 62970
rect 42450 62890 42510 62900
rect 42480 61260 42510 62890
rect 42450 61250 42510 61260
rect 42450 61180 42510 61190
rect 42330 59540 42390 59550
rect 42330 59470 42390 59480
rect 42210 57830 42270 57840
rect 42210 57760 42270 57770
rect 42090 56120 42150 56130
rect 42090 56050 42150 56060
rect 41970 52700 42030 52710
rect 41970 52630 42030 52640
rect 39720 39590 40340 39600
rect 39720 39570 40280 39590
rect 39600 39530 40160 39540
rect 39600 39510 40100 39530
rect 39480 39470 39980 39480
rect 39480 39450 39920 39470
rect 39360 39410 39800 39420
rect 39360 39390 39740 39410
rect 39240 39350 39620 39360
rect 39240 39330 39560 39350
rect 39120 39290 39440 39300
rect 39120 39270 39380 39290
rect 39000 39230 39260 39240
rect 39000 39210 39200 39230
rect 40280 39520 40340 39530
rect 41290 39590 41910 39600
rect 41350 39570 41910 39590
rect 42000 39540 42030 52630
rect 42120 51000 42150 56050
rect 42090 50990 42150 51000
rect 42090 50920 42150 50930
rect 41290 39520 41350 39530
rect 41470 39530 42030 39540
rect 40100 39460 40160 39470
rect 41530 39510 42030 39530
rect 42120 39480 42150 50920
rect 42240 49290 42270 57760
rect 42210 49280 42270 49290
rect 42210 49210 42270 49220
rect 41470 39460 41530 39470
rect 41650 39470 42150 39480
rect 39920 39400 39980 39410
rect 41710 39450 42150 39470
rect 42240 39420 42270 49210
rect 42360 47580 42390 59470
rect 42330 47570 42390 47580
rect 42330 47500 42390 47510
rect 41650 39400 41710 39410
rect 41830 39410 42270 39420
rect 39740 39340 39800 39350
rect 41890 39390 42270 39410
rect 42360 39360 42390 47500
rect 42480 45870 42510 61180
rect 42450 45860 42510 45870
rect 42450 45790 42510 45800
rect 42480 44160 42510 45790
rect 42450 44150 42510 44160
rect 42450 44080 42510 44090
rect 41830 39340 41890 39350
rect 42010 39350 42390 39360
rect 39560 39280 39620 39290
rect 42070 39330 42390 39350
rect 42480 39300 42510 44080
rect 42600 42450 42630 64600
rect 42570 42440 42630 42450
rect 42570 42370 42630 42380
rect 42600 40740 42630 42370
rect 42570 40730 42630 40740
rect 42570 40660 42630 40670
rect 42010 39280 42070 39290
rect 42190 39290 42510 39300
rect 39380 39220 39440 39230
rect 42250 39270 42510 39290
rect 42600 39240 42630 40660
rect 42660 66470 42730 67050
rect 42660 66210 42680 66470
rect 42720 66210 42730 66470
rect 43740 66470 43810 67050
rect 43190 66440 43270 66450
rect 42880 66402 43080 66408
rect 42770 66370 42850 66390
rect 42770 66310 42780 66370
rect 42840 66358 42850 66370
rect 42880 66368 42892 66402
rect 43068 66400 43080 66402
rect 43190 66400 43200 66440
rect 43068 66380 43200 66400
rect 43260 66400 43270 66440
rect 43378 66402 43578 66408
rect 43378 66400 43390 66402
rect 43260 66380 43390 66400
rect 43068 66370 43390 66380
rect 43068 66368 43080 66370
rect 42880 66362 43080 66368
rect 43378 66368 43390 66370
rect 43566 66368 43578 66402
rect 43378 66362 43578 66368
rect 43610 66370 43690 66390
rect 42842 66324 42850 66358
rect 42840 66310 42850 66324
rect 42770 66290 42850 66310
rect 42880 66314 43080 66320
rect 42880 66280 42892 66314
rect 43068 66310 43080 66314
rect 43378 66314 43578 66320
rect 43378 66310 43390 66314
rect 43068 66280 43390 66310
rect 43566 66280 43578 66314
rect 43610 66310 43620 66370
rect 43680 66310 43690 66370
rect 43610 66290 43690 66310
rect 42880 66274 43080 66280
rect 42660 66150 42730 66210
rect 42660 65910 42680 66150
rect 42720 65910 42730 66150
rect 43190 66270 43270 66280
rect 43378 66274 43578 66280
rect 43190 66210 43200 66270
rect 43260 66210 43270 66270
rect 43190 66160 43270 66210
rect 43190 66100 43200 66160
rect 43260 66100 43270 66160
rect 42880 66092 43080 66098
rect 42770 66060 42850 66080
rect 42770 66000 42780 66060
rect 42840 66048 42850 66060
rect 42880 66058 42892 66092
rect 43068 66090 43080 66092
rect 43190 66090 43270 66100
rect 43740 66230 43750 66470
rect 43790 66230 43810 66470
rect 43740 66150 43810 66230
rect 43378 66092 43578 66098
rect 43378 66090 43390 66092
rect 43068 66060 43390 66090
rect 43068 66058 43080 66060
rect 42880 66052 43080 66058
rect 43378 66058 43390 66060
rect 43566 66058 43578 66092
rect 43378 66052 43578 66058
rect 43610 66060 43690 66080
rect 42842 66014 42850 66048
rect 42840 66000 42850 66014
rect 42770 65980 42850 66000
rect 42880 66004 43080 66010
rect 42880 65970 42892 66004
rect 43068 66000 43080 66004
rect 43378 66004 43578 66010
rect 43378 66000 43390 66004
rect 43068 65990 43390 66000
rect 43068 65970 43200 65990
rect 42880 65964 43080 65970
rect 43190 65930 43200 65970
rect 43260 65970 43390 65990
rect 43566 65970 43578 66004
rect 43610 66000 43620 66060
rect 43680 66000 43690 66060
rect 43610 65980 43690 66000
rect 43260 65930 43270 65970
rect 43378 65964 43578 65970
rect 43190 65920 43270 65930
rect 42660 64760 42730 65910
rect 42660 64500 42680 64760
rect 42720 64500 42730 64760
rect 43740 65910 43750 66150
rect 43790 65910 43810 66150
rect 43740 64760 43810 65910
rect 43190 64730 43270 64740
rect 42880 64692 43080 64698
rect 42770 64660 42850 64680
rect 42770 64600 42780 64660
rect 42840 64648 42850 64660
rect 42880 64658 42892 64692
rect 43068 64690 43080 64692
rect 43190 64690 43200 64730
rect 43068 64670 43200 64690
rect 43260 64690 43270 64730
rect 43378 64692 43578 64698
rect 43378 64690 43390 64692
rect 43260 64670 43390 64690
rect 43068 64660 43390 64670
rect 43068 64658 43080 64660
rect 42880 64652 43080 64658
rect 43378 64658 43390 64660
rect 43566 64658 43578 64692
rect 43378 64652 43578 64658
rect 43610 64660 43690 64680
rect 42842 64614 42850 64648
rect 42840 64600 42850 64614
rect 42770 64580 42850 64600
rect 42880 64604 43080 64610
rect 42880 64570 42892 64604
rect 43068 64600 43080 64604
rect 43378 64604 43578 64610
rect 43378 64600 43390 64604
rect 43068 64570 43390 64600
rect 43566 64570 43578 64604
rect 43610 64600 43620 64660
rect 43680 64600 43690 64660
rect 43610 64580 43690 64600
rect 42880 64564 43080 64570
rect 42660 64440 42730 64500
rect 42660 64200 42680 64440
rect 42720 64200 42730 64440
rect 43190 64560 43270 64570
rect 43378 64564 43578 64570
rect 43190 64500 43200 64560
rect 43260 64500 43270 64560
rect 43190 64450 43270 64500
rect 43190 64390 43200 64450
rect 43260 64390 43270 64450
rect 42880 64382 43080 64388
rect 42770 64350 42850 64370
rect 42770 64290 42780 64350
rect 42840 64338 42850 64350
rect 42880 64348 42892 64382
rect 43068 64380 43080 64382
rect 43190 64380 43270 64390
rect 43740 64520 43750 64760
rect 43790 64520 43810 64760
rect 43740 64440 43810 64520
rect 43378 64382 43578 64388
rect 43378 64380 43390 64382
rect 43068 64350 43390 64380
rect 43068 64348 43080 64350
rect 42880 64342 43080 64348
rect 43378 64348 43390 64350
rect 43566 64348 43578 64382
rect 43378 64342 43578 64348
rect 43610 64350 43690 64370
rect 42842 64304 42850 64338
rect 42840 64290 42850 64304
rect 42770 64270 42850 64290
rect 42880 64294 43080 64300
rect 42880 64260 42892 64294
rect 43068 64290 43080 64294
rect 43378 64294 43578 64300
rect 43378 64290 43390 64294
rect 43068 64280 43390 64290
rect 43068 64260 43200 64280
rect 42880 64254 43080 64260
rect 43190 64220 43200 64260
rect 43260 64260 43390 64280
rect 43566 64260 43578 64294
rect 43610 64290 43620 64350
rect 43680 64290 43690 64350
rect 43610 64270 43690 64290
rect 43260 64220 43270 64260
rect 43378 64254 43578 64260
rect 43190 64210 43270 64220
rect 42660 63050 42730 64200
rect 42660 62790 42680 63050
rect 42720 62790 42730 63050
rect 43740 64200 43750 64440
rect 43790 64200 43810 64440
rect 43740 63050 43810 64200
rect 43190 63020 43270 63030
rect 42880 62982 43080 62988
rect 42770 62950 42850 62970
rect 42770 62890 42780 62950
rect 42840 62938 42850 62950
rect 42880 62948 42892 62982
rect 43068 62980 43080 62982
rect 43190 62980 43200 63020
rect 43068 62960 43200 62980
rect 43260 62980 43270 63020
rect 43378 62982 43578 62988
rect 43378 62980 43390 62982
rect 43260 62960 43390 62980
rect 43068 62950 43390 62960
rect 43068 62948 43080 62950
rect 42880 62942 43080 62948
rect 43378 62948 43390 62950
rect 43566 62948 43578 62982
rect 43378 62942 43578 62948
rect 43610 62950 43690 62970
rect 42842 62904 42850 62938
rect 42840 62890 42850 62904
rect 42770 62870 42850 62890
rect 42880 62894 43080 62900
rect 42880 62860 42892 62894
rect 43068 62890 43080 62894
rect 43378 62894 43578 62900
rect 43378 62890 43390 62894
rect 43068 62860 43390 62890
rect 43566 62860 43578 62894
rect 43610 62890 43620 62950
rect 43680 62890 43690 62950
rect 43610 62870 43690 62890
rect 42880 62854 43080 62860
rect 42660 62730 42730 62790
rect 42660 62490 42680 62730
rect 42720 62490 42730 62730
rect 43190 62850 43270 62860
rect 43378 62854 43578 62860
rect 43190 62790 43200 62850
rect 43260 62790 43270 62850
rect 43190 62740 43270 62790
rect 43190 62680 43200 62740
rect 43260 62680 43270 62740
rect 42880 62672 43080 62678
rect 42770 62640 42850 62660
rect 42770 62580 42780 62640
rect 42840 62628 42850 62640
rect 42880 62638 42892 62672
rect 43068 62670 43080 62672
rect 43190 62670 43270 62680
rect 43740 62810 43750 63050
rect 43790 62810 43810 63050
rect 43740 62730 43810 62810
rect 43378 62672 43578 62678
rect 43378 62670 43390 62672
rect 43068 62640 43390 62670
rect 43068 62638 43080 62640
rect 42880 62632 43080 62638
rect 43378 62638 43390 62640
rect 43566 62638 43578 62672
rect 43378 62632 43578 62638
rect 43610 62640 43690 62660
rect 42842 62594 42850 62628
rect 42840 62580 42850 62594
rect 42770 62560 42850 62580
rect 42880 62584 43080 62590
rect 42880 62550 42892 62584
rect 43068 62580 43080 62584
rect 43378 62584 43578 62590
rect 43378 62580 43390 62584
rect 43068 62570 43390 62580
rect 43068 62550 43200 62570
rect 42880 62544 43080 62550
rect 43190 62510 43200 62550
rect 43260 62550 43390 62570
rect 43566 62550 43578 62584
rect 43610 62580 43620 62640
rect 43680 62580 43690 62640
rect 43610 62560 43690 62580
rect 43260 62510 43270 62550
rect 43378 62544 43578 62550
rect 43190 62500 43270 62510
rect 42660 61340 42730 62490
rect 42660 61080 42680 61340
rect 42720 61080 42730 61340
rect 43740 62490 43750 62730
rect 43790 62490 43810 62730
rect 43740 61340 43810 62490
rect 43190 61310 43270 61320
rect 42880 61272 43080 61278
rect 42770 61240 42850 61260
rect 42770 61180 42780 61240
rect 42840 61228 42850 61240
rect 42880 61238 42892 61272
rect 43068 61270 43080 61272
rect 43190 61270 43200 61310
rect 43068 61250 43200 61270
rect 43260 61270 43270 61310
rect 43378 61272 43578 61278
rect 43378 61270 43390 61272
rect 43260 61250 43390 61270
rect 43068 61240 43390 61250
rect 43068 61238 43080 61240
rect 42880 61232 43080 61238
rect 43378 61238 43390 61240
rect 43566 61238 43578 61272
rect 43378 61232 43578 61238
rect 43610 61240 43690 61260
rect 42842 61194 42850 61228
rect 42840 61180 42850 61194
rect 42770 61160 42850 61180
rect 42880 61184 43080 61190
rect 42880 61150 42892 61184
rect 43068 61180 43080 61184
rect 43378 61184 43578 61190
rect 43378 61180 43390 61184
rect 43068 61150 43390 61180
rect 43566 61150 43578 61184
rect 43610 61180 43620 61240
rect 43680 61180 43690 61240
rect 43610 61160 43690 61180
rect 42880 61144 43080 61150
rect 42660 61020 42730 61080
rect 42660 60780 42680 61020
rect 42720 60780 42730 61020
rect 43190 61140 43270 61150
rect 43378 61144 43578 61150
rect 43190 61080 43200 61140
rect 43260 61080 43270 61140
rect 43190 61030 43270 61080
rect 43190 60970 43200 61030
rect 43260 60970 43270 61030
rect 42880 60962 43080 60968
rect 42770 60930 42850 60950
rect 42770 60870 42780 60930
rect 42840 60918 42850 60930
rect 42880 60928 42892 60962
rect 43068 60960 43080 60962
rect 43190 60960 43270 60970
rect 43740 61100 43750 61340
rect 43790 61100 43810 61340
rect 43740 61020 43810 61100
rect 43378 60962 43578 60968
rect 43378 60960 43390 60962
rect 43068 60930 43390 60960
rect 43068 60928 43080 60930
rect 42880 60922 43080 60928
rect 43378 60928 43390 60930
rect 43566 60928 43578 60962
rect 43378 60922 43578 60928
rect 43610 60930 43690 60950
rect 42842 60884 42850 60918
rect 42840 60870 42850 60884
rect 42770 60850 42850 60870
rect 42880 60874 43080 60880
rect 42880 60840 42892 60874
rect 43068 60870 43080 60874
rect 43378 60874 43578 60880
rect 43378 60870 43390 60874
rect 43068 60860 43390 60870
rect 43068 60840 43200 60860
rect 42880 60834 43080 60840
rect 43190 60800 43200 60840
rect 43260 60840 43390 60860
rect 43566 60840 43578 60874
rect 43610 60870 43620 60930
rect 43680 60870 43690 60930
rect 43610 60850 43690 60870
rect 43260 60800 43270 60840
rect 43378 60834 43578 60840
rect 43190 60790 43270 60800
rect 42660 59630 42730 60780
rect 42660 59370 42680 59630
rect 42720 59370 42730 59630
rect 43740 60780 43750 61020
rect 43790 60780 43810 61020
rect 43740 59630 43810 60780
rect 43190 59600 43270 59610
rect 42880 59562 43080 59568
rect 42770 59530 42850 59550
rect 42770 59470 42780 59530
rect 42840 59518 42850 59530
rect 42880 59528 42892 59562
rect 43068 59560 43080 59562
rect 43190 59560 43200 59600
rect 43068 59540 43200 59560
rect 43260 59560 43270 59600
rect 43378 59562 43578 59568
rect 43378 59560 43390 59562
rect 43260 59540 43390 59560
rect 43068 59530 43390 59540
rect 43068 59528 43080 59530
rect 42880 59522 43080 59528
rect 43378 59528 43390 59530
rect 43566 59528 43578 59562
rect 43378 59522 43578 59528
rect 43610 59530 43690 59550
rect 42842 59484 42850 59518
rect 42840 59470 42850 59484
rect 42770 59450 42850 59470
rect 42880 59474 43080 59480
rect 42880 59440 42892 59474
rect 43068 59470 43080 59474
rect 43378 59474 43578 59480
rect 43378 59470 43390 59474
rect 43068 59440 43390 59470
rect 43566 59440 43578 59474
rect 43610 59470 43620 59530
rect 43680 59470 43690 59530
rect 43610 59450 43690 59470
rect 42880 59434 43080 59440
rect 42660 59310 42730 59370
rect 42660 59070 42680 59310
rect 42720 59070 42730 59310
rect 43190 59430 43270 59440
rect 43378 59434 43578 59440
rect 43190 59370 43200 59430
rect 43260 59370 43270 59430
rect 43190 59320 43270 59370
rect 43190 59260 43200 59320
rect 43260 59260 43270 59320
rect 42880 59252 43080 59258
rect 42770 59220 42850 59240
rect 42770 59160 42780 59220
rect 42840 59208 42850 59220
rect 42880 59218 42892 59252
rect 43068 59250 43080 59252
rect 43190 59250 43270 59260
rect 43740 59390 43750 59630
rect 43790 59390 43810 59630
rect 43740 59310 43810 59390
rect 43378 59252 43578 59258
rect 43378 59250 43390 59252
rect 43068 59220 43390 59250
rect 43068 59218 43080 59220
rect 42880 59212 43080 59218
rect 43378 59218 43390 59220
rect 43566 59218 43578 59252
rect 43378 59212 43578 59218
rect 43610 59220 43690 59240
rect 42842 59174 42850 59208
rect 42840 59160 42850 59174
rect 42770 59140 42850 59160
rect 42880 59164 43080 59170
rect 42880 59130 42892 59164
rect 43068 59160 43080 59164
rect 43378 59164 43578 59170
rect 43378 59160 43390 59164
rect 43068 59150 43390 59160
rect 43068 59130 43200 59150
rect 42880 59124 43080 59130
rect 43190 59090 43200 59130
rect 43260 59130 43390 59150
rect 43566 59130 43578 59164
rect 43610 59160 43620 59220
rect 43680 59160 43690 59220
rect 43610 59140 43690 59160
rect 43260 59090 43270 59130
rect 43378 59124 43578 59130
rect 43190 59080 43270 59090
rect 42660 57920 42730 59070
rect 42660 57660 42680 57920
rect 42720 57660 42730 57920
rect 43740 59070 43750 59310
rect 43790 59070 43810 59310
rect 43740 57920 43810 59070
rect 43190 57890 43270 57900
rect 42880 57852 43080 57858
rect 42770 57820 42850 57840
rect 42770 57760 42780 57820
rect 42840 57808 42850 57820
rect 42880 57818 42892 57852
rect 43068 57850 43080 57852
rect 43190 57850 43200 57890
rect 43068 57830 43200 57850
rect 43260 57850 43270 57890
rect 43378 57852 43578 57858
rect 43378 57850 43390 57852
rect 43260 57830 43390 57850
rect 43068 57820 43390 57830
rect 43068 57818 43080 57820
rect 42880 57812 43080 57818
rect 43378 57818 43390 57820
rect 43566 57818 43578 57852
rect 43378 57812 43578 57818
rect 43610 57820 43690 57840
rect 42842 57774 42850 57808
rect 42840 57760 42850 57774
rect 42770 57740 42850 57760
rect 42880 57764 43080 57770
rect 42880 57730 42892 57764
rect 43068 57760 43080 57764
rect 43378 57764 43578 57770
rect 43378 57760 43390 57764
rect 43068 57730 43390 57760
rect 43566 57730 43578 57764
rect 43610 57760 43620 57820
rect 43680 57760 43690 57820
rect 43610 57740 43690 57760
rect 42880 57724 43080 57730
rect 42660 57600 42730 57660
rect 42660 57360 42680 57600
rect 42720 57360 42730 57600
rect 43190 57720 43270 57730
rect 43378 57724 43578 57730
rect 43190 57660 43200 57720
rect 43260 57660 43270 57720
rect 43190 57610 43270 57660
rect 43190 57550 43200 57610
rect 43260 57550 43270 57610
rect 42880 57542 43080 57548
rect 42770 57510 42850 57530
rect 42770 57450 42780 57510
rect 42840 57498 42850 57510
rect 42880 57508 42892 57542
rect 43068 57540 43080 57542
rect 43190 57540 43270 57550
rect 43740 57680 43750 57920
rect 43790 57680 43810 57920
rect 43740 57600 43810 57680
rect 43378 57542 43578 57548
rect 43378 57540 43390 57542
rect 43068 57510 43390 57540
rect 43068 57508 43080 57510
rect 42880 57502 43080 57508
rect 43378 57508 43390 57510
rect 43566 57508 43578 57542
rect 43378 57502 43578 57508
rect 43610 57510 43690 57530
rect 42842 57464 42850 57498
rect 42840 57450 42850 57464
rect 42770 57430 42850 57450
rect 42880 57454 43080 57460
rect 42880 57420 42892 57454
rect 43068 57450 43080 57454
rect 43378 57454 43578 57460
rect 43378 57450 43390 57454
rect 43068 57440 43390 57450
rect 43068 57420 43200 57440
rect 42880 57414 43080 57420
rect 43190 57380 43200 57420
rect 43260 57420 43390 57440
rect 43566 57420 43578 57454
rect 43610 57450 43620 57510
rect 43680 57450 43690 57510
rect 43610 57430 43690 57450
rect 43260 57380 43270 57420
rect 43378 57414 43578 57420
rect 43190 57370 43270 57380
rect 42660 56210 42730 57360
rect 42660 55950 42680 56210
rect 42720 55950 42730 56210
rect 43740 57360 43750 57600
rect 43790 57360 43810 57600
rect 43740 56210 43810 57360
rect 43190 56180 43270 56190
rect 42880 56142 43080 56148
rect 42770 56110 42850 56130
rect 42770 56050 42780 56110
rect 42840 56098 42850 56110
rect 42880 56108 42892 56142
rect 43068 56140 43080 56142
rect 43190 56140 43200 56180
rect 43068 56120 43200 56140
rect 43260 56140 43270 56180
rect 43378 56142 43578 56148
rect 43378 56140 43390 56142
rect 43260 56120 43390 56140
rect 43068 56110 43390 56120
rect 43068 56108 43080 56110
rect 42880 56102 43080 56108
rect 43378 56108 43390 56110
rect 43566 56108 43578 56142
rect 43378 56102 43578 56108
rect 43610 56110 43690 56130
rect 42842 56064 42850 56098
rect 42840 56050 42850 56064
rect 42770 56030 42850 56050
rect 42880 56054 43080 56060
rect 42880 56020 42892 56054
rect 43068 56050 43080 56054
rect 43378 56054 43578 56060
rect 43378 56050 43390 56054
rect 43068 56020 43390 56050
rect 43566 56020 43578 56054
rect 43610 56050 43620 56110
rect 43680 56050 43690 56110
rect 43610 56030 43690 56050
rect 42880 56014 43080 56020
rect 42660 55890 42730 55950
rect 42660 55650 42680 55890
rect 42720 55650 42730 55890
rect 43190 56010 43270 56020
rect 43378 56014 43578 56020
rect 43190 55950 43200 56010
rect 43260 55950 43270 56010
rect 43190 55900 43270 55950
rect 43190 55840 43200 55900
rect 43260 55840 43270 55900
rect 42880 55832 43080 55838
rect 42770 55800 42850 55820
rect 42770 55740 42780 55800
rect 42840 55788 42850 55800
rect 42880 55798 42892 55832
rect 43068 55830 43080 55832
rect 43190 55830 43270 55840
rect 43740 55970 43750 56210
rect 43790 55970 43810 56210
rect 43740 55890 43810 55970
rect 43378 55832 43578 55838
rect 43378 55830 43390 55832
rect 43068 55800 43390 55830
rect 43068 55798 43080 55800
rect 42880 55792 43080 55798
rect 43378 55798 43390 55800
rect 43566 55798 43578 55832
rect 43378 55792 43578 55798
rect 43610 55800 43690 55820
rect 42842 55754 42850 55788
rect 42840 55740 42850 55754
rect 42770 55720 42850 55740
rect 42880 55744 43080 55750
rect 42880 55710 42892 55744
rect 43068 55740 43080 55744
rect 43378 55744 43578 55750
rect 43378 55740 43390 55744
rect 43068 55730 43390 55740
rect 43068 55710 43200 55730
rect 42880 55704 43080 55710
rect 43190 55670 43200 55710
rect 43260 55710 43390 55730
rect 43566 55710 43578 55744
rect 43610 55740 43620 55800
rect 43680 55740 43690 55800
rect 43610 55720 43690 55740
rect 43260 55670 43270 55710
rect 43378 55704 43578 55710
rect 43190 55660 43270 55670
rect 42660 54500 42730 55650
rect 42660 54240 42680 54500
rect 42720 54240 42730 54500
rect 43740 55650 43750 55890
rect 43790 55650 43810 55890
rect 43740 54500 43810 55650
rect 43190 54470 43270 54480
rect 42880 54432 43080 54438
rect 42770 54400 42850 54420
rect 42770 54340 42780 54400
rect 42840 54388 42850 54400
rect 42880 54398 42892 54432
rect 43068 54430 43080 54432
rect 43190 54430 43200 54470
rect 43068 54410 43200 54430
rect 43260 54430 43270 54470
rect 43378 54432 43578 54438
rect 43378 54430 43390 54432
rect 43260 54410 43390 54430
rect 43068 54400 43390 54410
rect 43068 54398 43080 54400
rect 42880 54392 43080 54398
rect 43378 54398 43390 54400
rect 43566 54398 43578 54432
rect 43378 54392 43578 54398
rect 43610 54400 43690 54420
rect 42842 54354 42850 54388
rect 42840 54340 42850 54354
rect 42770 54320 42850 54340
rect 42880 54344 43080 54350
rect 42880 54310 42892 54344
rect 43068 54340 43080 54344
rect 43378 54344 43578 54350
rect 43378 54340 43390 54344
rect 43068 54310 43390 54340
rect 43566 54310 43578 54344
rect 43610 54340 43620 54400
rect 43680 54340 43690 54400
rect 43610 54320 43690 54340
rect 42880 54304 43080 54310
rect 42660 54180 42730 54240
rect 42660 53940 42680 54180
rect 42720 53940 42730 54180
rect 43190 54300 43270 54310
rect 43378 54304 43578 54310
rect 43190 54240 43200 54300
rect 43260 54240 43270 54300
rect 43190 54190 43270 54240
rect 43190 54130 43200 54190
rect 43260 54130 43270 54190
rect 42880 54122 43080 54128
rect 42770 54090 42850 54110
rect 42770 54030 42780 54090
rect 42840 54078 42850 54090
rect 42880 54088 42892 54122
rect 43068 54120 43080 54122
rect 43190 54120 43270 54130
rect 43740 54260 43750 54500
rect 43790 54260 43810 54500
rect 43740 54180 43810 54260
rect 43378 54122 43578 54128
rect 43378 54120 43390 54122
rect 43068 54090 43390 54120
rect 43068 54088 43080 54090
rect 42880 54082 43080 54088
rect 43378 54088 43390 54090
rect 43566 54088 43578 54122
rect 43378 54082 43578 54088
rect 43610 54090 43690 54110
rect 42842 54044 42850 54078
rect 42840 54030 42850 54044
rect 42770 54010 42850 54030
rect 42880 54034 43080 54040
rect 42880 54000 42892 54034
rect 43068 54030 43080 54034
rect 43378 54034 43578 54040
rect 43378 54030 43390 54034
rect 43068 54020 43390 54030
rect 43068 54000 43200 54020
rect 42880 53994 43080 54000
rect 43190 53960 43200 54000
rect 43260 54000 43390 54020
rect 43566 54000 43578 54034
rect 43610 54030 43620 54090
rect 43680 54030 43690 54090
rect 43610 54010 43690 54030
rect 43260 53960 43270 54000
rect 43378 53994 43578 54000
rect 43190 53950 43270 53960
rect 42660 52790 42730 53940
rect 42660 52530 42680 52790
rect 42720 52530 42730 52790
rect 43740 53940 43750 54180
rect 43790 53940 43810 54180
rect 43740 52790 43810 53940
rect 43190 52760 43270 52770
rect 42880 52722 43080 52728
rect 42770 52690 42850 52710
rect 42770 52630 42780 52690
rect 42840 52678 42850 52690
rect 42880 52688 42892 52722
rect 43068 52720 43080 52722
rect 43190 52720 43200 52760
rect 43068 52700 43200 52720
rect 43260 52720 43270 52760
rect 43378 52722 43578 52728
rect 43378 52720 43390 52722
rect 43260 52700 43390 52720
rect 43068 52690 43390 52700
rect 43068 52688 43080 52690
rect 42880 52682 43080 52688
rect 43378 52688 43390 52690
rect 43566 52688 43578 52722
rect 43378 52682 43578 52688
rect 43610 52690 43690 52710
rect 42842 52644 42850 52678
rect 42840 52630 42850 52644
rect 42770 52610 42850 52630
rect 42880 52634 43080 52640
rect 42880 52600 42892 52634
rect 43068 52630 43080 52634
rect 43378 52634 43578 52640
rect 43378 52630 43390 52634
rect 43068 52600 43390 52630
rect 43566 52600 43578 52634
rect 43610 52630 43620 52690
rect 43680 52630 43690 52690
rect 43610 52610 43690 52630
rect 42880 52594 43080 52600
rect 42660 52470 42730 52530
rect 42660 52230 42680 52470
rect 42720 52230 42730 52470
rect 43190 52590 43270 52600
rect 43378 52594 43578 52600
rect 43190 52530 43200 52590
rect 43260 52530 43270 52590
rect 43190 52480 43270 52530
rect 43190 52420 43200 52480
rect 43260 52420 43270 52480
rect 42880 52412 43080 52418
rect 42770 52380 42850 52400
rect 42770 52320 42780 52380
rect 42840 52368 42850 52380
rect 42880 52378 42892 52412
rect 43068 52410 43080 52412
rect 43190 52410 43270 52420
rect 43740 52550 43750 52790
rect 43790 52550 43810 52790
rect 43740 52470 43810 52550
rect 43378 52412 43578 52418
rect 43378 52410 43390 52412
rect 43068 52380 43390 52410
rect 43068 52378 43080 52380
rect 42880 52372 43080 52378
rect 43378 52378 43390 52380
rect 43566 52378 43578 52412
rect 43378 52372 43578 52378
rect 43610 52380 43690 52400
rect 42842 52334 42850 52368
rect 42840 52320 42850 52334
rect 42770 52300 42850 52320
rect 42880 52324 43080 52330
rect 42880 52290 42892 52324
rect 43068 52320 43080 52324
rect 43378 52324 43578 52330
rect 43378 52320 43390 52324
rect 43068 52310 43390 52320
rect 43068 52290 43200 52310
rect 42880 52284 43080 52290
rect 43190 52250 43200 52290
rect 43260 52290 43390 52310
rect 43566 52290 43578 52324
rect 43610 52320 43620 52380
rect 43680 52320 43690 52380
rect 43610 52300 43690 52320
rect 43260 52250 43270 52290
rect 43378 52284 43578 52290
rect 43190 52240 43270 52250
rect 42660 51080 42730 52230
rect 42660 50820 42680 51080
rect 42720 50820 42730 51080
rect 43740 52230 43750 52470
rect 43790 52230 43810 52470
rect 43740 51080 43810 52230
rect 43190 51050 43270 51060
rect 42880 51012 43080 51018
rect 42770 50980 42850 51000
rect 42770 50920 42780 50980
rect 42840 50968 42850 50980
rect 42880 50978 42892 51012
rect 43068 51010 43080 51012
rect 43190 51010 43200 51050
rect 43068 50990 43200 51010
rect 43260 51010 43270 51050
rect 43378 51012 43578 51018
rect 43378 51010 43390 51012
rect 43260 50990 43390 51010
rect 43068 50980 43390 50990
rect 43068 50978 43080 50980
rect 42880 50972 43080 50978
rect 43378 50978 43390 50980
rect 43566 50978 43578 51012
rect 43378 50972 43578 50978
rect 43610 50980 43690 51000
rect 42842 50934 42850 50968
rect 42840 50920 42850 50934
rect 42770 50900 42850 50920
rect 42880 50924 43080 50930
rect 42880 50890 42892 50924
rect 43068 50920 43080 50924
rect 43378 50924 43578 50930
rect 43378 50920 43390 50924
rect 43068 50890 43390 50920
rect 43566 50890 43578 50924
rect 43610 50920 43620 50980
rect 43680 50920 43690 50980
rect 43610 50900 43690 50920
rect 42880 50884 43080 50890
rect 42660 50760 42730 50820
rect 42660 50520 42680 50760
rect 42720 50520 42730 50760
rect 43190 50880 43270 50890
rect 43378 50884 43578 50890
rect 43190 50820 43200 50880
rect 43260 50820 43270 50880
rect 43190 50770 43270 50820
rect 43190 50710 43200 50770
rect 43260 50710 43270 50770
rect 42880 50702 43080 50708
rect 42770 50670 42850 50690
rect 42770 50610 42780 50670
rect 42840 50658 42850 50670
rect 42880 50668 42892 50702
rect 43068 50700 43080 50702
rect 43190 50700 43270 50710
rect 43740 50840 43750 51080
rect 43790 50840 43810 51080
rect 43740 50760 43810 50840
rect 43378 50702 43578 50708
rect 43378 50700 43390 50702
rect 43068 50670 43390 50700
rect 43068 50668 43080 50670
rect 42880 50662 43080 50668
rect 43378 50668 43390 50670
rect 43566 50668 43578 50702
rect 43378 50662 43578 50668
rect 43610 50670 43690 50690
rect 42842 50624 42850 50658
rect 42840 50610 42850 50624
rect 42770 50590 42850 50610
rect 42880 50614 43080 50620
rect 42880 50580 42892 50614
rect 43068 50610 43080 50614
rect 43378 50614 43578 50620
rect 43378 50610 43390 50614
rect 43068 50600 43390 50610
rect 43068 50580 43200 50600
rect 42880 50574 43080 50580
rect 43190 50540 43200 50580
rect 43260 50580 43390 50600
rect 43566 50580 43578 50614
rect 43610 50610 43620 50670
rect 43680 50610 43690 50670
rect 43610 50590 43690 50610
rect 43260 50540 43270 50580
rect 43378 50574 43578 50580
rect 43190 50530 43270 50540
rect 42660 49370 42730 50520
rect 42660 49110 42680 49370
rect 42720 49110 42730 49370
rect 43740 50520 43750 50760
rect 43790 50520 43810 50760
rect 43740 49370 43810 50520
rect 43190 49340 43270 49350
rect 42880 49302 43080 49308
rect 42770 49270 42850 49290
rect 42770 49210 42780 49270
rect 42840 49258 42850 49270
rect 42880 49268 42892 49302
rect 43068 49300 43080 49302
rect 43190 49300 43200 49340
rect 43068 49280 43200 49300
rect 43260 49300 43270 49340
rect 43378 49302 43578 49308
rect 43378 49300 43390 49302
rect 43260 49280 43390 49300
rect 43068 49270 43390 49280
rect 43068 49268 43080 49270
rect 42880 49262 43080 49268
rect 43378 49268 43390 49270
rect 43566 49268 43578 49302
rect 43378 49262 43578 49268
rect 43610 49270 43690 49290
rect 42842 49224 42850 49258
rect 42840 49210 42850 49224
rect 42770 49190 42850 49210
rect 42880 49214 43080 49220
rect 42880 49180 42892 49214
rect 43068 49210 43080 49214
rect 43378 49214 43578 49220
rect 43378 49210 43390 49214
rect 43068 49180 43390 49210
rect 43566 49180 43578 49214
rect 43610 49210 43620 49270
rect 43680 49210 43690 49270
rect 43610 49190 43690 49210
rect 42880 49174 43080 49180
rect 42660 49050 42730 49110
rect 42660 48810 42680 49050
rect 42720 48810 42730 49050
rect 43190 49170 43270 49180
rect 43378 49174 43578 49180
rect 43190 49110 43200 49170
rect 43260 49110 43270 49170
rect 43190 49060 43270 49110
rect 43190 49000 43200 49060
rect 43260 49000 43270 49060
rect 42880 48992 43080 48998
rect 42770 48960 42850 48980
rect 42770 48900 42780 48960
rect 42840 48948 42850 48960
rect 42880 48958 42892 48992
rect 43068 48990 43080 48992
rect 43190 48990 43270 49000
rect 43740 49130 43750 49370
rect 43790 49130 43810 49370
rect 43740 49050 43810 49130
rect 43378 48992 43578 48998
rect 43378 48990 43390 48992
rect 43068 48960 43390 48990
rect 43068 48958 43080 48960
rect 42880 48952 43080 48958
rect 43378 48958 43390 48960
rect 43566 48958 43578 48992
rect 43378 48952 43578 48958
rect 43610 48960 43690 48980
rect 42842 48914 42850 48948
rect 42840 48900 42850 48914
rect 42770 48880 42850 48900
rect 42880 48904 43080 48910
rect 42880 48870 42892 48904
rect 43068 48900 43080 48904
rect 43378 48904 43578 48910
rect 43378 48900 43390 48904
rect 43068 48890 43390 48900
rect 43068 48870 43200 48890
rect 42880 48864 43080 48870
rect 43190 48830 43200 48870
rect 43260 48870 43390 48890
rect 43566 48870 43578 48904
rect 43610 48900 43620 48960
rect 43680 48900 43690 48960
rect 43610 48880 43690 48900
rect 43260 48830 43270 48870
rect 43378 48864 43578 48870
rect 43190 48820 43270 48830
rect 42660 47660 42730 48810
rect 42660 47400 42680 47660
rect 42720 47400 42730 47660
rect 43740 48810 43750 49050
rect 43790 48810 43810 49050
rect 43740 47660 43810 48810
rect 43190 47630 43270 47640
rect 42880 47592 43080 47598
rect 42770 47560 42850 47580
rect 42770 47500 42780 47560
rect 42840 47548 42850 47560
rect 42880 47558 42892 47592
rect 43068 47590 43080 47592
rect 43190 47590 43200 47630
rect 43068 47570 43200 47590
rect 43260 47590 43270 47630
rect 43378 47592 43578 47598
rect 43378 47590 43390 47592
rect 43260 47570 43390 47590
rect 43068 47560 43390 47570
rect 43068 47558 43080 47560
rect 42880 47552 43080 47558
rect 43378 47558 43390 47560
rect 43566 47558 43578 47592
rect 43378 47552 43578 47558
rect 43610 47560 43690 47580
rect 42842 47514 42850 47548
rect 42840 47500 42850 47514
rect 42770 47480 42850 47500
rect 42880 47504 43080 47510
rect 42880 47470 42892 47504
rect 43068 47500 43080 47504
rect 43378 47504 43578 47510
rect 43378 47500 43390 47504
rect 43068 47470 43390 47500
rect 43566 47470 43578 47504
rect 43610 47500 43620 47560
rect 43680 47500 43690 47560
rect 43610 47480 43690 47500
rect 42880 47464 43080 47470
rect 42660 47340 42730 47400
rect 42660 47100 42680 47340
rect 42720 47100 42730 47340
rect 43190 47460 43270 47470
rect 43378 47464 43578 47470
rect 43190 47400 43200 47460
rect 43260 47400 43270 47460
rect 43190 47350 43270 47400
rect 43190 47290 43200 47350
rect 43260 47290 43270 47350
rect 42880 47282 43080 47288
rect 42770 47250 42850 47270
rect 42770 47190 42780 47250
rect 42840 47238 42850 47250
rect 42880 47248 42892 47282
rect 43068 47280 43080 47282
rect 43190 47280 43270 47290
rect 43740 47420 43750 47660
rect 43790 47420 43810 47660
rect 43740 47340 43810 47420
rect 43378 47282 43578 47288
rect 43378 47280 43390 47282
rect 43068 47250 43390 47280
rect 43068 47248 43080 47250
rect 42880 47242 43080 47248
rect 43378 47248 43390 47250
rect 43566 47248 43578 47282
rect 43378 47242 43578 47248
rect 43610 47250 43690 47270
rect 42842 47204 42850 47238
rect 42840 47190 42850 47204
rect 42770 47170 42850 47190
rect 42880 47194 43080 47200
rect 42880 47160 42892 47194
rect 43068 47190 43080 47194
rect 43378 47194 43578 47200
rect 43378 47190 43390 47194
rect 43068 47180 43390 47190
rect 43068 47160 43200 47180
rect 42880 47154 43080 47160
rect 43190 47120 43200 47160
rect 43260 47160 43390 47180
rect 43566 47160 43578 47194
rect 43610 47190 43620 47250
rect 43680 47190 43690 47250
rect 43610 47170 43690 47190
rect 43260 47120 43270 47160
rect 43378 47154 43578 47160
rect 43190 47110 43270 47120
rect 42660 45950 42730 47100
rect 42660 45690 42680 45950
rect 42720 45690 42730 45950
rect 43740 47100 43750 47340
rect 43790 47100 43810 47340
rect 43740 45950 43810 47100
rect 43190 45920 43270 45930
rect 42880 45882 43080 45888
rect 42770 45850 42850 45870
rect 42770 45790 42780 45850
rect 42840 45838 42850 45850
rect 42880 45848 42892 45882
rect 43068 45880 43080 45882
rect 43190 45880 43200 45920
rect 43068 45860 43200 45880
rect 43260 45880 43270 45920
rect 43378 45882 43578 45888
rect 43378 45880 43390 45882
rect 43260 45860 43390 45880
rect 43068 45850 43390 45860
rect 43068 45848 43080 45850
rect 42880 45842 43080 45848
rect 43378 45848 43390 45850
rect 43566 45848 43578 45882
rect 43378 45842 43578 45848
rect 43610 45850 43690 45870
rect 42842 45804 42850 45838
rect 42840 45790 42850 45804
rect 42770 45770 42850 45790
rect 42880 45794 43080 45800
rect 42880 45760 42892 45794
rect 43068 45790 43080 45794
rect 43378 45794 43578 45800
rect 43378 45790 43390 45794
rect 43068 45760 43390 45790
rect 43566 45760 43578 45794
rect 43610 45790 43620 45850
rect 43680 45790 43690 45850
rect 43610 45770 43690 45790
rect 42880 45754 43080 45760
rect 42660 45630 42730 45690
rect 42660 45390 42680 45630
rect 42720 45390 42730 45630
rect 43190 45750 43270 45760
rect 43378 45754 43578 45760
rect 43190 45690 43200 45750
rect 43260 45690 43270 45750
rect 43190 45640 43270 45690
rect 43190 45580 43200 45640
rect 43260 45580 43270 45640
rect 42880 45572 43080 45578
rect 42770 45540 42850 45560
rect 42770 45480 42780 45540
rect 42840 45528 42850 45540
rect 42880 45538 42892 45572
rect 43068 45570 43080 45572
rect 43190 45570 43270 45580
rect 43740 45710 43750 45950
rect 43790 45710 43810 45950
rect 43740 45630 43810 45710
rect 43378 45572 43578 45578
rect 43378 45570 43390 45572
rect 43068 45540 43390 45570
rect 43068 45538 43080 45540
rect 42880 45532 43080 45538
rect 43378 45538 43390 45540
rect 43566 45538 43578 45572
rect 43378 45532 43578 45538
rect 43610 45540 43690 45560
rect 42842 45494 42850 45528
rect 42840 45480 42850 45494
rect 42770 45460 42850 45480
rect 42880 45484 43080 45490
rect 42880 45450 42892 45484
rect 43068 45480 43080 45484
rect 43378 45484 43578 45490
rect 43378 45480 43390 45484
rect 43068 45470 43390 45480
rect 43068 45450 43200 45470
rect 42880 45444 43080 45450
rect 43190 45410 43200 45450
rect 43260 45450 43390 45470
rect 43566 45450 43578 45484
rect 43610 45480 43620 45540
rect 43680 45480 43690 45540
rect 43610 45460 43690 45480
rect 43260 45410 43270 45450
rect 43378 45444 43578 45450
rect 43190 45400 43270 45410
rect 42660 44240 42730 45390
rect 42660 43980 42680 44240
rect 42720 43980 42730 44240
rect 43740 45390 43750 45630
rect 43790 45390 43810 45630
rect 43740 44240 43810 45390
rect 43190 44210 43270 44220
rect 42880 44172 43080 44178
rect 42770 44140 42850 44160
rect 42770 44080 42780 44140
rect 42840 44128 42850 44140
rect 42880 44138 42892 44172
rect 43068 44170 43080 44172
rect 43190 44170 43200 44210
rect 43068 44150 43200 44170
rect 43260 44170 43270 44210
rect 43378 44172 43578 44178
rect 43378 44170 43390 44172
rect 43260 44150 43390 44170
rect 43068 44140 43390 44150
rect 43068 44138 43080 44140
rect 42880 44132 43080 44138
rect 43378 44138 43390 44140
rect 43566 44138 43578 44172
rect 43378 44132 43578 44138
rect 43610 44140 43690 44160
rect 42842 44094 42850 44128
rect 42840 44080 42850 44094
rect 42770 44060 42850 44080
rect 42880 44084 43080 44090
rect 42880 44050 42892 44084
rect 43068 44080 43080 44084
rect 43378 44084 43578 44090
rect 43378 44080 43390 44084
rect 43068 44050 43390 44080
rect 43566 44050 43578 44084
rect 43610 44080 43620 44140
rect 43680 44080 43690 44140
rect 43610 44060 43690 44080
rect 42880 44044 43080 44050
rect 42660 43920 42730 43980
rect 42660 43680 42680 43920
rect 42720 43680 42730 43920
rect 43190 44040 43270 44050
rect 43378 44044 43578 44050
rect 43190 43980 43200 44040
rect 43260 43980 43270 44040
rect 43190 43930 43270 43980
rect 43190 43870 43200 43930
rect 43260 43870 43270 43930
rect 42880 43862 43080 43868
rect 42770 43830 42850 43850
rect 42770 43770 42780 43830
rect 42840 43818 42850 43830
rect 42880 43828 42892 43862
rect 43068 43860 43080 43862
rect 43190 43860 43270 43870
rect 43740 44000 43750 44240
rect 43790 44000 43810 44240
rect 43740 43920 43810 44000
rect 43378 43862 43578 43868
rect 43378 43860 43390 43862
rect 43068 43830 43390 43860
rect 43068 43828 43080 43830
rect 42880 43822 43080 43828
rect 43378 43828 43390 43830
rect 43566 43828 43578 43862
rect 43378 43822 43578 43828
rect 43610 43830 43690 43850
rect 42842 43784 42850 43818
rect 42840 43770 42850 43784
rect 42770 43750 42850 43770
rect 42880 43774 43080 43780
rect 42880 43740 42892 43774
rect 43068 43770 43080 43774
rect 43378 43774 43578 43780
rect 43378 43770 43390 43774
rect 43068 43760 43390 43770
rect 43068 43740 43200 43760
rect 42880 43734 43080 43740
rect 43190 43700 43200 43740
rect 43260 43740 43390 43760
rect 43566 43740 43578 43774
rect 43610 43770 43620 43830
rect 43680 43770 43690 43830
rect 43610 43750 43690 43770
rect 43260 43700 43270 43740
rect 43378 43734 43578 43740
rect 43190 43690 43270 43700
rect 42660 42530 42730 43680
rect 42660 42270 42680 42530
rect 42720 42270 42730 42530
rect 43740 43680 43750 43920
rect 43790 43680 43810 43920
rect 43740 42530 43810 43680
rect 43190 42500 43270 42510
rect 42880 42462 43080 42468
rect 42770 42430 42850 42450
rect 42770 42370 42780 42430
rect 42840 42418 42850 42430
rect 42880 42428 42892 42462
rect 43068 42460 43080 42462
rect 43190 42460 43200 42500
rect 43068 42440 43200 42460
rect 43260 42460 43270 42500
rect 43378 42462 43578 42468
rect 43378 42460 43390 42462
rect 43260 42440 43390 42460
rect 43068 42430 43390 42440
rect 43068 42428 43080 42430
rect 42880 42422 43080 42428
rect 43378 42428 43390 42430
rect 43566 42428 43578 42462
rect 43378 42422 43578 42428
rect 43610 42430 43690 42450
rect 42842 42384 42850 42418
rect 42840 42370 42850 42384
rect 42770 42350 42850 42370
rect 42880 42374 43080 42380
rect 42880 42340 42892 42374
rect 43068 42370 43080 42374
rect 43378 42374 43578 42380
rect 43378 42370 43390 42374
rect 43068 42340 43390 42370
rect 43566 42340 43578 42374
rect 43610 42370 43620 42430
rect 43680 42370 43690 42430
rect 43610 42350 43690 42370
rect 42880 42334 43080 42340
rect 42660 42210 42730 42270
rect 42660 41970 42680 42210
rect 42720 41970 42730 42210
rect 43190 42330 43270 42340
rect 43378 42334 43578 42340
rect 43190 42270 43200 42330
rect 43260 42270 43270 42330
rect 43190 42220 43270 42270
rect 43190 42160 43200 42220
rect 43260 42160 43270 42220
rect 42880 42152 43080 42158
rect 42770 42120 42850 42140
rect 42770 42060 42780 42120
rect 42840 42108 42850 42120
rect 42880 42118 42892 42152
rect 43068 42150 43080 42152
rect 43190 42150 43270 42160
rect 43740 42290 43750 42530
rect 43790 42290 43810 42530
rect 43740 42210 43810 42290
rect 43378 42152 43578 42158
rect 43378 42150 43390 42152
rect 43068 42120 43390 42150
rect 43068 42118 43080 42120
rect 42880 42112 43080 42118
rect 43378 42118 43390 42120
rect 43566 42118 43578 42152
rect 43378 42112 43578 42118
rect 43610 42120 43690 42140
rect 42842 42074 42850 42108
rect 42840 42060 42850 42074
rect 42770 42040 42850 42060
rect 42880 42064 43080 42070
rect 42880 42030 42892 42064
rect 43068 42060 43080 42064
rect 43378 42064 43578 42070
rect 43378 42060 43390 42064
rect 43068 42050 43390 42060
rect 43068 42030 43200 42050
rect 42880 42024 43080 42030
rect 43190 41990 43200 42030
rect 43260 42030 43390 42050
rect 43566 42030 43578 42064
rect 43610 42060 43620 42120
rect 43680 42060 43690 42120
rect 43610 42040 43690 42060
rect 43260 41990 43270 42030
rect 43378 42024 43578 42030
rect 43190 41980 43270 41990
rect 42660 40820 42730 41970
rect 42660 40560 42680 40820
rect 42720 40560 42730 40820
rect 43740 41970 43750 42210
rect 43790 41970 43810 42210
rect 43740 40820 43810 41970
rect 43190 40790 43270 40800
rect 42880 40752 43080 40758
rect 42770 40720 42850 40740
rect 42770 40660 42780 40720
rect 42840 40708 42850 40720
rect 42880 40718 42892 40752
rect 43068 40750 43080 40752
rect 43190 40750 43200 40790
rect 43068 40730 43200 40750
rect 43260 40750 43270 40790
rect 43378 40752 43578 40758
rect 43378 40750 43390 40752
rect 43260 40730 43390 40750
rect 43068 40720 43390 40730
rect 43068 40718 43080 40720
rect 42880 40712 43080 40718
rect 43378 40718 43390 40720
rect 43566 40718 43578 40752
rect 43378 40712 43578 40718
rect 43610 40720 43690 40740
rect 42842 40674 42850 40708
rect 42840 40660 42850 40674
rect 42770 40640 42850 40660
rect 42880 40664 43080 40670
rect 42880 40630 42892 40664
rect 43068 40660 43080 40664
rect 43378 40664 43578 40670
rect 43378 40660 43390 40664
rect 43068 40630 43390 40660
rect 43566 40630 43578 40664
rect 43610 40660 43620 40720
rect 43680 40660 43690 40720
rect 43610 40640 43690 40660
rect 42880 40624 43080 40630
rect 42660 40500 42730 40560
rect 42660 40260 42680 40500
rect 42720 40260 42730 40500
rect 43190 40620 43270 40630
rect 43378 40624 43578 40630
rect 43190 40560 43200 40620
rect 43260 40560 43270 40620
rect 43190 40510 43270 40560
rect 43190 40450 43200 40510
rect 43260 40450 43270 40510
rect 42880 40442 43080 40448
rect 42770 40410 42850 40430
rect 42770 40350 42780 40410
rect 42840 40398 42850 40410
rect 42880 40408 42892 40442
rect 43068 40440 43080 40442
rect 43190 40440 43270 40450
rect 43740 40580 43750 40820
rect 43790 40580 43810 40820
rect 43740 40500 43810 40580
rect 43378 40442 43578 40448
rect 43378 40440 43390 40442
rect 43068 40410 43390 40440
rect 43068 40408 43080 40410
rect 42880 40402 43080 40408
rect 43378 40408 43390 40410
rect 43566 40408 43578 40442
rect 43378 40402 43578 40408
rect 43610 40410 43690 40430
rect 42842 40364 42850 40398
rect 42840 40350 42850 40364
rect 42770 40330 42850 40350
rect 42880 40354 43080 40360
rect 42880 40320 42892 40354
rect 43068 40350 43080 40354
rect 43378 40354 43578 40360
rect 43378 40350 43390 40354
rect 43068 40340 43390 40350
rect 43068 40320 43200 40340
rect 42880 40314 43080 40320
rect 43190 40280 43200 40320
rect 43260 40320 43390 40340
rect 43566 40320 43578 40354
rect 43610 40350 43620 40410
rect 43680 40350 43690 40410
rect 43610 40330 43690 40350
rect 43260 40280 43270 40320
rect 43378 40314 43578 40320
rect 43190 40270 43270 40280
rect 42660 39690 42730 40260
rect 43740 40260 43750 40500
rect 43790 40260 43810 40500
rect 43740 39690 43810 40260
rect 42660 39680 42740 39690
rect 42660 39620 42670 39680
rect 42730 39620 42740 39680
rect 43730 39680 43810 39690
rect 43730 39620 43740 39680
rect 43800 39620 43810 39680
rect 43730 39610 43810 39620
rect 43840 66480 43870 67050
rect 43840 66470 43900 66480
rect 43840 66400 43900 66410
rect 43840 64770 43870 66400
rect 43930 65950 43960 67050
rect 43900 65940 43960 65950
rect 43900 65870 43960 65880
rect 43840 64760 43900 64770
rect 43840 64690 43900 64700
rect 43840 63060 43870 64690
rect 43930 64240 43960 65870
rect 43900 64230 43960 64240
rect 43900 64160 43960 64170
rect 43840 63050 43900 63060
rect 43840 62980 43900 62990
rect 43840 61350 43870 62980
rect 43930 62530 43960 64160
rect 43900 62520 43960 62530
rect 43900 62450 43960 62460
rect 43840 61340 43900 61350
rect 43840 61270 43900 61280
rect 43840 59640 43870 61270
rect 43930 60820 43960 62450
rect 43900 60810 43960 60820
rect 43900 60740 43960 60750
rect 43840 59630 43900 59640
rect 43840 59560 43900 59570
rect 43840 57930 43870 59560
rect 43930 59110 43960 60740
rect 43900 59100 43960 59110
rect 43900 59030 43960 59040
rect 43840 57920 43900 57930
rect 43840 57850 43900 57860
rect 43840 56220 43870 57850
rect 43930 57400 43960 59030
rect 43900 57390 43960 57400
rect 43900 57320 43960 57330
rect 43840 56210 43900 56220
rect 43840 56140 43900 56150
rect 43840 54510 43870 56140
rect 43930 55690 43960 57320
rect 43900 55680 43960 55690
rect 43900 55610 43960 55620
rect 43840 54500 43900 54510
rect 43840 54430 43900 54440
rect 43840 52800 43870 54430
rect 43930 53980 43960 55610
rect 43900 53970 43960 53980
rect 43900 53900 43960 53910
rect 43840 52790 43900 52800
rect 43840 52720 43900 52730
rect 43840 51090 43870 52720
rect 43930 52270 43960 53900
rect 43900 52260 43960 52270
rect 43900 52190 43960 52200
rect 43840 51080 43900 51090
rect 43840 51010 43900 51020
rect 43840 49380 43870 51010
rect 43930 50560 43960 52190
rect 43900 50550 43960 50560
rect 43900 50480 43960 50490
rect 43840 49370 43900 49380
rect 43840 49300 43900 49310
rect 43840 47670 43870 49300
rect 43930 48850 43960 50480
rect 43900 48840 43960 48850
rect 43900 48770 43960 48780
rect 43840 47660 43900 47670
rect 43840 47590 43900 47600
rect 43840 45960 43870 47590
rect 43930 47140 43960 48770
rect 43900 47130 43960 47140
rect 43900 47060 43960 47070
rect 43840 45950 43900 45960
rect 43840 45880 43900 45890
rect 43840 44250 43870 45880
rect 43930 45430 43960 47060
rect 43900 45420 43960 45430
rect 43900 45350 43960 45360
rect 43840 44240 43900 44250
rect 43840 44170 43900 44180
rect 43840 42540 43870 44170
rect 43930 43720 43960 45350
rect 43900 43710 43960 43720
rect 43900 43640 43960 43650
rect 43840 42530 43900 42540
rect 43840 42460 43900 42470
rect 43840 40830 43870 42460
rect 43930 42010 43960 43640
rect 43900 42000 43960 42010
rect 43900 41930 43960 41940
rect 43840 40820 43900 40830
rect 43840 40750 43900 40760
rect 42190 39220 42250 39230
rect 42370 39230 42630 39240
rect 39200 39160 39260 39170
rect 42430 39210 42630 39230
rect 42370 39160 42430 39170
rect 43840 38840 43870 40750
rect 43930 40300 43960 41930
rect 43900 40290 43960 40300
rect 43900 40220 43960 40230
rect 43930 39690 43960 40220
rect 43900 39680 43960 39690
rect 43900 39610 43960 39620
rect 43990 66390 44020 67050
rect 43990 66380 44050 66390
rect 43990 66310 44050 66320
rect 43990 64680 44020 66310
rect 43990 64670 44050 64680
rect 43990 64600 44050 64610
rect 43990 42440 44020 64600
rect 44110 62970 44140 67050
rect 44110 62960 44170 62970
rect 44110 62890 44170 62900
rect 44110 61260 44140 62890
rect 44110 61250 44170 61260
rect 44110 61180 44170 61190
rect 44110 45870 44140 61180
rect 44230 59550 44260 67050
rect 44230 59540 44290 59550
rect 44230 59470 44290 59480
rect 44230 47580 44260 59470
rect 44350 57840 44380 67050
rect 44350 57830 44410 57840
rect 44350 57760 44410 57770
rect 44350 49290 44380 57760
rect 44470 56130 44500 67050
rect 44470 56120 44530 56130
rect 44470 56050 44530 56060
rect 44470 51000 44500 56050
rect 44590 52710 44620 67050
rect 44710 54410 44740 67050
rect 44710 54400 44770 54410
rect 44710 54330 44770 54340
rect 44590 52700 44650 52710
rect 44590 52630 44650 52640
rect 44470 50990 44530 51000
rect 44470 50920 44530 50930
rect 44350 49280 44410 49290
rect 44350 49210 44410 49220
rect 44230 47570 44290 47580
rect 44230 47500 44290 47510
rect 44110 45860 44170 45870
rect 44110 45790 44170 45800
rect 44110 44150 44140 45790
rect 44110 44140 44170 44150
rect 44110 44070 44170 44080
rect 43990 42430 44050 42440
rect 43990 42360 44050 42370
rect 43990 40740 44020 42360
rect 43990 40730 44050 40740
rect 43990 40660 44050 40670
rect 43990 39240 44020 40660
rect 44110 39300 44140 44070
rect 44230 39360 44260 47500
rect 44350 39420 44380 49210
rect 44470 39480 44500 50920
rect 44590 39540 44620 52630
rect 44710 39600 44740 54330
rect 46870 39690 46900 67050
rect 46990 54420 47020 67050
rect 47110 56130 47140 67050
rect 47230 57840 47260 67050
rect 47350 59550 47380 67050
rect 47470 62970 47500 67050
rect 47590 66390 47620 67050
rect 47560 66380 47620 66390
rect 47560 66310 47620 66320
rect 47590 64680 47620 66310
rect 47560 64670 47620 64680
rect 47560 64600 47620 64610
rect 47440 62960 47500 62970
rect 47440 62890 47500 62900
rect 47470 61260 47500 62890
rect 47440 61250 47500 61260
rect 47440 61180 47500 61190
rect 47320 59540 47380 59550
rect 47320 59470 47380 59480
rect 47200 57830 47260 57840
rect 47200 57760 47260 57770
rect 47080 56120 47140 56130
rect 47080 56050 47140 56060
rect 46960 54410 47020 54420
rect 46960 54340 47020 54350
rect 46990 52710 47020 54340
rect 46960 52700 47020 52710
rect 46960 52630 47020 52640
rect 44710 39590 45330 39600
rect 44710 39570 45270 39590
rect 44590 39530 45150 39540
rect 44590 39510 45090 39530
rect 44470 39470 44970 39480
rect 44470 39450 44910 39470
rect 44350 39410 44790 39420
rect 44350 39390 44730 39410
rect 44230 39350 44610 39360
rect 44230 39330 44550 39350
rect 44110 39290 44430 39300
rect 44110 39270 44370 39290
rect 43990 39230 44250 39240
rect 43990 39210 44190 39230
rect 46990 39540 47020 52630
rect 47110 51000 47140 56050
rect 47080 50990 47140 51000
rect 47080 50920 47140 50930
rect 45270 39520 45330 39530
rect 46460 39530 47020 39540
rect 45090 39460 45150 39470
rect 46520 39510 47020 39530
rect 47110 39480 47140 50920
rect 47230 49290 47260 57760
rect 47200 49280 47260 49290
rect 47200 49210 47260 49220
rect 46460 39460 46520 39470
rect 46640 39470 47140 39480
rect 44910 39400 44970 39410
rect 46700 39450 47140 39470
rect 47230 39420 47260 49210
rect 47350 47580 47380 59470
rect 47320 47570 47380 47580
rect 47320 47500 47380 47510
rect 46640 39400 46700 39410
rect 46820 39410 47260 39420
rect 44730 39340 44790 39350
rect 46880 39390 47260 39410
rect 47350 39360 47380 47500
rect 47470 45870 47500 61180
rect 47440 45860 47500 45870
rect 47440 45790 47500 45800
rect 47470 44160 47500 45790
rect 47440 44150 47500 44160
rect 47440 44080 47500 44090
rect 46820 39340 46880 39350
rect 47000 39350 47380 39360
rect 44550 39280 44610 39290
rect 47060 39330 47380 39350
rect 47470 39300 47500 44080
rect 47590 42450 47620 64600
rect 47560 42440 47620 42450
rect 47560 42370 47620 42380
rect 47590 40740 47620 42370
rect 47560 40730 47620 40740
rect 47560 40660 47620 40670
rect 47000 39280 47060 39290
rect 47180 39290 47500 39300
rect 44370 39220 44430 39230
rect 47240 39270 47500 39290
rect 47590 39240 47620 40660
rect 47650 66470 47720 67050
rect 47650 66210 47670 66470
rect 47710 66210 47720 66470
rect 48730 66470 48800 67050
rect 48180 66440 48260 66450
rect 47870 66402 48070 66408
rect 47760 66370 47840 66390
rect 47760 66310 47770 66370
rect 47830 66358 47840 66370
rect 47870 66368 47882 66402
rect 48058 66400 48070 66402
rect 48180 66400 48190 66440
rect 48058 66380 48190 66400
rect 48250 66400 48260 66440
rect 48368 66402 48568 66408
rect 48368 66400 48380 66402
rect 48250 66380 48380 66400
rect 48058 66370 48380 66380
rect 48058 66368 48070 66370
rect 47870 66362 48070 66368
rect 48368 66368 48380 66370
rect 48556 66368 48568 66402
rect 48368 66362 48568 66368
rect 48600 66370 48680 66390
rect 47832 66324 47840 66358
rect 47830 66310 47840 66324
rect 47760 66290 47840 66310
rect 47870 66314 48070 66320
rect 47870 66280 47882 66314
rect 48058 66310 48070 66314
rect 48368 66314 48568 66320
rect 48368 66310 48380 66314
rect 48058 66280 48380 66310
rect 48556 66280 48568 66314
rect 48600 66310 48610 66370
rect 48670 66310 48680 66370
rect 48600 66290 48680 66310
rect 47870 66274 48070 66280
rect 47650 66150 47720 66210
rect 47650 65910 47670 66150
rect 47710 65910 47720 66150
rect 48180 66270 48260 66280
rect 48368 66274 48568 66280
rect 48180 66210 48190 66270
rect 48250 66210 48260 66270
rect 48180 66160 48260 66210
rect 48180 66100 48190 66160
rect 48250 66100 48260 66160
rect 47870 66092 48070 66098
rect 47760 66060 47840 66080
rect 47760 66000 47770 66060
rect 47830 66048 47840 66060
rect 47870 66058 47882 66092
rect 48058 66090 48070 66092
rect 48180 66090 48260 66100
rect 48730 66230 48740 66470
rect 48780 66230 48800 66470
rect 48730 66150 48800 66230
rect 48368 66092 48568 66098
rect 48368 66090 48380 66092
rect 48058 66060 48380 66090
rect 48058 66058 48070 66060
rect 47870 66052 48070 66058
rect 48368 66058 48380 66060
rect 48556 66058 48568 66092
rect 48368 66052 48568 66058
rect 48600 66060 48680 66080
rect 47832 66014 47840 66048
rect 47830 66000 47840 66014
rect 47760 65980 47840 66000
rect 47870 66004 48070 66010
rect 47870 65970 47882 66004
rect 48058 66000 48070 66004
rect 48368 66004 48568 66010
rect 48368 66000 48380 66004
rect 48058 65990 48380 66000
rect 48058 65970 48190 65990
rect 47870 65964 48070 65970
rect 48180 65930 48190 65970
rect 48250 65970 48380 65990
rect 48556 65970 48568 66004
rect 48600 66000 48610 66060
rect 48670 66000 48680 66060
rect 48600 65980 48680 66000
rect 48250 65930 48260 65970
rect 48368 65964 48568 65970
rect 48180 65920 48260 65930
rect 47650 64760 47720 65910
rect 47650 64500 47670 64760
rect 47710 64500 47720 64760
rect 48730 65910 48740 66150
rect 48780 65910 48800 66150
rect 48730 64760 48800 65910
rect 48180 64730 48260 64740
rect 47870 64692 48070 64698
rect 47760 64660 47840 64680
rect 47760 64600 47770 64660
rect 47830 64648 47840 64660
rect 47870 64658 47882 64692
rect 48058 64690 48070 64692
rect 48180 64690 48190 64730
rect 48058 64670 48190 64690
rect 48250 64690 48260 64730
rect 48368 64692 48568 64698
rect 48368 64690 48380 64692
rect 48250 64670 48380 64690
rect 48058 64660 48380 64670
rect 48058 64658 48070 64660
rect 47870 64652 48070 64658
rect 48368 64658 48380 64660
rect 48556 64658 48568 64692
rect 48368 64652 48568 64658
rect 48600 64660 48680 64680
rect 47832 64614 47840 64648
rect 47830 64600 47840 64614
rect 47760 64580 47840 64600
rect 47870 64604 48070 64610
rect 47870 64570 47882 64604
rect 48058 64600 48070 64604
rect 48368 64604 48568 64610
rect 48368 64600 48380 64604
rect 48058 64570 48380 64600
rect 48556 64570 48568 64604
rect 48600 64600 48610 64660
rect 48670 64600 48680 64660
rect 48600 64580 48680 64600
rect 47870 64564 48070 64570
rect 47650 64440 47720 64500
rect 47650 64200 47670 64440
rect 47710 64200 47720 64440
rect 48180 64560 48260 64570
rect 48368 64564 48568 64570
rect 48180 64500 48190 64560
rect 48250 64500 48260 64560
rect 48180 64450 48260 64500
rect 48180 64390 48190 64450
rect 48250 64390 48260 64450
rect 47870 64382 48070 64388
rect 47760 64350 47840 64370
rect 47760 64290 47770 64350
rect 47830 64338 47840 64350
rect 47870 64348 47882 64382
rect 48058 64380 48070 64382
rect 48180 64380 48260 64390
rect 48730 64520 48740 64760
rect 48780 64520 48800 64760
rect 48730 64440 48800 64520
rect 48368 64382 48568 64388
rect 48368 64380 48380 64382
rect 48058 64350 48380 64380
rect 48058 64348 48070 64350
rect 47870 64342 48070 64348
rect 48368 64348 48380 64350
rect 48556 64348 48568 64382
rect 48368 64342 48568 64348
rect 48600 64350 48680 64370
rect 47832 64304 47840 64338
rect 47830 64290 47840 64304
rect 47760 64270 47840 64290
rect 47870 64294 48070 64300
rect 47870 64260 47882 64294
rect 48058 64290 48070 64294
rect 48368 64294 48568 64300
rect 48368 64290 48380 64294
rect 48058 64280 48380 64290
rect 48058 64260 48190 64280
rect 47870 64254 48070 64260
rect 48180 64220 48190 64260
rect 48250 64260 48380 64280
rect 48556 64260 48568 64294
rect 48600 64290 48610 64350
rect 48670 64290 48680 64350
rect 48600 64270 48680 64290
rect 48250 64220 48260 64260
rect 48368 64254 48568 64260
rect 48180 64210 48260 64220
rect 47650 63050 47720 64200
rect 47650 62790 47670 63050
rect 47710 62790 47720 63050
rect 48730 64200 48740 64440
rect 48780 64200 48800 64440
rect 48730 63050 48800 64200
rect 48180 63020 48260 63030
rect 47870 62982 48070 62988
rect 47760 62950 47840 62970
rect 47760 62890 47770 62950
rect 47830 62938 47840 62950
rect 47870 62948 47882 62982
rect 48058 62980 48070 62982
rect 48180 62980 48190 63020
rect 48058 62960 48190 62980
rect 48250 62980 48260 63020
rect 48368 62982 48568 62988
rect 48368 62980 48380 62982
rect 48250 62960 48380 62980
rect 48058 62950 48380 62960
rect 48058 62948 48070 62950
rect 47870 62942 48070 62948
rect 48368 62948 48380 62950
rect 48556 62948 48568 62982
rect 48368 62942 48568 62948
rect 48600 62950 48680 62970
rect 47832 62904 47840 62938
rect 47830 62890 47840 62904
rect 47760 62870 47840 62890
rect 47870 62894 48070 62900
rect 47870 62860 47882 62894
rect 48058 62890 48070 62894
rect 48368 62894 48568 62900
rect 48368 62890 48380 62894
rect 48058 62860 48380 62890
rect 48556 62860 48568 62894
rect 48600 62890 48610 62950
rect 48670 62890 48680 62950
rect 48600 62870 48680 62890
rect 47870 62854 48070 62860
rect 47650 62730 47720 62790
rect 47650 62490 47670 62730
rect 47710 62490 47720 62730
rect 48180 62850 48260 62860
rect 48368 62854 48568 62860
rect 48180 62790 48190 62850
rect 48250 62790 48260 62850
rect 48180 62740 48260 62790
rect 48180 62680 48190 62740
rect 48250 62680 48260 62740
rect 47870 62672 48070 62678
rect 47760 62640 47840 62660
rect 47760 62580 47770 62640
rect 47830 62628 47840 62640
rect 47870 62638 47882 62672
rect 48058 62670 48070 62672
rect 48180 62670 48260 62680
rect 48730 62810 48740 63050
rect 48780 62810 48800 63050
rect 48730 62730 48800 62810
rect 48368 62672 48568 62678
rect 48368 62670 48380 62672
rect 48058 62640 48380 62670
rect 48058 62638 48070 62640
rect 47870 62632 48070 62638
rect 48368 62638 48380 62640
rect 48556 62638 48568 62672
rect 48368 62632 48568 62638
rect 48600 62640 48680 62660
rect 47832 62594 47840 62628
rect 47830 62580 47840 62594
rect 47760 62560 47840 62580
rect 47870 62584 48070 62590
rect 47870 62550 47882 62584
rect 48058 62580 48070 62584
rect 48368 62584 48568 62590
rect 48368 62580 48380 62584
rect 48058 62570 48380 62580
rect 48058 62550 48190 62570
rect 47870 62544 48070 62550
rect 48180 62510 48190 62550
rect 48250 62550 48380 62570
rect 48556 62550 48568 62584
rect 48600 62580 48610 62640
rect 48670 62580 48680 62640
rect 48600 62560 48680 62580
rect 48250 62510 48260 62550
rect 48368 62544 48568 62550
rect 48180 62500 48260 62510
rect 47650 61340 47720 62490
rect 47650 61080 47670 61340
rect 47710 61080 47720 61340
rect 48730 62490 48740 62730
rect 48780 62490 48800 62730
rect 48730 61340 48800 62490
rect 48180 61310 48260 61320
rect 47870 61272 48070 61278
rect 47760 61240 47840 61260
rect 47760 61180 47770 61240
rect 47830 61228 47840 61240
rect 47870 61238 47882 61272
rect 48058 61270 48070 61272
rect 48180 61270 48190 61310
rect 48058 61250 48190 61270
rect 48250 61270 48260 61310
rect 48368 61272 48568 61278
rect 48368 61270 48380 61272
rect 48250 61250 48380 61270
rect 48058 61240 48380 61250
rect 48058 61238 48070 61240
rect 47870 61232 48070 61238
rect 48368 61238 48380 61240
rect 48556 61238 48568 61272
rect 48368 61232 48568 61238
rect 48600 61240 48680 61260
rect 47832 61194 47840 61228
rect 47830 61180 47840 61194
rect 47760 61160 47840 61180
rect 47870 61184 48070 61190
rect 47870 61150 47882 61184
rect 48058 61180 48070 61184
rect 48368 61184 48568 61190
rect 48368 61180 48380 61184
rect 48058 61150 48380 61180
rect 48556 61150 48568 61184
rect 48600 61180 48610 61240
rect 48670 61180 48680 61240
rect 48600 61160 48680 61180
rect 47870 61144 48070 61150
rect 47650 61020 47720 61080
rect 47650 60780 47670 61020
rect 47710 60780 47720 61020
rect 48180 61140 48260 61150
rect 48368 61144 48568 61150
rect 48180 61080 48190 61140
rect 48250 61080 48260 61140
rect 48180 61030 48260 61080
rect 48180 60970 48190 61030
rect 48250 60970 48260 61030
rect 47870 60962 48070 60968
rect 47760 60930 47840 60950
rect 47760 60870 47770 60930
rect 47830 60918 47840 60930
rect 47870 60928 47882 60962
rect 48058 60960 48070 60962
rect 48180 60960 48260 60970
rect 48730 61100 48740 61340
rect 48780 61100 48800 61340
rect 48730 61020 48800 61100
rect 48368 60962 48568 60968
rect 48368 60960 48380 60962
rect 48058 60930 48380 60960
rect 48058 60928 48070 60930
rect 47870 60922 48070 60928
rect 48368 60928 48380 60930
rect 48556 60928 48568 60962
rect 48368 60922 48568 60928
rect 48600 60930 48680 60950
rect 47832 60884 47840 60918
rect 47830 60870 47840 60884
rect 47760 60850 47840 60870
rect 47870 60874 48070 60880
rect 47870 60840 47882 60874
rect 48058 60870 48070 60874
rect 48368 60874 48568 60880
rect 48368 60870 48380 60874
rect 48058 60860 48380 60870
rect 48058 60840 48190 60860
rect 47870 60834 48070 60840
rect 48180 60800 48190 60840
rect 48250 60840 48380 60860
rect 48556 60840 48568 60874
rect 48600 60870 48610 60930
rect 48670 60870 48680 60930
rect 48600 60850 48680 60870
rect 48250 60800 48260 60840
rect 48368 60834 48568 60840
rect 48180 60790 48260 60800
rect 47650 59630 47720 60780
rect 47650 59370 47670 59630
rect 47710 59370 47720 59630
rect 48730 60780 48740 61020
rect 48780 60780 48800 61020
rect 48730 59630 48800 60780
rect 48180 59600 48260 59610
rect 47870 59562 48070 59568
rect 47760 59530 47840 59550
rect 47760 59470 47770 59530
rect 47830 59518 47840 59530
rect 47870 59528 47882 59562
rect 48058 59560 48070 59562
rect 48180 59560 48190 59600
rect 48058 59540 48190 59560
rect 48250 59560 48260 59600
rect 48368 59562 48568 59568
rect 48368 59560 48380 59562
rect 48250 59540 48380 59560
rect 48058 59530 48380 59540
rect 48058 59528 48070 59530
rect 47870 59522 48070 59528
rect 48368 59528 48380 59530
rect 48556 59528 48568 59562
rect 48368 59522 48568 59528
rect 48600 59530 48680 59550
rect 47832 59484 47840 59518
rect 47830 59470 47840 59484
rect 47760 59450 47840 59470
rect 47870 59474 48070 59480
rect 47870 59440 47882 59474
rect 48058 59470 48070 59474
rect 48368 59474 48568 59480
rect 48368 59470 48380 59474
rect 48058 59440 48380 59470
rect 48556 59440 48568 59474
rect 48600 59470 48610 59530
rect 48670 59470 48680 59530
rect 48600 59450 48680 59470
rect 47870 59434 48070 59440
rect 47650 59310 47720 59370
rect 47650 59070 47670 59310
rect 47710 59070 47720 59310
rect 48180 59430 48260 59440
rect 48368 59434 48568 59440
rect 48180 59370 48190 59430
rect 48250 59370 48260 59430
rect 48180 59320 48260 59370
rect 48180 59260 48190 59320
rect 48250 59260 48260 59320
rect 47870 59252 48070 59258
rect 47760 59220 47840 59240
rect 47760 59160 47770 59220
rect 47830 59208 47840 59220
rect 47870 59218 47882 59252
rect 48058 59250 48070 59252
rect 48180 59250 48260 59260
rect 48730 59390 48740 59630
rect 48780 59390 48800 59630
rect 48730 59310 48800 59390
rect 48368 59252 48568 59258
rect 48368 59250 48380 59252
rect 48058 59220 48380 59250
rect 48058 59218 48070 59220
rect 47870 59212 48070 59218
rect 48368 59218 48380 59220
rect 48556 59218 48568 59252
rect 48368 59212 48568 59218
rect 48600 59220 48680 59240
rect 47832 59174 47840 59208
rect 47830 59160 47840 59174
rect 47760 59140 47840 59160
rect 47870 59164 48070 59170
rect 47870 59130 47882 59164
rect 48058 59160 48070 59164
rect 48368 59164 48568 59170
rect 48368 59160 48380 59164
rect 48058 59150 48380 59160
rect 48058 59130 48190 59150
rect 47870 59124 48070 59130
rect 48180 59090 48190 59130
rect 48250 59130 48380 59150
rect 48556 59130 48568 59164
rect 48600 59160 48610 59220
rect 48670 59160 48680 59220
rect 48600 59140 48680 59160
rect 48250 59090 48260 59130
rect 48368 59124 48568 59130
rect 48180 59080 48260 59090
rect 47650 57920 47720 59070
rect 47650 57660 47670 57920
rect 47710 57660 47720 57920
rect 48730 59070 48740 59310
rect 48780 59070 48800 59310
rect 48730 57920 48800 59070
rect 48180 57890 48260 57900
rect 47870 57852 48070 57858
rect 47760 57820 47840 57840
rect 47760 57760 47770 57820
rect 47830 57808 47840 57820
rect 47870 57818 47882 57852
rect 48058 57850 48070 57852
rect 48180 57850 48190 57890
rect 48058 57830 48190 57850
rect 48250 57850 48260 57890
rect 48368 57852 48568 57858
rect 48368 57850 48380 57852
rect 48250 57830 48380 57850
rect 48058 57820 48380 57830
rect 48058 57818 48070 57820
rect 47870 57812 48070 57818
rect 48368 57818 48380 57820
rect 48556 57818 48568 57852
rect 48368 57812 48568 57818
rect 48600 57820 48680 57840
rect 47832 57774 47840 57808
rect 47830 57760 47840 57774
rect 47760 57740 47840 57760
rect 47870 57764 48070 57770
rect 47870 57730 47882 57764
rect 48058 57760 48070 57764
rect 48368 57764 48568 57770
rect 48368 57760 48380 57764
rect 48058 57730 48380 57760
rect 48556 57730 48568 57764
rect 48600 57760 48610 57820
rect 48670 57760 48680 57820
rect 48600 57740 48680 57760
rect 47870 57724 48070 57730
rect 47650 57600 47720 57660
rect 47650 57360 47670 57600
rect 47710 57360 47720 57600
rect 48180 57720 48260 57730
rect 48368 57724 48568 57730
rect 48180 57660 48190 57720
rect 48250 57660 48260 57720
rect 48180 57610 48260 57660
rect 48180 57550 48190 57610
rect 48250 57550 48260 57610
rect 47870 57542 48070 57548
rect 47760 57510 47840 57530
rect 47760 57450 47770 57510
rect 47830 57498 47840 57510
rect 47870 57508 47882 57542
rect 48058 57540 48070 57542
rect 48180 57540 48260 57550
rect 48730 57680 48740 57920
rect 48780 57680 48800 57920
rect 48730 57600 48800 57680
rect 48368 57542 48568 57548
rect 48368 57540 48380 57542
rect 48058 57510 48380 57540
rect 48058 57508 48070 57510
rect 47870 57502 48070 57508
rect 48368 57508 48380 57510
rect 48556 57508 48568 57542
rect 48368 57502 48568 57508
rect 48600 57510 48680 57530
rect 47832 57464 47840 57498
rect 47830 57450 47840 57464
rect 47760 57430 47840 57450
rect 47870 57454 48070 57460
rect 47870 57420 47882 57454
rect 48058 57450 48070 57454
rect 48368 57454 48568 57460
rect 48368 57450 48380 57454
rect 48058 57440 48380 57450
rect 48058 57420 48190 57440
rect 47870 57414 48070 57420
rect 48180 57380 48190 57420
rect 48250 57420 48380 57440
rect 48556 57420 48568 57454
rect 48600 57450 48610 57510
rect 48670 57450 48680 57510
rect 48600 57430 48680 57450
rect 48250 57380 48260 57420
rect 48368 57414 48568 57420
rect 48180 57370 48260 57380
rect 47650 56210 47720 57360
rect 47650 55950 47670 56210
rect 47710 55950 47720 56210
rect 48730 57360 48740 57600
rect 48780 57360 48800 57600
rect 48730 56210 48800 57360
rect 48180 56180 48260 56190
rect 47870 56142 48070 56148
rect 47760 56110 47840 56130
rect 47760 56050 47770 56110
rect 47830 56098 47840 56110
rect 47870 56108 47882 56142
rect 48058 56140 48070 56142
rect 48180 56140 48190 56180
rect 48058 56120 48190 56140
rect 48250 56140 48260 56180
rect 48368 56142 48568 56148
rect 48368 56140 48380 56142
rect 48250 56120 48380 56140
rect 48058 56110 48380 56120
rect 48058 56108 48070 56110
rect 47870 56102 48070 56108
rect 48368 56108 48380 56110
rect 48556 56108 48568 56142
rect 48368 56102 48568 56108
rect 48600 56110 48680 56130
rect 47832 56064 47840 56098
rect 47830 56050 47840 56064
rect 47760 56030 47840 56050
rect 47870 56054 48070 56060
rect 47870 56020 47882 56054
rect 48058 56050 48070 56054
rect 48368 56054 48568 56060
rect 48368 56050 48380 56054
rect 48058 56020 48380 56050
rect 48556 56020 48568 56054
rect 48600 56050 48610 56110
rect 48670 56050 48680 56110
rect 48600 56030 48680 56050
rect 47870 56014 48070 56020
rect 47650 55890 47720 55950
rect 47650 55650 47670 55890
rect 47710 55650 47720 55890
rect 48180 56010 48260 56020
rect 48368 56014 48568 56020
rect 48180 55950 48190 56010
rect 48250 55950 48260 56010
rect 48180 55900 48260 55950
rect 48180 55840 48190 55900
rect 48250 55840 48260 55900
rect 47870 55832 48070 55838
rect 47760 55800 47840 55820
rect 47760 55740 47770 55800
rect 47830 55788 47840 55800
rect 47870 55798 47882 55832
rect 48058 55830 48070 55832
rect 48180 55830 48260 55840
rect 48730 55970 48740 56210
rect 48780 55970 48800 56210
rect 48730 55890 48800 55970
rect 48368 55832 48568 55838
rect 48368 55830 48380 55832
rect 48058 55800 48380 55830
rect 48058 55798 48070 55800
rect 47870 55792 48070 55798
rect 48368 55798 48380 55800
rect 48556 55798 48568 55832
rect 48368 55792 48568 55798
rect 48600 55800 48680 55820
rect 47832 55754 47840 55788
rect 47830 55740 47840 55754
rect 47760 55720 47840 55740
rect 47870 55744 48070 55750
rect 47870 55710 47882 55744
rect 48058 55740 48070 55744
rect 48368 55744 48568 55750
rect 48368 55740 48380 55744
rect 48058 55730 48380 55740
rect 48058 55710 48190 55730
rect 47870 55704 48070 55710
rect 48180 55670 48190 55710
rect 48250 55710 48380 55730
rect 48556 55710 48568 55744
rect 48600 55740 48610 55800
rect 48670 55740 48680 55800
rect 48600 55720 48680 55740
rect 48250 55670 48260 55710
rect 48368 55704 48568 55710
rect 48180 55660 48260 55670
rect 47650 54500 47720 55650
rect 47650 54240 47670 54500
rect 47710 54240 47720 54500
rect 48730 55650 48740 55890
rect 48780 55650 48800 55890
rect 48730 54500 48800 55650
rect 48180 54470 48260 54480
rect 47870 54432 48070 54438
rect 47760 54400 47840 54420
rect 47760 54340 47770 54400
rect 47830 54388 47840 54400
rect 47870 54398 47882 54432
rect 48058 54430 48070 54432
rect 48180 54430 48190 54470
rect 48058 54410 48190 54430
rect 48250 54430 48260 54470
rect 48368 54432 48568 54438
rect 48368 54430 48380 54432
rect 48250 54410 48380 54430
rect 48058 54400 48380 54410
rect 48058 54398 48070 54400
rect 47870 54392 48070 54398
rect 48368 54398 48380 54400
rect 48556 54398 48568 54432
rect 48368 54392 48568 54398
rect 48600 54400 48680 54420
rect 47832 54354 47840 54388
rect 47830 54340 47840 54354
rect 47760 54320 47840 54340
rect 47870 54344 48070 54350
rect 47870 54310 47882 54344
rect 48058 54340 48070 54344
rect 48368 54344 48568 54350
rect 48368 54340 48380 54344
rect 48058 54310 48380 54340
rect 48556 54310 48568 54344
rect 48600 54340 48610 54400
rect 48670 54340 48680 54400
rect 48600 54320 48680 54340
rect 47870 54304 48070 54310
rect 47650 54180 47720 54240
rect 47650 53940 47670 54180
rect 47710 53940 47720 54180
rect 48180 54300 48260 54310
rect 48368 54304 48568 54310
rect 48180 54240 48190 54300
rect 48250 54240 48260 54300
rect 48180 54190 48260 54240
rect 48180 54130 48190 54190
rect 48250 54130 48260 54190
rect 47870 54122 48070 54128
rect 47760 54090 47840 54110
rect 47760 54030 47770 54090
rect 47830 54078 47840 54090
rect 47870 54088 47882 54122
rect 48058 54120 48070 54122
rect 48180 54120 48260 54130
rect 48730 54260 48740 54500
rect 48780 54260 48800 54500
rect 48730 54180 48800 54260
rect 48368 54122 48568 54128
rect 48368 54120 48380 54122
rect 48058 54090 48380 54120
rect 48058 54088 48070 54090
rect 47870 54082 48070 54088
rect 48368 54088 48380 54090
rect 48556 54088 48568 54122
rect 48368 54082 48568 54088
rect 48600 54090 48680 54110
rect 47832 54044 47840 54078
rect 47830 54030 47840 54044
rect 47760 54010 47840 54030
rect 47870 54034 48070 54040
rect 47870 54000 47882 54034
rect 48058 54030 48070 54034
rect 48368 54034 48568 54040
rect 48368 54030 48380 54034
rect 48058 54020 48380 54030
rect 48058 54000 48190 54020
rect 47870 53994 48070 54000
rect 48180 53960 48190 54000
rect 48250 54000 48380 54020
rect 48556 54000 48568 54034
rect 48600 54030 48610 54090
rect 48670 54030 48680 54090
rect 48600 54010 48680 54030
rect 48250 53960 48260 54000
rect 48368 53994 48568 54000
rect 48180 53950 48260 53960
rect 47650 52790 47720 53940
rect 47650 52530 47670 52790
rect 47710 52530 47720 52790
rect 48730 53940 48740 54180
rect 48780 53940 48800 54180
rect 48730 52790 48800 53940
rect 48180 52760 48260 52770
rect 47870 52722 48070 52728
rect 47760 52690 47840 52710
rect 47760 52630 47770 52690
rect 47830 52678 47840 52690
rect 47870 52688 47882 52722
rect 48058 52720 48070 52722
rect 48180 52720 48190 52760
rect 48058 52700 48190 52720
rect 48250 52720 48260 52760
rect 48368 52722 48568 52728
rect 48368 52720 48380 52722
rect 48250 52700 48380 52720
rect 48058 52690 48380 52700
rect 48058 52688 48070 52690
rect 47870 52682 48070 52688
rect 48368 52688 48380 52690
rect 48556 52688 48568 52722
rect 48368 52682 48568 52688
rect 48600 52690 48680 52710
rect 47832 52644 47840 52678
rect 47830 52630 47840 52644
rect 47760 52610 47840 52630
rect 47870 52634 48070 52640
rect 47870 52600 47882 52634
rect 48058 52630 48070 52634
rect 48368 52634 48568 52640
rect 48368 52630 48380 52634
rect 48058 52600 48380 52630
rect 48556 52600 48568 52634
rect 48600 52630 48610 52690
rect 48670 52630 48680 52690
rect 48600 52610 48680 52630
rect 47870 52594 48070 52600
rect 47650 52470 47720 52530
rect 47650 52230 47670 52470
rect 47710 52230 47720 52470
rect 48180 52590 48260 52600
rect 48368 52594 48568 52600
rect 48180 52530 48190 52590
rect 48250 52530 48260 52590
rect 48180 52480 48260 52530
rect 48180 52420 48190 52480
rect 48250 52420 48260 52480
rect 47870 52412 48070 52418
rect 47760 52380 47840 52400
rect 47760 52320 47770 52380
rect 47830 52368 47840 52380
rect 47870 52378 47882 52412
rect 48058 52410 48070 52412
rect 48180 52410 48260 52420
rect 48730 52550 48740 52790
rect 48780 52550 48800 52790
rect 48730 52470 48800 52550
rect 48368 52412 48568 52418
rect 48368 52410 48380 52412
rect 48058 52380 48380 52410
rect 48058 52378 48070 52380
rect 47870 52372 48070 52378
rect 48368 52378 48380 52380
rect 48556 52378 48568 52412
rect 48368 52372 48568 52378
rect 48600 52380 48680 52400
rect 47832 52334 47840 52368
rect 47830 52320 47840 52334
rect 47760 52300 47840 52320
rect 47870 52324 48070 52330
rect 47870 52290 47882 52324
rect 48058 52320 48070 52324
rect 48368 52324 48568 52330
rect 48368 52320 48380 52324
rect 48058 52310 48380 52320
rect 48058 52290 48190 52310
rect 47870 52284 48070 52290
rect 48180 52250 48190 52290
rect 48250 52290 48380 52310
rect 48556 52290 48568 52324
rect 48600 52320 48610 52380
rect 48670 52320 48680 52380
rect 48600 52300 48680 52320
rect 48250 52250 48260 52290
rect 48368 52284 48568 52290
rect 48180 52240 48260 52250
rect 47650 51080 47720 52230
rect 47650 50820 47670 51080
rect 47710 50820 47720 51080
rect 48730 52230 48740 52470
rect 48780 52230 48800 52470
rect 48730 51080 48800 52230
rect 48180 51050 48260 51060
rect 47870 51012 48070 51018
rect 47760 50980 47840 51000
rect 47760 50920 47770 50980
rect 47830 50968 47840 50980
rect 47870 50978 47882 51012
rect 48058 51010 48070 51012
rect 48180 51010 48190 51050
rect 48058 50990 48190 51010
rect 48250 51010 48260 51050
rect 48368 51012 48568 51018
rect 48368 51010 48380 51012
rect 48250 50990 48380 51010
rect 48058 50980 48380 50990
rect 48058 50978 48070 50980
rect 47870 50972 48070 50978
rect 48368 50978 48380 50980
rect 48556 50978 48568 51012
rect 48368 50972 48568 50978
rect 48600 50980 48680 51000
rect 47832 50934 47840 50968
rect 47830 50920 47840 50934
rect 47760 50900 47840 50920
rect 47870 50924 48070 50930
rect 47870 50890 47882 50924
rect 48058 50920 48070 50924
rect 48368 50924 48568 50930
rect 48368 50920 48380 50924
rect 48058 50890 48380 50920
rect 48556 50890 48568 50924
rect 48600 50920 48610 50980
rect 48670 50920 48680 50980
rect 48600 50900 48680 50920
rect 47870 50884 48070 50890
rect 47650 50760 47720 50820
rect 47650 50520 47670 50760
rect 47710 50520 47720 50760
rect 48180 50880 48260 50890
rect 48368 50884 48568 50890
rect 48180 50820 48190 50880
rect 48250 50820 48260 50880
rect 48180 50770 48260 50820
rect 48180 50710 48190 50770
rect 48250 50710 48260 50770
rect 47870 50702 48070 50708
rect 47760 50670 47840 50690
rect 47760 50610 47770 50670
rect 47830 50658 47840 50670
rect 47870 50668 47882 50702
rect 48058 50700 48070 50702
rect 48180 50700 48260 50710
rect 48730 50840 48740 51080
rect 48780 50840 48800 51080
rect 48730 50760 48800 50840
rect 48368 50702 48568 50708
rect 48368 50700 48380 50702
rect 48058 50670 48380 50700
rect 48058 50668 48070 50670
rect 47870 50662 48070 50668
rect 48368 50668 48380 50670
rect 48556 50668 48568 50702
rect 48368 50662 48568 50668
rect 48600 50670 48680 50690
rect 47832 50624 47840 50658
rect 47830 50610 47840 50624
rect 47760 50590 47840 50610
rect 47870 50614 48070 50620
rect 47870 50580 47882 50614
rect 48058 50610 48070 50614
rect 48368 50614 48568 50620
rect 48368 50610 48380 50614
rect 48058 50600 48380 50610
rect 48058 50580 48190 50600
rect 47870 50574 48070 50580
rect 48180 50540 48190 50580
rect 48250 50580 48380 50600
rect 48556 50580 48568 50614
rect 48600 50610 48610 50670
rect 48670 50610 48680 50670
rect 48600 50590 48680 50610
rect 48250 50540 48260 50580
rect 48368 50574 48568 50580
rect 48180 50530 48260 50540
rect 47650 49370 47720 50520
rect 47650 49110 47670 49370
rect 47710 49110 47720 49370
rect 48730 50520 48740 50760
rect 48780 50520 48800 50760
rect 48730 49370 48800 50520
rect 48180 49340 48260 49350
rect 47870 49302 48070 49308
rect 47760 49270 47840 49290
rect 47760 49210 47770 49270
rect 47830 49258 47840 49270
rect 47870 49268 47882 49302
rect 48058 49300 48070 49302
rect 48180 49300 48190 49340
rect 48058 49280 48190 49300
rect 48250 49300 48260 49340
rect 48368 49302 48568 49308
rect 48368 49300 48380 49302
rect 48250 49280 48380 49300
rect 48058 49270 48380 49280
rect 48058 49268 48070 49270
rect 47870 49262 48070 49268
rect 48368 49268 48380 49270
rect 48556 49268 48568 49302
rect 48368 49262 48568 49268
rect 48600 49270 48680 49290
rect 47832 49224 47840 49258
rect 47830 49210 47840 49224
rect 47760 49190 47840 49210
rect 47870 49214 48070 49220
rect 47870 49180 47882 49214
rect 48058 49210 48070 49214
rect 48368 49214 48568 49220
rect 48368 49210 48380 49214
rect 48058 49180 48380 49210
rect 48556 49180 48568 49214
rect 48600 49210 48610 49270
rect 48670 49210 48680 49270
rect 48600 49190 48680 49210
rect 47870 49174 48070 49180
rect 47650 49050 47720 49110
rect 47650 48810 47670 49050
rect 47710 48810 47720 49050
rect 48180 49170 48260 49180
rect 48368 49174 48568 49180
rect 48180 49110 48190 49170
rect 48250 49110 48260 49170
rect 48180 49060 48260 49110
rect 48180 49000 48190 49060
rect 48250 49000 48260 49060
rect 47870 48992 48070 48998
rect 47760 48960 47840 48980
rect 47760 48900 47770 48960
rect 47830 48948 47840 48960
rect 47870 48958 47882 48992
rect 48058 48990 48070 48992
rect 48180 48990 48260 49000
rect 48730 49130 48740 49370
rect 48780 49130 48800 49370
rect 48730 49050 48800 49130
rect 48368 48992 48568 48998
rect 48368 48990 48380 48992
rect 48058 48960 48380 48990
rect 48058 48958 48070 48960
rect 47870 48952 48070 48958
rect 48368 48958 48380 48960
rect 48556 48958 48568 48992
rect 48368 48952 48568 48958
rect 48600 48960 48680 48980
rect 47832 48914 47840 48948
rect 47830 48900 47840 48914
rect 47760 48880 47840 48900
rect 47870 48904 48070 48910
rect 47870 48870 47882 48904
rect 48058 48900 48070 48904
rect 48368 48904 48568 48910
rect 48368 48900 48380 48904
rect 48058 48890 48380 48900
rect 48058 48870 48190 48890
rect 47870 48864 48070 48870
rect 48180 48830 48190 48870
rect 48250 48870 48380 48890
rect 48556 48870 48568 48904
rect 48600 48900 48610 48960
rect 48670 48900 48680 48960
rect 48600 48880 48680 48900
rect 48250 48830 48260 48870
rect 48368 48864 48568 48870
rect 48180 48820 48260 48830
rect 47650 47660 47720 48810
rect 47650 47400 47670 47660
rect 47710 47400 47720 47660
rect 48730 48810 48740 49050
rect 48780 48810 48800 49050
rect 48730 47660 48800 48810
rect 48180 47630 48260 47640
rect 47870 47592 48070 47598
rect 47760 47560 47840 47580
rect 47760 47500 47770 47560
rect 47830 47548 47840 47560
rect 47870 47558 47882 47592
rect 48058 47590 48070 47592
rect 48180 47590 48190 47630
rect 48058 47570 48190 47590
rect 48250 47590 48260 47630
rect 48368 47592 48568 47598
rect 48368 47590 48380 47592
rect 48250 47570 48380 47590
rect 48058 47560 48380 47570
rect 48058 47558 48070 47560
rect 47870 47552 48070 47558
rect 48368 47558 48380 47560
rect 48556 47558 48568 47592
rect 48368 47552 48568 47558
rect 48600 47560 48680 47580
rect 47832 47514 47840 47548
rect 47830 47500 47840 47514
rect 47760 47480 47840 47500
rect 47870 47504 48070 47510
rect 47870 47470 47882 47504
rect 48058 47500 48070 47504
rect 48368 47504 48568 47510
rect 48368 47500 48380 47504
rect 48058 47470 48380 47500
rect 48556 47470 48568 47504
rect 48600 47500 48610 47560
rect 48670 47500 48680 47560
rect 48600 47480 48680 47500
rect 47870 47464 48070 47470
rect 47650 47340 47720 47400
rect 47650 47100 47670 47340
rect 47710 47100 47720 47340
rect 48180 47460 48260 47470
rect 48368 47464 48568 47470
rect 48180 47400 48190 47460
rect 48250 47400 48260 47460
rect 48180 47350 48260 47400
rect 48180 47290 48190 47350
rect 48250 47290 48260 47350
rect 47870 47282 48070 47288
rect 47760 47250 47840 47270
rect 47760 47190 47770 47250
rect 47830 47238 47840 47250
rect 47870 47248 47882 47282
rect 48058 47280 48070 47282
rect 48180 47280 48260 47290
rect 48730 47420 48740 47660
rect 48780 47420 48800 47660
rect 48730 47340 48800 47420
rect 48368 47282 48568 47288
rect 48368 47280 48380 47282
rect 48058 47250 48380 47280
rect 48058 47248 48070 47250
rect 47870 47242 48070 47248
rect 48368 47248 48380 47250
rect 48556 47248 48568 47282
rect 48368 47242 48568 47248
rect 48600 47250 48680 47270
rect 47832 47204 47840 47238
rect 47830 47190 47840 47204
rect 47760 47170 47840 47190
rect 47870 47194 48070 47200
rect 47870 47160 47882 47194
rect 48058 47190 48070 47194
rect 48368 47194 48568 47200
rect 48368 47190 48380 47194
rect 48058 47180 48380 47190
rect 48058 47160 48190 47180
rect 47870 47154 48070 47160
rect 48180 47120 48190 47160
rect 48250 47160 48380 47180
rect 48556 47160 48568 47194
rect 48600 47190 48610 47250
rect 48670 47190 48680 47250
rect 48600 47170 48680 47190
rect 48250 47120 48260 47160
rect 48368 47154 48568 47160
rect 48180 47110 48260 47120
rect 47650 45950 47720 47100
rect 47650 45690 47670 45950
rect 47710 45690 47720 45950
rect 48730 47100 48740 47340
rect 48780 47100 48800 47340
rect 48730 45950 48800 47100
rect 48180 45920 48260 45930
rect 47870 45882 48070 45888
rect 47760 45850 47840 45870
rect 47760 45790 47770 45850
rect 47830 45838 47840 45850
rect 47870 45848 47882 45882
rect 48058 45880 48070 45882
rect 48180 45880 48190 45920
rect 48058 45860 48190 45880
rect 48250 45880 48260 45920
rect 48368 45882 48568 45888
rect 48368 45880 48380 45882
rect 48250 45860 48380 45880
rect 48058 45850 48380 45860
rect 48058 45848 48070 45850
rect 47870 45842 48070 45848
rect 48368 45848 48380 45850
rect 48556 45848 48568 45882
rect 48368 45842 48568 45848
rect 48600 45850 48680 45870
rect 47832 45804 47840 45838
rect 47830 45790 47840 45804
rect 47760 45770 47840 45790
rect 47870 45794 48070 45800
rect 47870 45760 47882 45794
rect 48058 45790 48070 45794
rect 48368 45794 48568 45800
rect 48368 45790 48380 45794
rect 48058 45760 48380 45790
rect 48556 45760 48568 45794
rect 48600 45790 48610 45850
rect 48670 45790 48680 45850
rect 48600 45770 48680 45790
rect 47870 45754 48070 45760
rect 47650 45630 47720 45690
rect 47650 45390 47670 45630
rect 47710 45390 47720 45630
rect 48180 45750 48260 45760
rect 48368 45754 48568 45760
rect 48180 45690 48190 45750
rect 48250 45690 48260 45750
rect 48180 45640 48260 45690
rect 48180 45580 48190 45640
rect 48250 45580 48260 45640
rect 47870 45572 48070 45578
rect 47760 45540 47840 45560
rect 47760 45480 47770 45540
rect 47830 45528 47840 45540
rect 47870 45538 47882 45572
rect 48058 45570 48070 45572
rect 48180 45570 48260 45580
rect 48730 45710 48740 45950
rect 48780 45710 48800 45950
rect 48730 45630 48800 45710
rect 48368 45572 48568 45578
rect 48368 45570 48380 45572
rect 48058 45540 48380 45570
rect 48058 45538 48070 45540
rect 47870 45532 48070 45538
rect 48368 45538 48380 45540
rect 48556 45538 48568 45572
rect 48368 45532 48568 45538
rect 48600 45540 48680 45560
rect 47832 45494 47840 45528
rect 47830 45480 47840 45494
rect 47760 45460 47840 45480
rect 47870 45484 48070 45490
rect 47870 45450 47882 45484
rect 48058 45480 48070 45484
rect 48368 45484 48568 45490
rect 48368 45480 48380 45484
rect 48058 45470 48380 45480
rect 48058 45450 48190 45470
rect 47870 45444 48070 45450
rect 48180 45410 48190 45450
rect 48250 45450 48380 45470
rect 48556 45450 48568 45484
rect 48600 45480 48610 45540
rect 48670 45480 48680 45540
rect 48600 45460 48680 45480
rect 48250 45410 48260 45450
rect 48368 45444 48568 45450
rect 48180 45400 48260 45410
rect 47650 44240 47720 45390
rect 47650 43980 47670 44240
rect 47710 43980 47720 44240
rect 48730 45390 48740 45630
rect 48780 45390 48800 45630
rect 48730 44240 48800 45390
rect 48180 44210 48260 44220
rect 47870 44172 48070 44178
rect 47760 44140 47840 44160
rect 47760 44080 47770 44140
rect 47830 44128 47840 44140
rect 47870 44138 47882 44172
rect 48058 44170 48070 44172
rect 48180 44170 48190 44210
rect 48058 44150 48190 44170
rect 48250 44170 48260 44210
rect 48368 44172 48568 44178
rect 48368 44170 48380 44172
rect 48250 44150 48380 44170
rect 48058 44140 48380 44150
rect 48058 44138 48070 44140
rect 47870 44132 48070 44138
rect 48368 44138 48380 44140
rect 48556 44138 48568 44172
rect 48368 44132 48568 44138
rect 48600 44140 48680 44160
rect 47832 44094 47840 44128
rect 47830 44080 47840 44094
rect 47760 44060 47840 44080
rect 47870 44084 48070 44090
rect 47870 44050 47882 44084
rect 48058 44080 48070 44084
rect 48368 44084 48568 44090
rect 48368 44080 48380 44084
rect 48058 44050 48380 44080
rect 48556 44050 48568 44084
rect 48600 44080 48610 44140
rect 48670 44080 48680 44140
rect 48600 44060 48680 44080
rect 47870 44044 48070 44050
rect 47650 43920 47720 43980
rect 47650 43680 47670 43920
rect 47710 43680 47720 43920
rect 48180 44040 48260 44050
rect 48368 44044 48568 44050
rect 48180 43980 48190 44040
rect 48250 43980 48260 44040
rect 48180 43930 48260 43980
rect 48180 43870 48190 43930
rect 48250 43870 48260 43930
rect 47870 43862 48070 43868
rect 47760 43830 47840 43850
rect 47760 43770 47770 43830
rect 47830 43818 47840 43830
rect 47870 43828 47882 43862
rect 48058 43860 48070 43862
rect 48180 43860 48260 43870
rect 48730 44000 48740 44240
rect 48780 44000 48800 44240
rect 48730 43920 48800 44000
rect 48368 43862 48568 43868
rect 48368 43860 48380 43862
rect 48058 43830 48380 43860
rect 48058 43828 48070 43830
rect 47870 43822 48070 43828
rect 48368 43828 48380 43830
rect 48556 43828 48568 43862
rect 48368 43822 48568 43828
rect 48600 43830 48680 43850
rect 47832 43784 47840 43818
rect 47830 43770 47840 43784
rect 47760 43750 47840 43770
rect 47870 43774 48070 43780
rect 47870 43740 47882 43774
rect 48058 43770 48070 43774
rect 48368 43774 48568 43780
rect 48368 43770 48380 43774
rect 48058 43760 48380 43770
rect 48058 43740 48190 43760
rect 47870 43734 48070 43740
rect 48180 43700 48190 43740
rect 48250 43740 48380 43760
rect 48556 43740 48568 43774
rect 48600 43770 48610 43830
rect 48670 43770 48680 43830
rect 48600 43750 48680 43770
rect 48250 43700 48260 43740
rect 48368 43734 48568 43740
rect 48180 43690 48260 43700
rect 47650 42530 47720 43680
rect 47650 42270 47670 42530
rect 47710 42270 47720 42530
rect 48730 43680 48740 43920
rect 48780 43680 48800 43920
rect 48730 42530 48800 43680
rect 48180 42500 48260 42510
rect 47870 42462 48070 42468
rect 47760 42430 47840 42450
rect 47760 42370 47770 42430
rect 47830 42418 47840 42430
rect 47870 42428 47882 42462
rect 48058 42460 48070 42462
rect 48180 42460 48190 42500
rect 48058 42440 48190 42460
rect 48250 42460 48260 42500
rect 48368 42462 48568 42468
rect 48368 42460 48380 42462
rect 48250 42440 48380 42460
rect 48058 42430 48380 42440
rect 48058 42428 48070 42430
rect 47870 42422 48070 42428
rect 48368 42428 48380 42430
rect 48556 42428 48568 42462
rect 48368 42422 48568 42428
rect 48600 42430 48680 42450
rect 47832 42384 47840 42418
rect 47830 42370 47840 42384
rect 47760 42350 47840 42370
rect 47870 42374 48070 42380
rect 47870 42340 47882 42374
rect 48058 42370 48070 42374
rect 48368 42374 48568 42380
rect 48368 42370 48380 42374
rect 48058 42340 48380 42370
rect 48556 42340 48568 42374
rect 48600 42370 48610 42430
rect 48670 42370 48680 42430
rect 48600 42350 48680 42370
rect 47870 42334 48070 42340
rect 47650 42210 47720 42270
rect 47650 41970 47670 42210
rect 47710 41970 47720 42210
rect 48180 42330 48260 42340
rect 48368 42334 48568 42340
rect 48180 42270 48190 42330
rect 48250 42270 48260 42330
rect 48180 42220 48260 42270
rect 48180 42160 48190 42220
rect 48250 42160 48260 42220
rect 47870 42152 48070 42158
rect 47760 42120 47840 42140
rect 47760 42060 47770 42120
rect 47830 42108 47840 42120
rect 47870 42118 47882 42152
rect 48058 42150 48070 42152
rect 48180 42150 48260 42160
rect 48730 42290 48740 42530
rect 48780 42290 48800 42530
rect 48730 42210 48800 42290
rect 48368 42152 48568 42158
rect 48368 42150 48380 42152
rect 48058 42120 48380 42150
rect 48058 42118 48070 42120
rect 47870 42112 48070 42118
rect 48368 42118 48380 42120
rect 48556 42118 48568 42152
rect 48368 42112 48568 42118
rect 48600 42120 48680 42140
rect 47832 42074 47840 42108
rect 47830 42060 47840 42074
rect 47760 42040 47840 42060
rect 47870 42064 48070 42070
rect 47870 42030 47882 42064
rect 48058 42060 48070 42064
rect 48368 42064 48568 42070
rect 48368 42060 48380 42064
rect 48058 42050 48380 42060
rect 48058 42030 48190 42050
rect 47870 42024 48070 42030
rect 48180 41990 48190 42030
rect 48250 42030 48380 42050
rect 48556 42030 48568 42064
rect 48600 42060 48610 42120
rect 48670 42060 48680 42120
rect 48600 42040 48680 42060
rect 48250 41990 48260 42030
rect 48368 42024 48568 42030
rect 48180 41980 48260 41990
rect 47650 40820 47720 41970
rect 47650 40560 47670 40820
rect 47710 40560 47720 40820
rect 48730 41970 48740 42210
rect 48780 41970 48800 42210
rect 48730 40820 48800 41970
rect 48180 40790 48260 40800
rect 47870 40752 48070 40758
rect 47760 40720 47840 40740
rect 47760 40660 47770 40720
rect 47830 40708 47840 40720
rect 47870 40718 47882 40752
rect 48058 40750 48070 40752
rect 48180 40750 48190 40790
rect 48058 40730 48190 40750
rect 48250 40750 48260 40790
rect 48368 40752 48568 40758
rect 48368 40750 48380 40752
rect 48250 40730 48380 40750
rect 48058 40720 48380 40730
rect 48058 40718 48070 40720
rect 47870 40712 48070 40718
rect 48368 40718 48380 40720
rect 48556 40718 48568 40752
rect 48368 40712 48568 40718
rect 48600 40720 48680 40740
rect 47832 40674 47840 40708
rect 47830 40660 47840 40674
rect 47760 40640 47840 40660
rect 47870 40664 48070 40670
rect 47870 40630 47882 40664
rect 48058 40660 48070 40664
rect 48368 40664 48568 40670
rect 48368 40660 48380 40664
rect 48058 40630 48380 40660
rect 48556 40630 48568 40664
rect 48600 40660 48610 40720
rect 48670 40660 48680 40720
rect 48600 40640 48680 40660
rect 47870 40624 48070 40630
rect 47650 40500 47720 40560
rect 47650 40260 47670 40500
rect 47710 40260 47720 40500
rect 48180 40620 48260 40630
rect 48368 40624 48568 40630
rect 48180 40560 48190 40620
rect 48250 40560 48260 40620
rect 48180 40510 48260 40560
rect 48180 40450 48190 40510
rect 48250 40450 48260 40510
rect 47870 40442 48070 40448
rect 47760 40410 47840 40430
rect 47760 40350 47770 40410
rect 47830 40398 47840 40410
rect 47870 40408 47882 40442
rect 48058 40440 48070 40442
rect 48180 40440 48260 40450
rect 48730 40580 48740 40820
rect 48780 40580 48800 40820
rect 48730 40500 48800 40580
rect 48368 40442 48568 40448
rect 48368 40440 48380 40442
rect 48058 40410 48380 40440
rect 48058 40408 48070 40410
rect 47870 40402 48070 40408
rect 48368 40408 48380 40410
rect 48556 40408 48568 40442
rect 48368 40402 48568 40408
rect 48600 40410 48680 40430
rect 47832 40364 47840 40398
rect 47830 40350 47840 40364
rect 47760 40330 47840 40350
rect 47870 40354 48070 40360
rect 47870 40320 47882 40354
rect 48058 40350 48070 40354
rect 48368 40354 48568 40360
rect 48368 40350 48380 40354
rect 48058 40340 48380 40350
rect 48058 40320 48190 40340
rect 47870 40314 48070 40320
rect 48180 40280 48190 40320
rect 48250 40320 48380 40340
rect 48556 40320 48568 40354
rect 48600 40350 48610 40410
rect 48670 40350 48680 40410
rect 48600 40330 48680 40350
rect 48250 40280 48260 40320
rect 48368 40314 48568 40320
rect 48180 40270 48260 40280
rect 47650 39690 47720 40260
rect 48730 40260 48740 40500
rect 48780 40260 48800 40500
rect 48730 39690 48800 40260
rect 47650 39680 47730 39690
rect 47650 39620 47660 39680
rect 47720 39620 47730 39680
rect 48720 39680 48800 39690
rect 48720 39620 48730 39680
rect 48790 39620 48800 39680
rect 48720 39610 48800 39620
rect 48830 66480 48860 67050
rect 48830 66470 48890 66480
rect 48830 66400 48890 66410
rect 48830 64770 48860 66400
rect 48920 65950 48950 67050
rect 48890 65940 48950 65950
rect 48890 65870 48950 65880
rect 48830 64760 48890 64770
rect 48830 64690 48890 64700
rect 48830 63060 48860 64690
rect 48920 64240 48950 65870
rect 48890 64230 48950 64240
rect 48890 64160 48950 64170
rect 48830 63050 48890 63060
rect 48830 62980 48890 62990
rect 48830 61350 48860 62980
rect 48920 62530 48950 64160
rect 48890 62520 48950 62530
rect 48890 62450 48950 62460
rect 48830 61340 48890 61350
rect 48830 61270 48890 61280
rect 48830 59640 48860 61270
rect 48920 60820 48950 62450
rect 48890 60810 48950 60820
rect 48890 60740 48950 60750
rect 48830 59630 48890 59640
rect 48830 59560 48890 59570
rect 48830 57930 48860 59560
rect 48920 59110 48950 60740
rect 48890 59100 48950 59110
rect 48890 59030 48950 59040
rect 48830 57920 48890 57930
rect 48830 57850 48890 57860
rect 48830 56220 48860 57850
rect 48920 57400 48950 59030
rect 48890 57390 48950 57400
rect 48890 57320 48950 57330
rect 48830 56210 48890 56220
rect 48830 56140 48890 56150
rect 48830 54510 48860 56140
rect 48920 55690 48950 57320
rect 48890 55680 48950 55690
rect 48890 55610 48950 55620
rect 48830 54500 48890 54510
rect 48830 54430 48890 54440
rect 48830 52800 48860 54430
rect 48920 53980 48950 55610
rect 48890 53970 48950 53980
rect 48890 53900 48950 53910
rect 48830 52790 48890 52800
rect 48830 52720 48890 52730
rect 48830 51090 48860 52720
rect 48920 52270 48950 53900
rect 48890 52260 48950 52270
rect 48890 52190 48950 52200
rect 48830 51080 48890 51090
rect 48830 51010 48890 51020
rect 48830 49380 48860 51010
rect 48920 50560 48950 52190
rect 48890 50550 48950 50560
rect 48890 50480 48950 50490
rect 48830 49370 48890 49380
rect 48830 49300 48890 49310
rect 48830 47670 48860 49300
rect 48920 48850 48950 50480
rect 48890 48840 48950 48850
rect 48890 48770 48950 48780
rect 48830 47660 48890 47670
rect 48830 47590 48890 47600
rect 48830 45960 48860 47590
rect 48920 47140 48950 48770
rect 48890 47130 48950 47140
rect 48890 47060 48950 47070
rect 48830 45950 48890 45960
rect 48830 45880 48890 45890
rect 48830 44250 48860 45880
rect 48920 45430 48950 47060
rect 48890 45420 48950 45430
rect 48890 45350 48950 45360
rect 48830 44240 48890 44250
rect 48830 44170 48890 44180
rect 48830 42540 48860 44170
rect 48920 43720 48950 45350
rect 48890 43710 48950 43720
rect 48890 43640 48950 43650
rect 48830 42530 48890 42540
rect 48830 42460 48890 42470
rect 48830 40830 48860 42460
rect 48920 42010 48950 43640
rect 48890 42000 48950 42010
rect 48890 41930 48950 41940
rect 48830 40820 48890 40830
rect 48830 40750 48890 40760
rect 47180 39220 47240 39230
rect 47360 39230 47620 39240
rect 44190 39160 44250 39170
rect 47420 39210 47620 39230
rect 47360 39160 47420 39170
rect 48830 38840 48860 40750
rect 48920 40300 48950 41930
rect 48890 40290 48950 40300
rect 48890 40220 48950 40230
rect 48920 39690 48950 40220
rect 48890 39680 48950 39690
rect 48890 39610 48950 39620
rect 48980 66390 49010 67050
rect 48980 66380 49040 66390
rect 48980 66310 49040 66320
rect 48980 64680 49010 66310
rect 48980 64670 49040 64680
rect 48980 64600 49040 64610
rect 48980 42450 49010 64600
rect 49100 62970 49130 67050
rect 49100 62960 49160 62970
rect 49100 62890 49160 62900
rect 49100 61260 49130 62890
rect 49100 61250 49160 61260
rect 49100 61180 49160 61190
rect 49100 45870 49130 61180
rect 49220 59550 49250 67050
rect 49220 59540 49280 59550
rect 49220 59470 49280 59480
rect 49220 47580 49250 59470
rect 49340 57840 49370 67050
rect 49340 57830 49400 57840
rect 49340 57760 49400 57770
rect 49340 49290 49370 57760
rect 49460 56130 49490 67050
rect 49460 56120 49520 56130
rect 49460 56050 49520 56060
rect 49460 51000 49490 56050
rect 49580 54420 49610 67050
rect 49580 54410 49640 54420
rect 49580 54340 49640 54350
rect 49580 52710 49610 54340
rect 49580 52700 49640 52710
rect 49580 52630 49640 52640
rect 49460 50990 49520 51000
rect 49460 50920 49520 50930
rect 49340 49280 49400 49290
rect 49340 49210 49400 49220
rect 49220 47570 49280 47580
rect 49220 47500 49280 47510
rect 49100 45860 49160 45870
rect 49100 45790 49160 45800
rect 49100 44160 49130 45790
rect 49100 44150 49160 44160
rect 49100 44080 49160 44090
rect 48980 42440 49040 42450
rect 48980 42370 49040 42380
rect 48980 40740 49010 42370
rect 48980 40730 49040 40740
rect 48980 40660 49040 40670
rect 48980 39240 49010 40660
rect 49100 39300 49130 44080
rect 49220 39360 49250 47500
rect 49340 39420 49370 49210
rect 49460 39480 49490 50920
rect 49580 39540 49610 52630
rect 49700 39690 49730 67050
rect 51860 39690 51890 67050
rect 51980 39690 52010 67050
rect 52100 39690 52130 67050
rect 52220 57840 52250 67050
rect 52340 59550 52370 67050
rect 52460 62970 52490 67050
rect 52580 66390 52610 67050
rect 52550 66380 52610 66390
rect 52550 66310 52610 66320
rect 52580 64680 52610 66310
rect 52550 64670 52610 64680
rect 52550 64600 52610 64610
rect 52430 62960 52490 62970
rect 52430 62890 52490 62900
rect 52460 61250 52490 62890
rect 52430 61240 52490 61250
rect 52430 61170 52490 61180
rect 52310 59540 52370 59550
rect 52310 59470 52370 59480
rect 52190 57830 52250 57840
rect 52190 57760 52250 57770
rect 52220 56130 52250 57760
rect 52190 56120 52250 56130
rect 52190 56050 52250 56060
rect 52220 54420 52250 56050
rect 52190 54410 52250 54420
rect 52190 54340 52250 54350
rect 52220 52710 52250 54340
rect 52190 52700 52250 52710
rect 52190 52630 52250 52640
rect 52220 51000 52250 52630
rect 52190 50990 52250 51000
rect 52190 50920 52250 50930
rect 52220 49290 52250 50920
rect 52190 49280 52250 49290
rect 52190 49210 52250 49220
rect 49580 39530 50140 39540
rect 49580 39510 50080 39530
rect 49460 39470 49960 39480
rect 49460 39450 49900 39470
rect 49340 39410 49780 39420
rect 49340 39390 49720 39410
rect 49220 39350 49600 39360
rect 49220 39330 49540 39350
rect 49100 39290 49420 39300
rect 49100 39270 49360 39290
rect 48980 39230 49240 39240
rect 48980 39210 49180 39230
rect 50080 39460 50140 39470
rect 52220 39420 52250 49210
rect 52340 47580 52370 59470
rect 52310 47570 52370 47580
rect 52310 47500 52370 47510
rect 49900 39400 49960 39410
rect 51810 39410 52250 39420
rect 49720 39340 49780 39350
rect 51870 39390 52250 39410
rect 52340 39360 52370 47500
rect 52460 45870 52490 61170
rect 52430 45860 52490 45870
rect 52430 45790 52490 45800
rect 52460 44160 52490 45790
rect 52430 44150 52490 44160
rect 52430 44080 52490 44090
rect 51810 39340 51870 39350
rect 51990 39350 52370 39360
rect 49540 39280 49600 39290
rect 52050 39330 52370 39350
rect 52460 39300 52490 44080
rect 52580 42450 52610 64600
rect 52550 42440 52610 42450
rect 52550 42370 52610 42380
rect 52580 40740 52610 42370
rect 52550 40730 52610 40740
rect 52550 40660 52610 40670
rect 51990 39280 52050 39290
rect 52170 39290 52490 39300
rect 49360 39220 49420 39230
rect 52230 39270 52490 39290
rect 52580 39240 52610 40660
rect 52640 66470 52710 67050
rect 52640 66210 52660 66470
rect 52700 66210 52710 66470
rect 53720 66470 53790 67050
rect 53170 66440 53250 66450
rect 52860 66402 53060 66408
rect 52750 66370 52830 66390
rect 52750 66310 52760 66370
rect 52820 66358 52830 66370
rect 52860 66368 52872 66402
rect 53048 66400 53060 66402
rect 53170 66400 53180 66440
rect 53048 66380 53180 66400
rect 53240 66400 53250 66440
rect 53358 66402 53558 66408
rect 53358 66400 53370 66402
rect 53240 66380 53370 66400
rect 53048 66370 53370 66380
rect 53048 66368 53060 66370
rect 52860 66362 53060 66368
rect 53358 66368 53370 66370
rect 53546 66368 53558 66402
rect 53358 66362 53558 66368
rect 53590 66370 53670 66390
rect 52822 66324 52830 66358
rect 52820 66310 52830 66324
rect 52750 66290 52830 66310
rect 52860 66314 53060 66320
rect 52860 66280 52872 66314
rect 53048 66310 53060 66314
rect 53358 66314 53558 66320
rect 53358 66310 53370 66314
rect 53048 66280 53370 66310
rect 53546 66280 53558 66314
rect 53590 66310 53600 66370
rect 53660 66310 53670 66370
rect 53590 66290 53670 66310
rect 52860 66274 53060 66280
rect 52640 66150 52710 66210
rect 52640 65910 52660 66150
rect 52700 65910 52710 66150
rect 53170 66270 53250 66280
rect 53358 66274 53558 66280
rect 53170 66210 53180 66270
rect 53240 66210 53250 66270
rect 53170 66160 53250 66210
rect 53170 66100 53180 66160
rect 53240 66100 53250 66160
rect 52860 66092 53060 66098
rect 52750 66060 52830 66080
rect 52750 66000 52760 66060
rect 52820 66048 52830 66060
rect 52860 66058 52872 66092
rect 53048 66090 53060 66092
rect 53170 66090 53250 66100
rect 53720 66230 53730 66470
rect 53770 66230 53790 66470
rect 53720 66150 53790 66230
rect 53358 66092 53558 66098
rect 53358 66090 53370 66092
rect 53048 66060 53370 66090
rect 53048 66058 53060 66060
rect 52860 66052 53060 66058
rect 53358 66058 53370 66060
rect 53546 66058 53558 66092
rect 53358 66052 53558 66058
rect 53590 66060 53670 66080
rect 52822 66014 52830 66048
rect 52820 66000 52830 66014
rect 52750 65980 52830 66000
rect 52860 66004 53060 66010
rect 52860 65970 52872 66004
rect 53048 66000 53060 66004
rect 53358 66004 53558 66010
rect 53358 66000 53370 66004
rect 53048 65990 53370 66000
rect 53048 65970 53180 65990
rect 52860 65964 53060 65970
rect 53170 65930 53180 65970
rect 53240 65970 53370 65990
rect 53546 65970 53558 66004
rect 53590 66000 53600 66060
rect 53660 66000 53670 66060
rect 53590 65980 53670 66000
rect 53240 65930 53250 65970
rect 53358 65964 53558 65970
rect 53170 65920 53250 65930
rect 52640 64760 52710 65910
rect 52640 64500 52660 64760
rect 52700 64500 52710 64760
rect 53720 65910 53730 66150
rect 53770 65910 53790 66150
rect 53720 64760 53790 65910
rect 53170 64730 53250 64740
rect 52860 64692 53060 64698
rect 52750 64660 52830 64680
rect 52750 64600 52760 64660
rect 52820 64648 52830 64660
rect 52860 64658 52872 64692
rect 53048 64690 53060 64692
rect 53170 64690 53180 64730
rect 53048 64670 53180 64690
rect 53240 64690 53250 64730
rect 53358 64692 53558 64698
rect 53358 64690 53370 64692
rect 53240 64670 53370 64690
rect 53048 64660 53370 64670
rect 53048 64658 53060 64660
rect 52860 64652 53060 64658
rect 53358 64658 53370 64660
rect 53546 64658 53558 64692
rect 53358 64652 53558 64658
rect 53590 64660 53670 64680
rect 52822 64614 52830 64648
rect 52820 64600 52830 64614
rect 52750 64580 52830 64600
rect 52860 64604 53060 64610
rect 52860 64570 52872 64604
rect 53048 64600 53060 64604
rect 53358 64604 53558 64610
rect 53358 64600 53370 64604
rect 53048 64570 53370 64600
rect 53546 64570 53558 64604
rect 53590 64600 53600 64660
rect 53660 64600 53670 64660
rect 53590 64580 53670 64600
rect 52860 64564 53060 64570
rect 52640 64440 52710 64500
rect 52640 64200 52660 64440
rect 52700 64200 52710 64440
rect 53170 64560 53250 64570
rect 53358 64564 53558 64570
rect 53170 64500 53180 64560
rect 53240 64500 53250 64560
rect 53170 64450 53250 64500
rect 53170 64390 53180 64450
rect 53240 64390 53250 64450
rect 52860 64382 53060 64388
rect 52750 64350 52830 64370
rect 52750 64290 52760 64350
rect 52820 64338 52830 64350
rect 52860 64348 52872 64382
rect 53048 64380 53060 64382
rect 53170 64380 53250 64390
rect 53720 64520 53730 64760
rect 53770 64520 53790 64760
rect 53720 64440 53790 64520
rect 53358 64382 53558 64388
rect 53358 64380 53370 64382
rect 53048 64350 53370 64380
rect 53048 64348 53060 64350
rect 52860 64342 53060 64348
rect 53358 64348 53370 64350
rect 53546 64348 53558 64382
rect 53358 64342 53558 64348
rect 53590 64350 53670 64370
rect 52822 64304 52830 64338
rect 52820 64290 52830 64304
rect 52750 64270 52830 64290
rect 52860 64294 53060 64300
rect 52860 64260 52872 64294
rect 53048 64290 53060 64294
rect 53358 64294 53558 64300
rect 53358 64290 53370 64294
rect 53048 64280 53370 64290
rect 53048 64260 53180 64280
rect 52860 64254 53060 64260
rect 53170 64220 53180 64260
rect 53240 64260 53370 64280
rect 53546 64260 53558 64294
rect 53590 64290 53600 64350
rect 53660 64290 53670 64350
rect 53590 64270 53670 64290
rect 53240 64220 53250 64260
rect 53358 64254 53558 64260
rect 53170 64210 53250 64220
rect 52640 63050 52710 64200
rect 52640 62790 52660 63050
rect 52700 62790 52710 63050
rect 53720 64200 53730 64440
rect 53770 64200 53790 64440
rect 53720 63050 53790 64200
rect 53170 63020 53250 63030
rect 52860 62982 53060 62988
rect 52750 62950 52830 62970
rect 52750 62890 52760 62950
rect 52820 62938 52830 62950
rect 52860 62948 52872 62982
rect 53048 62980 53060 62982
rect 53170 62980 53180 63020
rect 53048 62960 53180 62980
rect 53240 62980 53250 63020
rect 53358 62982 53558 62988
rect 53358 62980 53370 62982
rect 53240 62960 53370 62980
rect 53048 62950 53370 62960
rect 53048 62948 53060 62950
rect 52860 62942 53060 62948
rect 53358 62948 53370 62950
rect 53546 62948 53558 62982
rect 53358 62942 53558 62948
rect 53590 62950 53670 62970
rect 52822 62904 52830 62938
rect 52820 62890 52830 62904
rect 52750 62870 52830 62890
rect 52860 62894 53060 62900
rect 52860 62860 52872 62894
rect 53048 62890 53060 62894
rect 53358 62894 53558 62900
rect 53358 62890 53370 62894
rect 53048 62860 53370 62890
rect 53546 62860 53558 62894
rect 53590 62890 53600 62950
rect 53660 62890 53670 62950
rect 53590 62870 53670 62890
rect 52860 62854 53060 62860
rect 52640 62730 52710 62790
rect 52640 62490 52660 62730
rect 52700 62490 52710 62730
rect 53170 62850 53250 62860
rect 53358 62854 53558 62860
rect 53170 62790 53180 62850
rect 53240 62790 53250 62850
rect 53170 62740 53250 62790
rect 53170 62680 53180 62740
rect 53240 62680 53250 62740
rect 52860 62672 53060 62678
rect 52750 62640 52830 62660
rect 52750 62580 52760 62640
rect 52820 62628 52830 62640
rect 52860 62638 52872 62672
rect 53048 62670 53060 62672
rect 53170 62670 53250 62680
rect 53720 62810 53730 63050
rect 53770 62810 53790 63050
rect 53720 62730 53790 62810
rect 53358 62672 53558 62678
rect 53358 62670 53370 62672
rect 53048 62640 53370 62670
rect 53048 62638 53060 62640
rect 52860 62632 53060 62638
rect 53358 62638 53370 62640
rect 53546 62638 53558 62672
rect 53358 62632 53558 62638
rect 53590 62640 53670 62660
rect 52822 62594 52830 62628
rect 52820 62580 52830 62594
rect 52750 62560 52830 62580
rect 52860 62584 53060 62590
rect 52860 62550 52872 62584
rect 53048 62580 53060 62584
rect 53358 62584 53558 62590
rect 53358 62580 53370 62584
rect 53048 62570 53370 62580
rect 53048 62550 53180 62570
rect 52860 62544 53060 62550
rect 53170 62510 53180 62550
rect 53240 62550 53370 62570
rect 53546 62550 53558 62584
rect 53590 62580 53600 62640
rect 53660 62580 53670 62640
rect 53590 62560 53670 62580
rect 53240 62510 53250 62550
rect 53358 62544 53558 62550
rect 53170 62500 53250 62510
rect 52640 61340 52710 62490
rect 52640 61080 52660 61340
rect 52700 61080 52710 61340
rect 53720 62490 53730 62730
rect 53770 62490 53790 62730
rect 53720 61340 53790 62490
rect 53170 61310 53250 61320
rect 52860 61272 53060 61278
rect 52750 61240 52830 61260
rect 52750 61180 52760 61240
rect 52820 61228 52830 61240
rect 52860 61238 52872 61272
rect 53048 61270 53060 61272
rect 53170 61270 53180 61310
rect 53048 61250 53180 61270
rect 53240 61270 53250 61310
rect 53358 61272 53558 61278
rect 53358 61270 53370 61272
rect 53240 61250 53370 61270
rect 53048 61240 53370 61250
rect 53048 61238 53060 61240
rect 52860 61232 53060 61238
rect 53358 61238 53370 61240
rect 53546 61238 53558 61272
rect 53358 61232 53558 61238
rect 53590 61240 53670 61260
rect 52822 61194 52830 61228
rect 52820 61180 52830 61194
rect 52750 61160 52830 61180
rect 52860 61184 53060 61190
rect 52860 61150 52872 61184
rect 53048 61180 53060 61184
rect 53358 61184 53558 61190
rect 53358 61180 53370 61184
rect 53048 61150 53370 61180
rect 53546 61150 53558 61184
rect 53590 61180 53600 61240
rect 53660 61180 53670 61240
rect 53590 61160 53670 61180
rect 52860 61144 53060 61150
rect 52640 61020 52710 61080
rect 52640 60780 52660 61020
rect 52700 60780 52710 61020
rect 53170 61140 53250 61150
rect 53358 61144 53558 61150
rect 53170 61080 53180 61140
rect 53240 61080 53250 61140
rect 53170 61030 53250 61080
rect 53170 60970 53180 61030
rect 53240 60970 53250 61030
rect 52860 60962 53060 60968
rect 52750 60930 52830 60950
rect 52750 60870 52760 60930
rect 52820 60918 52830 60930
rect 52860 60928 52872 60962
rect 53048 60960 53060 60962
rect 53170 60960 53250 60970
rect 53720 61100 53730 61340
rect 53770 61100 53790 61340
rect 53720 61020 53790 61100
rect 53358 60962 53558 60968
rect 53358 60960 53370 60962
rect 53048 60930 53370 60960
rect 53048 60928 53060 60930
rect 52860 60922 53060 60928
rect 53358 60928 53370 60930
rect 53546 60928 53558 60962
rect 53358 60922 53558 60928
rect 53590 60930 53670 60950
rect 52822 60884 52830 60918
rect 52820 60870 52830 60884
rect 52750 60850 52830 60870
rect 52860 60874 53060 60880
rect 52860 60840 52872 60874
rect 53048 60870 53060 60874
rect 53358 60874 53558 60880
rect 53358 60870 53370 60874
rect 53048 60860 53370 60870
rect 53048 60840 53180 60860
rect 52860 60834 53060 60840
rect 53170 60800 53180 60840
rect 53240 60840 53370 60860
rect 53546 60840 53558 60874
rect 53590 60870 53600 60930
rect 53660 60870 53670 60930
rect 53590 60850 53670 60870
rect 53240 60800 53250 60840
rect 53358 60834 53558 60840
rect 53170 60790 53250 60800
rect 52640 59630 52710 60780
rect 52640 59370 52660 59630
rect 52700 59370 52710 59630
rect 53720 60780 53730 61020
rect 53770 60780 53790 61020
rect 53720 59630 53790 60780
rect 53170 59600 53250 59610
rect 52860 59562 53060 59568
rect 52750 59530 52830 59550
rect 52750 59470 52760 59530
rect 52820 59518 52830 59530
rect 52860 59528 52872 59562
rect 53048 59560 53060 59562
rect 53170 59560 53180 59600
rect 53048 59540 53180 59560
rect 53240 59560 53250 59600
rect 53358 59562 53558 59568
rect 53358 59560 53370 59562
rect 53240 59540 53370 59560
rect 53048 59530 53370 59540
rect 53048 59528 53060 59530
rect 52860 59522 53060 59528
rect 53358 59528 53370 59530
rect 53546 59528 53558 59562
rect 53358 59522 53558 59528
rect 53590 59530 53670 59550
rect 52822 59484 52830 59518
rect 52820 59470 52830 59484
rect 52750 59450 52830 59470
rect 52860 59474 53060 59480
rect 52860 59440 52872 59474
rect 53048 59470 53060 59474
rect 53358 59474 53558 59480
rect 53358 59470 53370 59474
rect 53048 59440 53370 59470
rect 53546 59440 53558 59474
rect 53590 59470 53600 59530
rect 53660 59470 53670 59530
rect 53590 59450 53670 59470
rect 52860 59434 53060 59440
rect 52640 59310 52710 59370
rect 52640 59070 52660 59310
rect 52700 59070 52710 59310
rect 53170 59430 53250 59440
rect 53358 59434 53558 59440
rect 53170 59370 53180 59430
rect 53240 59370 53250 59430
rect 53170 59320 53250 59370
rect 53170 59260 53180 59320
rect 53240 59260 53250 59320
rect 52860 59252 53060 59258
rect 52750 59220 52830 59240
rect 52750 59160 52760 59220
rect 52820 59208 52830 59220
rect 52860 59218 52872 59252
rect 53048 59250 53060 59252
rect 53170 59250 53250 59260
rect 53720 59390 53730 59630
rect 53770 59390 53790 59630
rect 53720 59310 53790 59390
rect 53358 59252 53558 59258
rect 53358 59250 53370 59252
rect 53048 59220 53370 59250
rect 53048 59218 53060 59220
rect 52860 59212 53060 59218
rect 53358 59218 53370 59220
rect 53546 59218 53558 59252
rect 53358 59212 53558 59218
rect 53590 59220 53670 59240
rect 52822 59174 52830 59208
rect 52820 59160 52830 59174
rect 52750 59140 52830 59160
rect 52860 59164 53060 59170
rect 52860 59130 52872 59164
rect 53048 59160 53060 59164
rect 53358 59164 53558 59170
rect 53358 59160 53370 59164
rect 53048 59150 53370 59160
rect 53048 59130 53180 59150
rect 52860 59124 53060 59130
rect 53170 59090 53180 59130
rect 53240 59130 53370 59150
rect 53546 59130 53558 59164
rect 53590 59160 53600 59220
rect 53660 59160 53670 59220
rect 53590 59140 53670 59160
rect 53240 59090 53250 59130
rect 53358 59124 53558 59130
rect 53170 59080 53250 59090
rect 52640 57920 52710 59070
rect 52640 57660 52660 57920
rect 52700 57660 52710 57920
rect 53720 59070 53730 59310
rect 53770 59070 53790 59310
rect 53720 57920 53790 59070
rect 53170 57890 53250 57900
rect 52860 57852 53060 57858
rect 52750 57820 52830 57840
rect 52750 57760 52760 57820
rect 52820 57808 52830 57820
rect 52860 57818 52872 57852
rect 53048 57850 53060 57852
rect 53170 57850 53180 57890
rect 53048 57830 53180 57850
rect 53240 57850 53250 57890
rect 53358 57852 53558 57858
rect 53358 57850 53370 57852
rect 53240 57830 53370 57850
rect 53048 57820 53370 57830
rect 53048 57818 53060 57820
rect 52860 57812 53060 57818
rect 53358 57818 53370 57820
rect 53546 57818 53558 57852
rect 53358 57812 53558 57818
rect 53590 57820 53670 57840
rect 52822 57774 52830 57808
rect 52820 57760 52830 57774
rect 52750 57740 52830 57760
rect 52860 57764 53060 57770
rect 52860 57730 52872 57764
rect 53048 57760 53060 57764
rect 53358 57764 53558 57770
rect 53358 57760 53370 57764
rect 53048 57730 53370 57760
rect 53546 57730 53558 57764
rect 53590 57760 53600 57820
rect 53660 57760 53670 57820
rect 53590 57740 53670 57760
rect 52860 57724 53060 57730
rect 52640 57600 52710 57660
rect 52640 57360 52660 57600
rect 52700 57360 52710 57600
rect 53170 57720 53250 57730
rect 53358 57724 53558 57730
rect 53170 57660 53180 57720
rect 53240 57660 53250 57720
rect 53170 57610 53250 57660
rect 53170 57550 53180 57610
rect 53240 57550 53250 57610
rect 52860 57542 53060 57548
rect 52750 57510 52830 57530
rect 52750 57450 52760 57510
rect 52820 57498 52830 57510
rect 52860 57508 52872 57542
rect 53048 57540 53060 57542
rect 53170 57540 53250 57550
rect 53720 57680 53730 57920
rect 53770 57680 53790 57920
rect 53720 57600 53790 57680
rect 53358 57542 53558 57548
rect 53358 57540 53370 57542
rect 53048 57510 53370 57540
rect 53048 57508 53060 57510
rect 52860 57502 53060 57508
rect 53358 57508 53370 57510
rect 53546 57508 53558 57542
rect 53358 57502 53558 57508
rect 53590 57510 53670 57530
rect 52822 57464 52830 57498
rect 52820 57450 52830 57464
rect 52750 57430 52830 57450
rect 52860 57454 53060 57460
rect 52860 57420 52872 57454
rect 53048 57450 53060 57454
rect 53358 57454 53558 57460
rect 53358 57450 53370 57454
rect 53048 57440 53370 57450
rect 53048 57420 53180 57440
rect 52860 57414 53060 57420
rect 53170 57380 53180 57420
rect 53240 57420 53370 57440
rect 53546 57420 53558 57454
rect 53590 57450 53600 57510
rect 53660 57450 53670 57510
rect 53590 57430 53670 57450
rect 53240 57380 53250 57420
rect 53358 57414 53558 57420
rect 53170 57370 53250 57380
rect 52640 56210 52710 57360
rect 52640 55950 52660 56210
rect 52700 55950 52710 56210
rect 53720 57360 53730 57600
rect 53770 57360 53790 57600
rect 53720 56210 53790 57360
rect 53170 56180 53250 56190
rect 52860 56142 53060 56148
rect 52750 56110 52830 56130
rect 52750 56050 52760 56110
rect 52820 56098 52830 56110
rect 52860 56108 52872 56142
rect 53048 56140 53060 56142
rect 53170 56140 53180 56180
rect 53048 56120 53180 56140
rect 53240 56140 53250 56180
rect 53358 56142 53558 56148
rect 53358 56140 53370 56142
rect 53240 56120 53370 56140
rect 53048 56110 53370 56120
rect 53048 56108 53060 56110
rect 52860 56102 53060 56108
rect 53358 56108 53370 56110
rect 53546 56108 53558 56142
rect 53358 56102 53558 56108
rect 53590 56110 53670 56130
rect 52822 56064 52830 56098
rect 52820 56050 52830 56064
rect 52750 56030 52830 56050
rect 52860 56054 53060 56060
rect 52860 56020 52872 56054
rect 53048 56050 53060 56054
rect 53358 56054 53558 56060
rect 53358 56050 53370 56054
rect 53048 56020 53370 56050
rect 53546 56020 53558 56054
rect 53590 56050 53600 56110
rect 53660 56050 53670 56110
rect 53590 56030 53670 56050
rect 52860 56014 53060 56020
rect 52640 55890 52710 55950
rect 52640 55650 52660 55890
rect 52700 55650 52710 55890
rect 53170 56010 53250 56020
rect 53358 56014 53558 56020
rect 53170 55950 53180 56010
rect 53240 55950 53250 56010
rect 53170 55900 53250 55950
rect 53170 55840 53180 55900
rect 53240 55840 53250 55900
rect 52860 55832 53060 55838
rect 52750 55800 52830 55820
rect 52750 55740 52760 55800
rect 52820 55788 52830 55800
rect 52860 55798 52872 55832
rect 53048 55830 53060 55832
rect 53170 55830 53250 55840
rect 53720 55970 53730 56210
rect 53770 55970 53790 56210
rect 53720 55890 53790 55970
rect 53358 55832 53558 55838
rect 53358 55830 53370 55832
rect 53048 55800 53370 55830
rect 53048 55798 53060 55800
rect 52860 55792 53060 55798
rect 53358 55798 53370 55800
rect 53546 55798 53558 55832
rect 53358 55792 53558 55798
rect 53590 55800 53670 55820
rect 52822 55754 52830 55788
rect 52820 55740 52830 55754
rect 52750 55720 52830 55740
rect 52860 55744 53060 55750
rect 52860 55710 52872 55744
rect 53048 55740 53060 55744
rect 53358 55744 53558 55750
rect 53358 55740 53370 55744
rect 53048 55730 53370 55740
rect 53048 55710 53180 55730
rect 52860 55704 53060 55710
rect 53170 55670 53180 55710
rect 53240 55710 53370 55730
rect 53546 55710 53558 55744
rect 53590 55740 53600 55800
rect 53660 55740 53670 55800
rect 53590 55720 53670 55740
rect 53240 55670 53250 55710
rect 53358 55704 53558 55710
rect 53170 55660 53250 55670
rect 52640 54500 52710 55650
rect 52640 54240 52660 54500
rect 52700 54240 52710 54500
rect 53720 55650 53730 55890
rect 53770 55650 53790 55890
rect 53720 54500 53790 55650
rect 53170 54470 53250 54480
rect 52860 54432 53060 54438
rect 52750 54400 52830 54420
rect 52750 54340 52760 54400
rect 52820 54388 52830 54400
rect 52860 54398 52872 54432
rect 53048 54430 53060 54432
rect 53170 54430 53180 54470
rect 53048 54410 53180 54430
rect 53240 54430 53250 54470
rect 53358 54432 53558 54438
rect 53358 54430 53370 54432
rect 53240 54410 53370 54430
rect 53048 54400 53370 54410
rect 53048 54398 53060 54400
rect 52860 54392 53060 54398
rect 53358 54398 53370 54400
rect 53546 54398 53558 54432
rect 53358 54392 53558 54398
rect 53590 54400 53670 54420
rect 52822 54354 52830 54388
rect 52820 54340 52830 54354
rect 52750 54320 52830 54340
rect 52860 54344 53060 54350
rect 52860 54310 52872 54344
rect 53048 54340 53060 54344
rect 53358 54344 53558 54350
rect 53358 54340 53370 54344
rect 53048 54310 53370 54340
rect 53546 54310 53558 54344
rect 53590 54340 53600 54400
rect 53660 54340 53670 54400
rect 53590 54320 53670 54340
rect 52860 54304 53060 54310
rect 52640 54180 52710 54240
rect 52640 53940 52660 54180
rect 52700 53940 52710 54180
rect 53170 54300 53250 54310
rect 53358 54304 53558 54310
rect 53170 54240 53180 54300
rect 53240 54240 53250 54300
rect 53170 54190 53250 54240
rect 53170 54130 53180 54190
rect 53240 54130 53250 54190
rect 52860 54122 53060 54128
rect 52750 54090 52830 54110
rect 52750 54030 52760 54090
rect 52820 54078 52830 54090
rect 52860 54088 52872 54122
rect 53048 54120 53060 54122
rect 53170 54120 53250 54130
rect 53720 54260 53730 54500
rect 53770 54260 53790 54500
rect 53720 54180 53790 54260
rect 53358 54122 53558 54128
rect 53358 54120 53370 54122
rect 53048 54090 53370 54120
rect 53048 54088 53060 54090
rect 52860 54082 53060 54088
rect 53358 54088 53370 54090
rect 53546 54088 53558 54122
rect 53358 54082 53558 54088
rect 53590 54090 53670 54110
rect 52822 54044 52830 54078
rect 52820 54030 52830 54044
rect 52750 54010 52830 54030
rect 52860 54034 53060 54040
rect 52860 54000 52872 54034
rect 53048 54030 53060 54034
rect 53358 54034 53558 54040
rect 53358 54030 53370 54034
rect 53048 54020 53370 54030
rect 53048 54000 53180 54020
rect 52860 53994 53060 54000
rect 53170 53960 53180 54000
rect 53240 54000 53370 54020
rect 53546 54000 53558 54034
rect 53590 54030 53600 54090
rect 53660 54030 53670 54090
rect 53590 54010 53670 54030
rect 53240 53960 53250 54000
rect 53358 53994 53558 54000
rect 53170 53950 53250 53960
rect 52640 52790 52710 53940
rect 52640 52530 52660 52790
rect 52700 52530 52710 52790
rect 53720 53940 53730 54180
rect 53770 53940 53790 54180
rect 53720 52790 53790 53940
rect 53170 52760 53250 52770
rect 52860 52722 53060 52728
rect 52750 52690 52830 52710
rect 52750 52630 52760 52690
rect 52820 52678 52830 52690
rect 52860 52688 52872 52722
rect 53048 52720 53060 52722
rect 53170 52720 53180 52760
rect 53048 52700 53180 52720
rect 53240 52720 53250 52760
rect 53358 52722 53558 52728
rect 53358 52720 53370 52722
rect 53240 52700 53370 52720
rect 53048 52690 53370 52700
rect 53048 52688 53060 52690
rect 52860 52682 53060 52688
rect 53358 52688 53370 52690
rect 53546 52688 53558 52722
rect 53358 52682 53558 52688
rect 53590 52690 53670 52710
rect 52822 52644 52830 52678
rect 52820 52630 52830 52644
rect 52750 52610 52830 52630
rect 52860 52634 53060 52640
rect 52860 52600 52872 52634
rect 53048 52630 53060 52634
rect 53358 52634 53558 52640
rect 53358 52630 53370 52634
rect 53048 52600 53370 52630
rect 53546 52600 53558 52634
rect 53590 52630 53600 52690
rect 53660 52630 53670 52690
rect 53590 52610 53670 52630
rect 52860 52594 53060 52600
rect 52640 52470 52710 52530
rect 52640 52230 52660 52470
rect 52700 52230 52710 52470
rect 53170 52590 53250 52600
rect 53358 52594 53558 52600
rect 53170 52530 53180 52590
rect 53240 52530 53250 52590
rect 53170 52480 53250 52530
rect 53170 52420 53180 52480
rect 53240 52420 53250 52480
rect 52860 52412 53060 52418
rect 52750 52380 52830 52400
rect 52750 52320 52760 52380
rect 52820 52368 52830 52380
rect 52860 52378 52872 52412
rect 53048 52410 53060 52412
rect 53170 52410 53250 52420
rect 53720 52550 53730 52790
rect 53770 52550 53790 52790
rect 53720 52470 53790 52550
rect 53358 52412 53558 52418
rect 53358 52410 53370 52412
rect 53048 52380 53370 52410
rect 53048 52378 53060 52380
rect 52860 52372 53060 52378
rect 53358 52378 53370 52380
rect 53546 52378 53558 52412
rect 53358 52372 53558 52378
rect 53590 52380 53670 52400
rect 52822 52334 52830 52368
rect 52820 52320 52830 52334
rect 52750 52300 52830 52320
rect 52860 52324 53060 52330
rect 52860 52290 52872 52324
rect 53048 52320 53060 52324
rect 53358 52324 53558 52330
rect 53358 52320 53370 52324
rect 53048 52310 53370 52320
rect 53048 52290 53180 52310
rect 52860 52284 53060 52290
rect 53170 52250 53180 52290
rect 53240 52290 53370 52310
rect 53546 52290 53558 52324
rect 53590 52320 53600 52380
rect 53660 52320 53670 52380
rect 53590 52300 53670 52320
rect 53240 52250 53250 52290
rect 53358 52284 53558 52290
rect 53170 52240 53250 52250
rect 52640 51080 52710 52230
rect 52640 50820 52660 51080
rect 52700 50820 52710 51080
rect 53720 52230 53730 52470
rect 53770 52230 53790 52470
rect 53720 51080 53790 52230
rect 53170 51050 53250 51060
rect 52860 51012 53060 51018
rect 52750 50980 52830 51000
rect 52750 50920 52760 50980
rect 52820 50968 52830 50980
rect 52860 50978 52872 51012
rect 53048 51010 53060 51012
rect 53170 51010 53180 51050
rect 53048 50990 53180 51010
rect 53240 51010 53250 51050
rect 53358 51012 53558 51018
rect 53358 51010 53370 51012
rect 53240 50990 53370 51010
rect 53048 50980 53370 50990
rect 53048 50978 53060 50980
rect 52860 50972 53060 50978
rect 53358 50978 53370 50980
rect 53546 50978 53558 51012
rect 53358 50972 53558 50978
rect 53590 50980 53670 51000
rect 52822 50934 52830 50968
rect 52820 50920 52830 50934
rect 52750 50900 52830 50920
rect 52860 50924 53060 50930
rect 52860 50890 52872 50924
rect 53048 50920 53060 50924
rect 53358 50924 53558 50930
rect 53358 50920 53370 50924
rect 53048 50890 53370 50920
rect 53546 50890 53558 50924
rect 53590 50920 53600 50980
rect 53660 50920 53670 50980
rect 53590 50900 53670 50920
rect 52860 50884 53060 50890
rect 52640 50760 52710 50820
rect 52640 50520 52660 50760
rect 52700 50520 52710 50760
rect 53170 50880 53250 50890
rect 53358 50884 53558 50890
rect 53170 50820 53180 50880
rect 53240 50820 53250 50880
rect 53170 50770 53250 50820
rect 53170 50710 53180 50770
rect 53240 50710 53250 50770
rect 52860 50702 53060 50708
rect 52750 50670 52830 50690
rect 52750 50610 52760 50670
rect 52820 50658 52830 50670
rect 52860 50668 52872 50702
rect 53048 50700 53060 50702
rect 53170 50700 53250 50710
rect 53720 50840 53730 51080
rect 53770 50840 53790 51080
rect 53720 50760 53790 50840
rect 53358 50702 53558 50708
rect 53358 50700 53370 50702
rect 53048 50670 53370 50700
rect 53048 50668 53060 50670
rect 52860 50662 53060 50668
rect 53358 50668 53370 50670
rect 53546 50668 53558 50702
rect 53358 50662 53558 50668
rect 53590 50670 53670 50690
rect 52822 50624 52830 50658
rect 52820 50610 52830 50624
rect 52750 50590 52830 50610
rect 52860 50614 53060 50620
rect 52860 50580 52872 50614
rect 53048 50610 53060 50614
rect 53358 50614 53558 50620
rect 53358 50610 53370 50614
rect 53048 50600 53370 50610
rect 53048 50580 53180 50600
rect 52860 50574 53060 50580
rect 53170 50540 53180 50580
rect 53240 50580 53370 50600
rect 53546 50580 53558 50614
rect 53590 50610 53600 50670
rect 53660 50610 53670 50670
rect 53590 50590 53670 50610
rect 53240 50540 53250 50580
rect 53358 50574 53558 50580
rect 53170 50530 53250 50540
rect 52640 49370 52710 50520
rect 52640 49110 52660 49370
rect 52700 49110 52710 49370
rect 53720 50520 53730 50760
rect 53770 50520 53790 50760
rect 53720 49370 53790 50520
rect 53170 49340 53250 49350
rect 52860 49302 53060 49308
rect 52750 49270 52830 49290
rect 52750 49210 52760 49270
rect 52820 49258 52830 49270
rect 52860 49268 52872 49302
rect 53048 49300 53060 49302
rect 53170 49300 53180 49340
rect 53048 49280 53180 49300
rect 53240 49300 53250 49340
rect 53358 49302 53558 49308
rect 53358 49300 53370 49302
rect 53240 49280 53370 49300
rect 53048 49270 53370 49280
rect 53048 49268 53060 49270
rect 52860 49262 53060 49268
rect 53358 49268 53370 49270
rect 53546 49268 53558 49302
rect 53358 49262 53558 49268
rect 53590 49270 53670 49290
rect 52822 49224 52830 49258
rect 52820 49210 52830 49224
rect 52750 49190 52830 49210
rect 52860 49214 53060 49220
rect 52860 49180 52872 49214
rect 53048 49210 53060 49214
rect 53358 49214 53558 49220
rect 53358 49210 53370 49214
rect 53048 49180 53370 49210
rect 53546 49180 53558 49214
rect 53590 49210 53600 49270
rect 53660 49210 53670 49270
rect 53590 49190 53670 49210
rect 52860 49174 53060 49180
rect 52640 49050 52710 49110
rect 52640 48810 52660 49050
rect 52700 48810 52710 49050
rect 53170 49170 53250 49180
rect 53358 49174 53558 49180
rect 53170 49110 53180 49170
rect 53240 49110 53250 49170
rect 53170 49060 53250 49110
rect 53170 49000 53180 49060
rect 53240 49000 53250 49060
rect 52860 48992 53060 48998
rect 52750 48960 52830 48980
rect 52750 48900 52760 48960
rect 52820 48948 52830 48960
rect 52860 48958 52872 48992
rect 53048 48990 53060 48992
rect 53170 48990 53250 49000
rect 53720 49130 53730 49370
rect 53770 49130 53790 49370
rect 53720 49050 53790 49130
rect 53358 48992 53558 48998
rect 53358 48990 53370 48992
rect 53048 48960 53370 48990
rect 53048 48958 53060 48960
rect 52860 48952 53060 48958
rect 53358 48958 53370 48960
rect 53546 48958 53558 48992
rect 53358 48952 53558 48958
rect 53590 48960 53670 48980
rect 52822 48914 52830 48948
rect 52820 48900 52830 48914
rect 52750 48880 52830 48900
rect 52860 48904 53060 48910
rect 52860 48870 52872 48904
rect 53048 48900 53060 48904
rect 53358 48904 53558 48910
rect 53358 48900 53370 48904
rect 53048 48890 53370 48900
rect 53048 48870 53180 48890
rect 52860 48864 53060 48870
rect 53170 48830 53180 48870
rect 53240 48870 53370 48890
rect 53546 48870 53558 48904
rect 53590 48900 53600 48960
rect 53660 48900 53670 48960
rect 53590 48880 53670 48900
rect 53240 48830 53250 48870
rect 53358 48864 53558 48870
rect 53170 48820 53250 48830
rect 52640 47660 52710 48810
rect 52640 47400 52660 47660
rect 52700 47400 52710 47660
rect 53720 48810 53730 49050
rect 53770 48810 53790 49050
rect 53720 47660 53790 48810
rect 53170 47630 53250 47640
rect 52860 47592 53060 47598
rect 52750 47560 52830 47580
rect 52750 47500 52760 47560
rect 52820 47548 52830 47560
rect 52860 47558 52872 47592
rect 53048 47590 53060 47592
rect 53170 47590 53180 47630
rect 53048 47570 53180 47590
rect 53240 47590 53250 47630
rect 53358 47592 53558 47598
rect 53358 47590 53370 47592
rect 53240 47570 53370 47590
rect 53048 47560 53370 47570
rect 53048 47558 53060 47560
rect 52860 47552 53060 47558
rect 53358 47558 53370 47560
rect 53546 47558 53558 47592
rect 53358 47552 53558 47558
rect 53590 47560 53670 47580
rect 52822 47514 52830 47548
rect 52820 47500 52830 47514
rect 52750 47480 52830 47500
rect 52860 47504 53060 47510
rect 52860 47470 52872 47504
rect 53048 47500 53060 47504
rect 53358 47504 53558 47510
rect 53358 47500 53370 47504
rect 53048 47470 53370 47500
rect 53546 47470 53558 47504
rect 53590 47500 53600 47560
rect 53660 47500 53670 47560
rect 53590 47480 53670 47500
rect 52860 47464 53060 47470
rect 52640 47340 52710 47400
rect 52640 47100 52660 47340
rect 52700 47100 52710 47340
rect 53170 47460 53250 47470
rect 53358 47464 53558 47470
rect 53170 47400 53180 47460
rect 53240 47400 53250 47460
rect 53170 47350 53250 47400
rect 53170 47290 53180 47350
rect 53240 47290 53250 47350
rect 52860 47282 53060 47288
rect 52750 47250 52830 47270
rect 52750 47190 52760 47250
rect 52820 47238 52830 47250
rect 52860 47248 52872 47282
rect 53048 47280 53060 47282
rect 53170 47280 53250 47290
rect 53720 47420 53730 47660
rect 53770 47420 53790 47660
rect 53720 47340 53790 47420
rect 53358 47282 53558 47288
rect 53358 47280 53370 47282
rect 53048 47250 53370 47280
rect 53048 47248 53060 47250
rect 52860 47242 53060 47248
rect 53358 47248 53370 47250
rect 53546 47248 53558 47282
rect 53358 47242 53558 47248
rect 53590 47250 53670 47270
rect 52822 47204 52830 47238
rect 52820 47190 52830 47204
rect 52750 47170 52830 47190
rect 52860 47194 53060 47200
rect 52860 47160 52872 47194
rect 53048 47190 53060 47194
rect 53358 47194 53558 47200
rect 53358 47190 53370 47194
rect 53048 47180 53370 47190
rect 53048 47160 53180 47180
rect 52860 47154 53060 47160
rect 53170 47120 53180 47160
rect 53240 47160 53370 47180
rect 53546 47160 53558 47194
rect 53590 47190 53600 47250
rect 53660 47190 53670 47250
rect 53590 47170 53670 47190
rect 53240 47120 53250 47160
rect 53358 47154 53558 47160
rect 53170 47110 53250 47120
rect 52640 45950 52710 47100
rect 52640 45690 52660 45950
rect 52700 45690 52710 45950
rect 53720 47100 53730 47340
rect 53770 47100 53790 47340
rect 53720 45950 53790 47100
rect 53170 45920 53250 45930
rect 52860 45882 53060 45888
rect 52750 45850 52830 45870
rect 52750 45790 52760 45850
rect 52820 45838 52830 45850
rect 52860 45848 52872 45882
rect 53048 45880 53060 45882
rect 53170 45880 53180 45920
rect 53048 45860 53180 45880
rect 53240 45880 53250 45920
rect 53358 45882 53558 45888
rect 53358 45880 53370 45882
rect 53240 45860 53370 45880
rect 53048 45850 53370 45860
rect 53048 45848 53060 45850
rect 52860 45842 53060 45848
rect 53358 45848 53370 45850
rect 53546 45848 53558 45882
rect 53358 45842 53558 45848
rect 53590 45850 53670 45870
rect 52822 45804 52830 45838
rect 52820 45790 52830 45804
rect 52750 45770 52830 45790
rect 52860 45794 53060 45800
rect 52860 45760 52872 45794
rect 53048 45790 53060 45794
rect 53358 45794 53558 45800
rect 53358 45790 53370 45794
rect 53048 45760 53370 45790
rect 53546 45760 53558 45794
rect 53590 45790 53600 45850
rect 53660 45790 53670 45850
rect 53590 45770 53670 45790
rect 52860 45754 53060 45760
rect 52640 45630 52710 45690
rect 52640 45390 52660 45630
rect 52700 45390 52710 45630
rect 53170 45750 53250 45760
rect 53358 45754 53558 45760
rect 53170 45690 53180 45750
rect 53240 45690 53250 45750
rect 53170 45640 53250 45690
rect 53170 45580 53180 45640
rect 53240 45580 53250 45640
rect 52860 45572 53060 45578
rect 52750 45540 52830 45560
rect 52750 45480 52760 45540
rect 52820 45528 52830 45540
rect 52860 45538 52872 45572
rect 53048 45570 53060 45572
rect 53170 45570 53250 45580
rect 53720 45710 53730 45950
rect 53770 45710 53790 45950
rect 53720 45630 53790 45710
rect 53358 45572 53558 45578
rect 53358 45570 53370 45572
rect 53048 45540 53370 45570
rect 53048 45538 53060 45540
rect 52860 45532 53060 45538
rect 53358 45538 53370 45540
rect 53546 45538 53558 45572
rect 53358 45532 53558 45538
rect 53590 45540 53670 45560
rect 52822 45494 52830 45528
rect 52820 45480 52830 45494
rect 52750 45460 52830 45480
rect 52860 45484 53060 45490
rect 52860 45450 52872 45484
rect 53048 45480 53060 45484
rect 53358 45484 53558 45490
rect 53358 45480 53370 45484
rect 53048 45470 53370 45480
rect 53048 45450 53180 45470
rect 52860 45444 53060 45450
rect 53170 45410 53180 45450
rect 53240 45450 53370 45470
rect 53546 45450 53558 45484
rect 53590 45480 53600 45540
rect 53660 45480 53670 45540
rect 53590 45460 53670 45480
rect 53240 45410 53250 45450
rect 53358 45444 53558 45450
rect 53170 45400 53250 45410
rect 52640 44240 52710 45390
rect 52640 43980 52660 44240
rect 52700 43980 52710 44240
rect 53720 45390 53730 45630
rect 53770 45390 53790 45630
rect 53720 44240 53790 45390
rect 53170 44210 53250 44220
rect 52860 44172 53060 44178
rect 52750 44140 52830 44160
rect 52750 44080 52760 44140
rect 52820 44128 52830 44140
rect 52860 44138 52872 44172
rect 53048 44170 53060 44172
rect 53170 44170 53180 44210
rect 53048 44150 53180 44170
rect 53240 44170 53250 44210
rect 53358 44172 53558 44178
rect 53358 44170 53370 44172
rect 53240 44150 53370 44170
rect 53048 44140 53370 44150
rect 53048 44138 53060 44140
rect 52860 44132 53060 44138
rect 53358 44138 53370 44140
rect 53546 44138 53558 44172
rect 53358 44132 53558 44138
rect 53590 44140 53670 44160
rect 52822 44094 52830 44128
rect 52820 44080 52830 44094
rect 52750 44060 52830 44080
rect 52860 44084 53060 44090
rect 52860 44050 52872 44084
rect 53048 44080 53060 44084
rect 53358 44084 53558 44090
rect 53358 44080 53370 44084
rect 53048 44050 53370 44080
rect 53546 44050 53558 44084
rect 53590 44080 53600 44140
rect 53660 44080 53670 44140
rect 53590 44060 53670 44080
rect 52860 44044 53060 44050
rect 52640 43920 52710 43980
rect 52640 43680 52660 43920
rect 52700 43680 52710 43920
rect 53170 44040 53250 44050
rect 53358 44044 53558 44050
rect 53170 43980 53180 44040
rect 53240 43980 53250 44040
rect 53170 43930 53250 43980
rect 53170 43870 53180 43930
rect 53240 43870 53250 43930
rect 52860 43862 53060 43868
rect 52750 43830 52830 43850
rect 52750 43770 52760 43830
rect 52820 43818 52830 43830
rect 52860 43828 52872 43862
rect 53048 43860 53060 43862
rect 53170 43860 53250 43870
rect 53720 44000 53730 44240
rect 53770 44000 53790 44240
rect 53720 43920 53790 44000
rect 53358 43862 53558 43868
rect 53358 43860 53370 43862
rect 53048 43830 53370 43860
rect 53048 43828 53060 43830
rect 52860 43822 53060 43828
rect 53358 43828 53370 43830
rect 53546 43828 53558 43862
rect 53358 43822 53558 43828
rect 53590 43830 53670 43850
rect 52822 43784 52830 43818
rect 52820 43770 52830 43784
rect 52750 43750 52830 43770
rect 52860 43774 53060 43780
rect 52860 43740 52872 43774
rect 53048 43770 53060 43774
rect 53358 43774 53558 43780
rect 53358 43770 53370 43774
rect 53048 43760 53370 43770
rect 53048 43740 53180 43760
rect 52860 43734 53060 43740
rect 53170 43700 53180 43740
rect 53240 43740 53370 43760
rect 53546 43740 53558 43774
rect 53590 43770 53600 43830
rect 53660 43770 53670 43830
rect 53590 43750 53670 43770
rect 53240 43700 53250 43740
rect 53358 43734 53558 43740
rect 53170 43690 53250 43700
rect 52640 42530 52710 43680
rect 52640 42270 52660 42530
rect 52700 42270 52710 42530
rect 53720 43680 53730 43920
rect 53770 43680 53790 43920
rect 53720 42530 53790 43680
rect 53170 42500 53250 42510
rect 52860 42462 53060 42468
rect 52750 42430 52830 42450
rect 52750 42370 52760 42430
rect 52820 42418 52830 42430
rect 52860 42428 52872 42462
rect 53048 42460 53060 42462
rect 53170 42460 53180 42500
rect 53048 42440 53180 42460
rect 53240 42460 53250 42500
rect 53358 42462 53558 42468
rect 53358 42460 53370 42462
rect 53240 42440 53370 42460
rect 53048 42430 53370 42440
rect 53048 42428 53060 42430
rect 52860 42422 53060 42428
rect 53358 42428 53370 42430
rect 53546 42428 53558 42462
rect 53358 42422 53558 42428
rect 53590 42430 53670 42450
rect 52822 42384 52830 42418
rect 52820 42370 52830 42384
rect 52750 42350 52830 42370
rect 52860 42374 53060 42380
rect 52860 42340 52872 42374
rect 53048 42370 53060 42374
rect 53358 42374 53558 42380
rect 53358 42370 53370 42374
rect 53048 42340 53370 42370
rect 53546 42340 53558 42374
rect 53590 42370 53600 42430
rect 53660 42370 53670 42430
rect 53590 42350 53670 42370
rect 52860 42334 53060 42340
rect 52640 42210 52710 42270
rect 52640 41970 52660 42210
rect 52700 41970 52710 42210
rect 53170 42330 53250 42340
rect 53358 42334 53558 42340
rect 53170 42270 53180 42330
rect 53240 42270 53250 42330
rect 53170 42220 53250 42270
rect 53170 42160 53180 42220
rect 53240 42160 53250 42220
rect 52860 42152 53060 42158
rect 52750 42120 52830 42140
rect 52750 42060 52760 42120
rect 52820 42108 52830 42120
rect 52860 42118 52872 42152
rect 53048 42150 53060 42152
rect 53170 42150 53250 42160
rect 53720 42290 53730 42530
rect 53770 42290 53790 42530
rect 53720 42210 53790 42290
rect 53358 42152 53558 42158
rect 53358 42150 53370 42152
rect 53048 42120 53370 42150
rect 53048 42118 53060 42120
rect 52860 42112 53060 42118
rect 53358 42118 53370 42120
rect 53546 42118 53558 42152
rect 53358 42112 53558 42118
rect 53590 42120 53670 42140
rect 52822 42074 52830 42108
rect 52820 42060 52830 42074
rect 52750 42040 52830 42060
rect 52860 42064 53060 42070
rect 52860 42030 52872 42064
rect 53048 42060 53060 42064
rect 53358 42064 53558 42070
rect 53358 42060 53370 42064
rect 53048 42050 53370 42060
rect 53048 42030 53180 42050
rect 52860 42024 53060 42030
rect 53170 41990 53180 42030
rect 53240 42030 53370 42050
rect 53546 42030 53558 42064
rect 53590 42060 53600 42120
rect 53660 42060 53670 42120
rect 53590 42040 53670 42060
rect 53240 41990 53250 42030
rect 53358 42024 53558 42030
rect 53170 41980 53250 41990
rect 52640 40820 52710 41970
rect 52640 40560 52660 40820
rect 52700 40560 52710 40820
rect 53720 41970 53730 42210
rect 53770 41970 53790 42210
rect 53720 40820 53790 41970
rect 53170 40790 53250 40800
rect 52860 40752 53060 40758
rect 52750 40720 52830 40740
rect 52750 40660 52760 40720
rect 52820 40708 52830 40720
rect 52860 40718 52872 40752
rect 53048 40750 53060 40752
rect 53170 40750 53180 40790
rect 53048 40730 53180 40750
rect 53240 40750 53250 40790
rect 53358 40752 53558 40758
rect 53358 40750 53370 40752
rect 53240 40730 53370 40750
rect 53048 40720 53370 40730
rect 53048 40718 53060 40720
rect 52860 40712 53060 40718
rect 53358 40718 53370 40720
rect 53546 40718 53558 40752
rect 53358 40712 53558 40718
rect 53590 40720 53670 40740
rect 52822 40674 52830 40708
rect 52820 40660 52830 40674
rect 52750 40640 52830 40660
rect 52860 40664 53060 40670
rect 52860 40630 52872 40664
rect 53048 40660 53060 40664
rect 53358 40664 53558 40670
rect 53358 40660 53370 40664
rect 53048 40630 53370 40660
rect 53546 40630 53558 40664
rect 53590 40660 53600 40720
rect 53660 40660 53670 40720
rect 53590 40640 53670 40660
rect 52860 40624 53060 40630
rect 52640 40500 52710 40560
rect 52640 40260 52660 40500
rect 52700 40260 52710 40500
rect 53170 40620 53250 40630
rect 53358 40624 53558 40630
rect 53170 40560 53180 40620
rect 53240 40560 53250 40620
rect 53170 40510 53250 40560
rect 53170 40450 53180 40510
rect 53240 40450 53250 40510
rect 52860 40442 53060 40448
rect 52750 40410 52830 40430
rect 52750 40350 52760 40410
rect 52820 40398 52830 40410
rect 52860 40408 52872 40442
rect 53048 40440 53060 40442
rect 53170 40440 53250 40450
rect 53720 40580 53730 40820
rect 53770 40580 53790 40820
rect 53720 40500 53790 40580
rect 53358 40442 53558 40448
rect 53358 40440 53370 40442
rect 53048 40410 53370 40440
rect 53048 40408 53060 40410
rect 52860 40402 53060 40408
rect 53358 40408 53370 40410
rect 53546 40408 53558 40442
rect 53358 40402 53558 40408
rect 53590 40410 53670 40430
rect 52822 40364 52830 40398
rect 52820 40350 52830 40364
rect 52750 40330 52830 40350
rect 52860 40354 53060 40360
rect 52860 40320 52872 40354
rect 53048 40350 53060 40354
rect 53358 40354 53558 40360
rect 53358 40350 53370 40354
rect 53048 40340 53370 40350
rect 53048 40320 53180 40340
rect 52860 40314 53060 40320
rect 53170 40280 53180 40320
rect 53240 40320 53370 40340
rect 53546 40320 53558 40354
rect 53590 40350 53600 40410
rect 53660 40350 53670 40410
rect 53590 40330 53670 40350
rect 53240 40280 53250 40320
rect 53358 40314 53558 40320
rect 53170 40270 53250 40280
rect 52640 39690 52710 40260
rect 53720 40260 53730 40500
rect 53770 40260 53790 40500
rect 53720 39690 53790 40260
rect 52640 39680 52720 39690
rect 52640 39620 52650 39680
rect 52710 39620 52720 39680
rect 53710 39680 53790 39690
rect 53710 39620 53720 39680
rect 53780 39620 53790 39680
rect 53710 39610 53790 39620
rect 53820 66480 53850 67050
rect 53820 66470 53880 66480
rect 53820 66400 53880 66410
rect 53820 64770 53850 66400
rect 53910 65950 53940 67050
rect 53880 65940 53940 65950
rect 53880 65870 53940 65880
rect 53820 64760 53880 64770
rect 53820 64690 53880 64700
rect 53820 63060 53850 64690
rect 53910 64240 53940 65870
rect 53880 64230 53940 64240
rect 53880 64160 53940 64170
rect 53820 63050 53880 63060
rect 53820 62980 53880 62990
rect 53820 61350 53850 62980
rect 53910 62530 53940 64160
rect 53880 62520 53940 62530
rect 53880 62450 53940 62460
rect 53820 61340 53880 61350
rect 53820 61270 53880 61280
rect 53820 59640 53850 61270
rect 53910 60820 53940 62450
rect 53880 60810 53940 60820
rect 53880 60740 53940 60750
rect 53820 59630 53880 59640
rect 53820 59560 53880 59570
rect 53820 57930 53850 59560
rect 53910 59110 53940 60740
rect 53880 59100 53940 59110
rect 53880 59030 53940 59040
rect 53820 57920 53880 57930
rect 53820 57850 53880 57860
rect 53820 56220 53850 57850
rect 53910 57400 53940 59030
rect 53880 57390 53940 57400
rect 53880 57320 53940 57330
rect 53820 56210 53880 56220
rect 53820 56140 53880 56150
rect 53820 54510 53850 56140
rect 53910 55690 53940 57320
rect 53880 55680 53940 55690
rect 53880 55610 53940 55620
rect 53820 54500 53880 54510
rect 53820 54430 53880 54440
rect 53820 52800 53850 54430
rect 53910 53980 53940 55610
rect 53880 53970 53940 53980
rect 53880 53900 53940 53910
rect 53820 52790 53880 52800
rect 53820 52720 53880 52730
rect 53820 51090 53850 52720
rect 53910 52270 53940 53900
rect 53880 52260 53940 52270
rect 53880 52190 53940 52200
rect 53820 51080 53880 51090
rect 53820 51010 53880 51020
rect 53820 49380 53850 51010
rect 53910 50560 53940 52190
rect 53880 50550 53940 50560
rect 53880 50480 53940 50490
rect 53820 49370 53880 49380
rect 53820 49300 53880 49310
rect 53820 47670 53850 49300
rect 53910 48850 53940 50480
rect 53880 48840 53940 48850
rect 53880 48770 53940 48780
rect 53820 47660 53880 47670
rect 53820 47590 53880 47600
rect 53820 45960 53850 47590
rect 53910 47140 53940 48770
rect 53880 47130 53940 47140
rect 53880 47060 53940 47070
rect 53820 45950 53880 45960
rect 53820 45880 53880 45890
rect 53820 44250 53850 45880
rect 53910 45430 53940 47060
rect 53880 45420 53940 45430
rect 53880 45350 53940 45360
rect 53820 44240 53880 44250
rect 53820 44170 53880 44180
rect 53820 42540 53850 44170
rect 53910 43720 53940 45350
rect 53880 43710 53940 43720
rect 53880 43640 53940 43650
rect 53820 42530 53880 42540
rect 53820 42460 53880 42470
rect 53820 40830 53850 42460
rect 53910 42010 53940 43640
rect 53880 42000 53940 42010
rect 53880 41930 53940 41940
rect 53820 40820 53880 40830
rect 53820 40750 53880 40760
rect 52170 39220 52230 39230
rect 52350 39230 52610 39240
rect 49180 39160 49240 39170
rect 52410 39210 52610 39230
rect 52350 39160 52410 39170
rect 53820 38840 53850 40750
rect 53910 40300 53940 41930
rect 53880 40290 53940 40300
rect 53880 40220 53940 40230
rect 53910 39690 53940 40220
rect 53880 39680 53940 39690
rect 53880 39610 53940 39620
rect 53970 66390 54000 67050
rect 53970 66380 54030 66390
rect 53970 66310 54030 66320
rect 53970 64680 54000 66310
rect 53970 64670 54030 64680
rect 53970 64600 54030 64610
rect 53970 42450 54000 64600
rect 54090 62970 54120 67050
rect 54090 62960 54150 62970
rect 54090 62890 54150 62900
rect 54090 61250 54120 62890
rect 54090 61240 54150 61250
rect 54090 61170 54150 61180
rect 54090 45870 54120 61170
rect 54210 59550 54240 67050
rect 54210 59540 54270 59550
rect 54210 59470 54270 59480
rect 54210 47580 54240 59470
rect 54330 57840 54360 67050
rect 54330 57830 54390 57840
rect 54330 57760 54390 57770
rect 54330 56130 54360 57760
rect 54330 56120 54390 56130
rect 54330 56050 54390 56060
rect 54330 54420 54360 56050
rect 54330 54410 54390 54420
rect 54330 54340 54390 54350
rect 54330 52710 54360 54340
rect 54330 52700 54390 52710
rect 54330 52630 54390 52640
rect 54330 51000 54360 52630
rect 54330 50990 54390 51000
rect 54330 50920 54390 50930
rect 54330 49290 54360 50920
rect 54330 49280 54390 49290
rect 54330 49210 54390 49220
rect 54210 47570 54270 47580
rect 54210 47500 54270 47510
rect 54090 45860 54150 45870
rect 54090 45790 54150 45800
rect 54090 44160 54120 45790
rect 54090 44150 54150 44160
rect 54090 44080 54150 44090
rect 53970 42440 54030 42450
rect 53970 42370 54030 42380
rect 53970 40740 54000 42370
rect 53970 40730 54030 40740
rect 53970 40660 54030 40670
rect 53970 39240 54000 40660
rect 54090 39300 54120 44080
rect 54210 39360 54240 47500
rect 54330 39420 54360 49210
rect 54450 39690 54480 67050
rect 54570 39690 54600 67050
rect 54690 39690 54720 67050
rect 56850 39690 56880 67050
rect 56970 39690 57000 67050
rect 57090 39690 57120 67050
rect 57210 57840 57240 67050
rect 57330 59550 57360 67050
rect 57450 62970 57480 67050
rect 57570 66390 57600 67050
rect 57540 66380 57600 66390
rect 57540 66310 57600 66320
rect 57570 64680 57600 66310
rect 57540 64670 57600 64680
rect 57540 64600 57600 64610
rect 57420 62960 57480 62970
rect 57420 62890 57480 62900
rect 57450 61250 57480 62890
rect 57420 61240 57480 61250
rect 57420 61170 57480 61180
rect 57300 59540 57360 59550
rect 57300 59470 57360 59480
rect 57180 57830 57240 57840
rect 57180 57760 57240 57770
rect 57210 56130 57240 57760
rect 57180 56120 57240 56130
rect 57180 56050 57240 56060
rect 57210 54420 57240 56050
rect 57180 54410 57240 54420
rect 57180 54340 57240 54350
rect 57210 52710 57240 54340
rect 57180 52700 57240 52710
rect 57180 52630 57240 52640
rect 57210 51000 57240 52630
rect 57180 50990 57240 51000
rect 57180 50920 57240 50930
rect 57210 49290 57240 50920
rect 57180 49280 57240 49290
rect 57180 49210 57240 49220
rect 57210 39420 57240 49210
rect 57330 47580 57360 59470
rect 57300 47570 57360 47580
rect 57300 47500 57360 47510
rect 54330 39410 54770 39420
rect 54330 39390 54710 39410
rect 54210 39350 54590 39360
rect 54210 39330 54530 39350
rect 54090 39290 54410 39300
rect 54090 39270 54350 39290
rect 53970 39230 54230 39240
rect 53970 39210 54170 39230
rect 54710 39340 54770 39350
rect 56800 39410 57240 39420
rect 56860 39390 57240 39410
rect 57330 39360 57360 47500
rect 57450 45870 57480 61170
rect 57420 45860 57480 45870
rect 57420 45790 57480 45800
rect 57450 44160 57480 45790
rect 57420 44150 57480 44160
rect 57420 44080 57480 44090
rect 56800 39340 56860 39350
rect 56980 39350 57360 39360
rect 54530 39280 54590 39290
rect 57040 39330 57360 39350
rect 57450 39300 57480 44080
rect 57570 42450 57600 64600
rect 57540 42440 57600 42450
rect 57540 42370 57600 42380
rect 57570 40740 57600 42370
rect 57540 40730 57600 40740
rect 57540 40660 57600 40670
rect 56980 39280 57040 39290
rect 57160 39290 57480 39300
rect 54350 39220 54410 39230
rect 57220 39270 57480 39290
rect 57570 39240 57600 40660
rect 57630 66470 57700 67050
rect 57630 66210 57650 66470
rect 57690 66210 57700 66470
rect 58710 66470 58780 67050
rect 58160 66440 58240 66450
rect 57850 66402 58050 66408
rect 57740 66370 57820 66390
rect 57740 66310 57750 66370
rect 57810 66358 57820 66370
rect 57850 66368 57862 66402
rect 58038 66400 58050 66402
rect 58160 66400 58170 66440
rect 58038 66380 58170 66400
rect 58230 66400 58240 66440
rect 58348 66402 58548 66408
rect 58348 66400 58360 66402
rect 58230 66380 58360 66400
rect 58038 66370 58360 66380
rect 58038 66368 58050 66370
rect 57850 66362 58050 66368
rect 58348 66368 58360 66370
rect 58536 66368 58548 66402
rect 58348 66362 58548 66368
rect 58580 66370 58660 66390
rect 57812 66324 57820 66358
rect 57810 66310 57820 66324
rect 57740 66290 57820 66310
rect 57850 66314 58050 66320
rect 57850 66280 57862 66314
rect 58038 66310 58050 66314
rect 58348 66314 58548 66320
rect 58348 66310 58360 66314
rect 58038 66280 58360 66310
rect 58536 66280 58548 66314
rect 58580 66310 58590 66370
rect 58650 66310 58660 66370
rect 58580 66290 58660 66310
rect 57850 66274 58050 66280
rect 57630 66150 57700 66210
rect 57630 65910 57650 66150
rect 57690 65910 57700 66150
rect 58160 66270 58240 66280
rect 58348 66274 58548 66280
rect 58160 66210 58170 66270
rect 58230 66210 58240 66270
rect 58160 66160 58240 66210
rect 58160 66100 58170 66160
rect 58230 66100 58240 66160
rect 57850 66092 58050 66098
rect 57740 66060 57820 66080
rect 57740 66000 57750 66060
rect 57810 66048 57820 66060
rect 57850 66058 57862 66092
rect 58038 66090 58050 66092
rect 58160 66090 58240 66100
rect 58710 66230 58720 66470
rect 58760 66230 58780 66470
rect 58710 66150 58780 66230
rect 58348 66092 58548 66098
rect 58348 66090 58360 66092
rect 58038 66060 58360 66090
rect 58038 66058 58050 66060
rect 57850 66052 58050 66058
rect 58348 66058 58360 66060
rect 58536 66058 58548 66092
rect 58348 66052 58548 66058
rect 58580 66060 58660 66080
rect 57812 66014 57820 66048
rect 57810 66000 57820 66014
rect 57740 65980 57820 66000
rect 57850 66004 58050 66010
rect 57850 65970 57862 66004
rect 58038 66000 58050 66004
rect 58348 66004 58548 66010
rect 58348 66000 58360 66004
rect 58038 65990 58360 66000
rect 58038 65970 58170 65990
rect 57850 65964 58050 65970
rect 58160 65930 58170 65970
rect 58230 65970 58360 65990
rect 58536 65970 58548 66004
rect 58580 66000 58590 66060
rect 58650 66000 58660 66060
rect 58580 65980 58660 66000
rect 58230 65930 58240 65970
rect 58348 65964 58548 65970
rect 58160 65920 58240 65930
rect 57630 64760 57700 65910
rect 57630 64500 57650 64760
rect 57690 64500 57700 64760
rect 58710 65910 58720 66150
rect 58760 65910 58780 66150
rect 58710 64760 58780 65910
rect 58160 64730 58240 64740
rect 57850 64692 58050 64698
rect 57740 64660 57820 64680
rect 57740 64600 57750 64660
rect 57810 64648 57820 64660
rect 57850 64658 57862 64692
rect 58038 64690 58050 64692
rect 58160 64690 58170 64730
rect 58038 64670 58170 64690
rect 58230 64690 58240 64730
rect 58348 64692 58548 64698
rect 58348 64690 58360 64692
rect 58230 64670 58360 64690
rect 58038 64660 58360 64670
rect 58038 64658 58050 64660
rect 57850 64652 58050 64658
rect 58348 64658 58360 64660
rect 58536 64658 58548 64692
rect 58348 64652 58548 64658
rect 58580 64660 58660 64680
rect 57812 64614 57820 64648
rect 57810 64600 57820 64614
rect 57740 64580 57820 64600
rect 57850 64604 58050 64610
rect 57850 64570 57862 64604
rect 58038 64600 58050 64604
rect 58348 64604 58548 64610
rect 58348 64600 58360 64604
rect 58038 64570 58360 64600
rect 58536 64570 58548 64604
rect 58580 64600 58590 64660
rect 58650 64600 58660 64660
rect 58580 64580 58660 64600
rect 57850 64564 58050 64570
rect 57630 64440 57700 64500
rect 57630 64200 57650 64440
rect 57690 64200 57700 64440
rect 58160 64560 58240 64570
rect 58348 64564 58548 64570
rect 58160 64500 58170 64560
rect 58230 64500 58240 64560
rect 58160 64450 58240 64500
rect 58160 64390 58170 64450
rect 58230 64390 58240 64450
rect 57850 64382 58050 64388
rect 57740 64350 57820 64370
rect 57740 64290 57750 64350
rect 57810 64338 57820 64350
rect 57850 64348 57862 64382
rect 58038 64380 58050 64382
rect 58160 64380 58240 64390
rect 58710 64520 58720 64760
rect 58760 64520 58780 64760
rect 58710 64440 58780 64520
rect 58348 64382 58548 64388
rect 58348 64380 58360 64382
rect 58038 64350 58360 64380
rect 58038 64348 58050 64350
rect 57850 64342 58050 64348
rect 58348 64348 58360 64350
rect 58536 64348 58548 64382
rect 58348 64342 58548 64348
rect 58580 64350 58660 64370
rect 57812 64304 57820 64338
rect 57810 64290 57820 64304
rect 57740 64270 57820 64290
rect 57850 64294 58050 64300
rect 57850 64260 57862 64294
rect 58038 64290 58050 64294
rect 58348 64294 58548 64300
rect 58348 64290 58360 64294
rect 58038 64280 58360 64290
rect 58038 64260 58170 64280
rect 57850 64254 58050 64260
rect 58160 64220 58170 64260
rect 58230 64260 58360 64280
rect 58536 64260 58548 64294
rect 58580 64290 58590 64350
rect 58650 64290 58660 64350
rect 58580 64270 58660 64290
rect 58230 64220 58240 64260
rect 58348 64254 58548 64260
rect 58160 64210 58240 64220
rect 57630 63050 57700 64200
rect 57630 62790 57650 63050
rect 57690 62790 57700 63050
rect 58710 64200 58720 64440
rect 58760 64200 58780 64440
rect 58710 63050 58780 64200
rect 58160 63020 58240 63030
rect 57850 62982 58050 62988
rect 57740 62950 57820 62970
rect 57740 62890 57750 62950
rect 57810 62938 57820 62950
rect 57850 62948 57862 62982
rect 58038 62980 58050 62982
rect 58160 62980 58170 63020
rect 58038 62960 58170 62980
rect 58230 62980 58240 63020
rect 58348 62982 58548 62988
rect 58348 62980 58360 62982
rect 58230 62960 58360 62980
rect 58038 62950 58360 62960
rect 58038 62948 58050 62950
rect 57850 62942 58050 62948
rect 58348 62948 58360 62950
rect 58536 62948 58548 62982
rect 58348 62942 58548 62948
rect 58580 62950 58660 62970
rect 57812 62904 57820 62938
rect 57810 62890 57820 62904
rect 57740 62870 57820 62890
rect 57850 62894 58050 62900
rect 57850 62860 57862 62894
rect 58038 62890 58050 62894
rect 58348 62894 58548 62900
rect 58348 62890 58360 62894
rect 58038 62860 58360 62890
rect 58536 62860 58548 62894
rect 58580 62890 58590 62950
rect 58650 62890 58660 62950
rect 58580 62870 58660 62890
rect 57850 62854 58050 62860
rect 57630 62730 57700 62790
rect 57630 62490 57650 62730
rect 57690 62490 57700 62730
rect 58160 62850 58240 62860
rect 58348 62854 58548 62860
rect 58160 62790 58170 62850
rect 58230 62790 58240 62850
rect 58160 62740 58240 62790
rect 58160 62680 58170 62740
rect 58230 62680 58240 62740
rect 57850 62672 58050 62678
rect 57740 62640 57820 62660
rect 57740 62580 57750 62640
rect 57810 62628 57820 62640
rect 57850 62638 57862 62672
rect 58038 62670 58050 62672
rect 58160 62670 58240 62680
rect 58710 62810 58720 63050
rect 58760 62810 58780 63050
rect 58710 62730 58780 62810
rect 58348 62672 58548 62678
rect 58348 62670 58360 62672
rect 58038 62640 58360 62670
rect 58038 62638 58050 62640
rect 57850 62632 58050 62638
rect 58348 62638 58360 62640
rect 58536 62638 58548 62672
rect 58348 62632 58548 62638
rect 58580 62640 58660 62660
rect 57812 62594 57820 62628
rect 57810 62580 57820 62594
rect 57740 62560 57820 62580
rect 57850 62584 58050 62590
rect 57850 62550 57862 62584
rect 58038 62580 58050 62584
rect 58348 62584 58548 62590
rect 58348 62580 58360 62584
rect 58038 62570 58360 62580
rect 58038 62550 58170 62570
rect 57850 62544 58050 62550
rect 58160 62510 58170 62550
rect 58230 62550 58360 62570
rect 58536 62550 58548 62584
rect 58580 62580 58590 62640
rect 58650 62580 58660 62640
rect 58580 62560 58660 62580
rect 58230 62510 58240 62550
rect 58348 62544 58548 62550
rect 58160 62500 58240 62510
rect 57630 61340 57700 62490
rect 57630 61080 57650 61340
rect 57690 61080 57700 61340
rect 58710 62490 58720 62730
rect 58760 62490 58780 62730
rect 58710 61340 58780 62490
rect 58160 61310 58240 61320
rect 57850 61272 58050 61278
rect 57740 61240 57820 61260
rect 57740 61180 57750 61240
rect 57810 61228 57820 61240
rect 57850 61238 57862 61272
rect 58038 61270 58050 61272
rect 58160 61270 58170 61310
rect 58038 61250 58170 61270
rect 58230 61270 58240 61310
rect 58348 61272 58548 61278
rect 58348 61270 58360 61272
rect 58230 61250 58360 61270
rect 58038 61240 58360 61250
rect 58038 61238 58050 61240
rect 57850 61232 58050 61238
rect 58348 61238 58360 61240
rect 58536 61238 58548 61272
rect 58348 61232 58548 61238
rect 58580 61240 58660 61260
rect 57812 61194 57820 61228
rect 57810 61180 57820 61194
rect 57740 61160 57820 61180
rect 57850 61184 58050 61190
rect 57850 61150 57862 61184
rect 58038 61180 58050 61184
rect 58348 61184 58548 61190
rect 58348 61180 58360 61184
rect 58038 61150 58360 61180
rect 58536 61150 58548 61184
rect 58580 61180 58590 61240
rect 58650 61180 58660 61240
rect 58580 61160 58660 61180
rect 57850 61144 58050 61150
rect 57630 61020 57700 61080
rect 57630 60780 57650 61020
rect 57690 60780 57700 61020
rect 58160 61140 58240 61150
rect 58348 61144 58548 61150
rect 58160 61080 58170 61140
rect 58230 61080 58240 61140
rect 58160 61030 58240 61080
rect 58160 60970 58170 61030
rect 58230 60970 58240 61030
rect 57850 60962 58050 60968
rect 57740 60930 57820 60950
rect 57740 60870 57750 60930
rect 57810 60918 57820 60930
rect 57850 60928 57862 60962
rect 58038 60960 58050 60962
rect 58160 60960 58240 60970
rect 58710 61100 58720 61340
rect 58760 61100 58780 61340
rect 58710 61020 58780 61100
rect 58348 60962 58548 60968
rect 58348 60960 58360 60962
rect 58038 60930 58360 60960
rect 58038 60928 58050 60930
rect 57850 60922 58050 60928
rect 58348 60928 58360 60930
rect 58536 60928 58548 60962
rect 58348 60922 58548 60928
rect 58580 60930 58660 60950
rect 57812 60884 57820 60918
rect 57810 60870 57820 60884
rect 57740 60850 57820 60870
rect 57850 60874 58050 60880
rect 57850 60840 57862 60874
rect 58038 60870 58050 60874
rect 58348 60874 58548 60880
rect 58348 60870 58360 60874
rect 58038 60860 58360 60870
rect 58038 60840 58170 60860
rect 57850 60834 58050 60840
rect 58160 60800 58170 60840
rect 58230 60840 58360 60860
rect 58536 60840 58548 60874
rect 58580 60870 58590 60930
rect 58650 60870 58660 60930
rect 58580 60850 58660 60870
rect 58230 60800 58240 60840
rect 58348 60834 58548 60840
rect 58160 60790 58240 60800
rect 57630 59630 57700 60780
rect 57630 59370 57650 59630
rect 57690 59370 57700 59630
rect 58710 60780 58720 61020
rect 58760 60780 58780 61020
rect 58710 59630 58780 60780
rect 58160 59600 58240 59610
rect 57850 59562 58050 59568
rect 57740 59530 57820 59550
rect 57740 59470 57750 59530
rect 57810 59518 57820 59530
rect 57850 59528 57862 59562
rect 58038 59560 58050 59562
rect 58160 59560 58170 59600
rect 58038 59540 58170 59560
rect 58230 59560 58240 59600
rect 58348 59562 58548 59568
rect 58348 59560 58360 59562
rect 58230 59540 58360 59560
rect 58038 59530 58360 59540
rect 58038 59528 58050 59530
rect 57850 59522 58050 59528
rect 58348 59528 58360 59530
rect 58536 59528 58548 59562
rect 58348 59522 58548 59528
rect 58580 59530 58660 59550
rect 57812 59484 57820 59518
rect 57810 59470 57820 59484
rect 57740 59450 57820 59470
rect 57850 59474 58050 59480
rect 57850 59440 57862 59474
rect 58038 59470 58050 59474
rect 58348 59474 58548 59480
rect 58348 59470 58360 59474
rect 58038 59440 58360 59470
rect 58536 59440 58548 59474
rect 58580 59470 58590 59530
rect 58650 59470 58660 59530
rect 58580 59450 58660 59470
rect 57850 59434 58050 59440
rect 57630 59310 57700 59370
rect 57630 59070 57650 59310
rect 57690 59070 57700 59310
rect 58160 59430 58240 59440
rect 58348 59434 58548 59440
rect 58160 59370 58170 59430
rect 58230 59370 58240 59430
rect 58160 59320 58240 59370
rect 58160 59260 58170 59320
rect 58230 59260 58240 59320
rect 57850 59252 58050 59258
rect 57740 59220 57820 59240
rect 57740 59160 57750 59220
rect 57810 59208 57820 59220
rect 57850 59218 57862 59252
rect 58038 59250 58050 59252
rect 58160 59250 58240 59260
rect 58710 59390 58720 59630
rect 58760 59390 58780 59630
rect 58710 59310 58780 59390
rect 58348 59252 58548 59258
rect 58348 59250 58360 59252
rect 58038 59220 58360 59250
rect 58038 59218 58050 59220
rect 57850 59212 58050 59218
rect 58348 59218 58360 59220
rect 58536 59218 58548 59252
rect 58348 59212 58548 59218
rect 58580 59220 58660 59240
rect 57812 59174 57820 59208
rect 57810 59160 57820 59174
rect 57740 59140 57820 59160
rect 57850 59164 58050 59170
rect 57850 59130 57862 59164
rect 58038 59160 58050 59164
rect 58348 59164 58548 59170
rect 58348 59160 58360 59164
rect 58038 59150 58360 59160
rect 58038 59130 58170 59150
rect 57850 59124 58050 59130
rect 58160 59090 58170 59130
rect 58230 59130 58360 59150
rect 58536 59130 58548 59164
rect 58580 59160 58590 59220
rect 58650 59160 58660 59220
rect 58580 59140 58660 59160
rect 58230 59090 58240 59130
rect 58348 59124 58548 59130
rect 58160 59080 58240 59090
rect 57630 57920 57700 59070
rect 57630 57660 57650 57920
rect 57690 57660 57700 57920
rect 58710 59070 58720 59310
rect 58760 59070 58780 59310
rect 58710 57920 58780 59070
rect 58160 57890 58240 57900
rect 57850 57852 58050 57858
rect 57740 57820 57820 57840
rect 57740 57760 57750 57820
rect 57810 57808 57820 57820
rect 57850 57818 57862 57852
rect 58038 57850 58050 57852
rect 58160 57850 58170 57890
rect 58038 57830 58170 57850
rect 58230 57850 58240 57890
rect 58348 57852 58548 57858
rect 58348 57850 58360 57852
rect 58230 57830 58360 57850
rect 58038 57820 58360 57830
rect 58038 57818 58050 57820
rect 57850 57812 58050 57818
rect 58348 57818 58360 57820
rect 58536 57818 58548 57852
rect 58348 57812 58548 57818
rect 58580 57820 58660 57840
rect 57812 57774 57820 57808
rect 57810 57760 57820 57774
rect 57740 57740 57820 57760
rect 57850 57764 58050 57770
rect 57850 57730 57862 57764
rect 58038 57760 58050 57764
rect 58348 57764 58548 57770
rect 58348 57760 58360 57764
rect 58038 57730 58360 57760
rect 58536 57730 58548 57764
rect 58580 57760 58590 57820
rect 58650 57760 58660 57820
rect 58580 57740 58660 57760
rect 57850 57724 58050 57730
rect 57630 57600 57700 57660
rect 57630 57360 57650 57600
rect 57690 57360 57700 57600
rect 58160 57720 58240 57730
rect 58348 57724 58548 57730
rect 58160 57660 58170 57720
rect 58230 57660 58240 57720
rect 58160 57610 58240 57660
rect 58160 57550 58170 57610
rect 58230 57550 58240 57610
rect 57850 57542 58050 57548
rect 57740 57510 57820 57530
rect 57740 57450 57750 57510
rect 57810 57498 57820 57510
rect 57850 57508 57862 57542
rect 58038 57540 58050 57542
rect 58160 57540 58240 57550
rect 58710 57680 58720 57920
rect 58760 57680 58780 57920
rect 58710 57600 58780 57680
rect 58348 57542 58548 57548
rect 58348 57540 58360 57542
rect 58038 57510 58360 57540
rect 58038 57508 58050 57510
rect 57850 57502 58050 57508
rect 58348 57508 58360 57510
rect 58536 57508 58548 57542
rect 58348 57502 58548 57508
rect 58580 57510 58660 57530
rect 57812 57464 57820 57498
rect 57810 57450 57820 57464
rect 57740 57430 57820 57450
rect 57850 57454 58050 57460
rect 57850 57420 57862 57454
rect 58038 57450 58050 57454
rect 58348 57454 58548 57460
rect 58348 57450 58360 57454
rect 58038 57440 58360 57450
rect 58038 57420 58170 57440
rect 57850 57414 58050 57420
rect 58160 57380 58170 57420
rect 58230 57420 58360 57440
rect 58536 57420 58548 57454
rect 58580 57450 58590 57510
rect 58650 57450 58660 57510
rect 58580 57430 58660 57450
rect 58230 57380 58240 57420
rect 58348 57414 58548 57420
rect 58160 57370 58240 57380
rect 57630 56210 57700 57360
rect 57630 55950 57650 56210
rect 57690 55950 57700 56210
rect 58710 57360 58720 57600
rect 58760 57360 58780 57600
rect 58710 56210 58780 57360
rect 58160 56180 58240 56190
rect 57850 56142 58050 56148
rect 57740 56110 57820 56130
rect 57740 56050 57750 56110
rect 57810 56098 57820 56110
rect 57850 56108 57862 56142
rect 58038 56140 58050 56142
rect 58160 56140 58170 56180
rect 58038 56120 58170 56140
rect 58230 56140 58240 56180
rect 58348 56142 58548 56148
rect 58348 56140 58360 56142
rect 58230 56120 58360 56140
rect 58038 56110 58360 56120
rect 58038 56108 58050 56110
rect 57850 56102 58050 56108
rect 58348 56108 58360 56110
rect 58536 56108 58548 56142
rect 58348 56102 58548 56108
rect 58580 56110 58660 56130
rect 57812 56064 57820 56098
rect 57810 56050 57820 56064
rect 57740 56030 57820 56050
rect 57850 56054 58050 56060
rect 57850 56020 57862 56054
rect 58038 56050 58050 56054
rect 58348 56054 58548 56060
rect 58348 56050 58360 56054
rect 58038 56020 58360 56050
rect 58536 56020 58548 56054
rect 58580 56050 58590 56110
rect 58650 56050 58660 56110
rect 58580 56030 58660 56050
rect 57850 56014 58050 56020
rect 57630 55890 57700 55950
rect 57630 55650 57650 55890
rect 57690 55650 57700 55890
rect 58160 56010 58240 56020
rect 58348 56014 58548 56020
rect 58160 55950 58170 56010
rect 58230 55950 58240 56010
rect 58160 55900 58240 55950
rect 58160 55840 58170 55900
rect 58230 55840 58240 55900
rect 57850 55832 58050 55838
rect 57740 55800 57820 55820
rect 57740 55740 57750 55800
rect 57810 55788 57820 55800
rect 57850 55798 57862 55832
rect 58038 55830 58050 55832
rect 58160 55830 58240 55840
rect 58710 55970 58720 56210
rect 58760 55970 58780 56210
rect 58710 55890 58780 55970
rect 58348 55832 58548 55838
rect 58348 55830 58360 55832
rect 58038 55800 58360 55830
rect 58038 55798 58050 55800
rect 57850 55792 58050 55798
rect 58348 55798 58360 55800
rect 58536 55798 58548 55832
rect 58348 55792 58548 55798
rect 58580 55800 58660 55820
rect 57812 55754 57820 55788
rect 57810 55740 57820 55754
rect 57740 55720 57820 55740
rect 57850 55744 58050 55750
rect 57850 55710 57862 55744
rect 58038 55740 58050 55744
rect 58348 55744 58548 55750
rect 58348 55740 58360 55744
rect 58038 55730 58360 55740
rect 58038 55710 58170 55730
rect 57850 55704 58050 55710
rect 58160 55670 58170 55710
rect 58230 55710 58360 55730
rect 58536 55710 58548 55744
rect 58580 55740 58590 55800
rect 58650 55740 58660 55800
rect 58580 55720 58660 55740
rect 58230 55670 58240 55710
rect 58348 55704 58548 55710
rect 58160 55660 58240 55670
rect 57630 54500 57700 55650
rect 57630 54240 57650 54500
rect 57690 54240 57700 54500
rect 58710 55650 58720 55890
rect 58760 55650 58780 55890
rect 58710 54500 58780 55650
rect 58160 54470 58240 54480
rect 57850 54432 58050 54438
rect 57740 54400 57820 54420
rect 57740 54340 57750 54400
rect 57810 54388 57820 54400
rect 57850 54398 57862 54432
rect 58038 54430 58050 54432
rect 58160 54430 58170 54470
rect 58038 54410 58170 54430
rect 58230 54430 58240 54470
rect 58348 54432 58548 54438
rect 58348 54430 58360 54432
rect 58230 54410 58360 54430
rect 58038 54400 58360 54410
rect 58038 54398 58050 54400
rect 57850 54392 58050 54398
rect 58348 54398 58360 54400
rect 58536 54398 58548 54432
rect 58348 54392 58548 54398
rect 58580 54400 58660 54420
rect 57812 54354 57820 54388
rect 57810 54340 57820 54354
rect 57740 54320 57820 54340
rect 57850 54344 58050 54350
rect 57850 54310 57862 54344
rect 58038 54340 58050 54344
rect 58348 54344 58548 54350
rect 58348 54340 58360 54344
rect 58038 54310 58360 54340
rect 58536 54310 58548 54344
rect 58580 54340 58590 54400
rect 58650 54340 58660 54400
rect 58580 54320 58660 54340
rect 57850 54304 58050 54310
rect 57630 54180 57700 54240
rect 57630 53940 57650 54180
rect 57690 53940 57700 54180
rect 58160 54300 58240 54310
rect 58348 54304 58548 54310
rect 58160 54240 58170 54300
rect 58230 54240 58240 54300
rect 58160 54190 58240 54240
rect 58160 54130 58170 54190
rect 58230 54130 58240 54190
rect 57850 54122 58050 54128
rect 57740 54090 57820 54110
rect 57740 54030 57750 54090
rect 57810 54078 57820 54090
rect 57850 54088 57862 54122
rect 58038 54120 58050 54122
rect 58160 54120 58240 54130
rect 58710 54260 58720 54500
rect 58760 54260 58780 54500
rect 58710 54180 58780 54260
rect 58348 54122 58548 54128
rect 58348 54120 58360 54122
rect 58038 54090 58360 54120
rect 58038 54088 58050 54090
rect 57850 54082 58050 54088
rect 58348 54088 58360 54090
rect 58536 54088 58548 54122
rect 58348 54082 58548 54088
rect 58580 54090 58660 54110
rect 57812 54044 57820 54078
rect 57810 54030 57820 54044
rect 57740 54010 57820 54030
rect 57850 54034 58050 54040
rect 57850 54000 57862 54034
rect 58038 54030 58050 54034
rect 58348 54034 58548 54040
rect 58348 54030 58360 54034
rect 58038 54020 58360 54030
rect 58038 54000 58170 54020
rect 57850 53994 58050 54000
rect 58160 53960 58170 54000
rect 58230 54000 58360 54020
rect 58536 54000 58548 54034
rect 58580 54030 58590 54090
rect 58650 54030 58660 54090
rect 58580 54010 58660 54030
rect 58230 53960 58240 54000
rect 58348 53994 58548 54000
rect 58160 53950 58240 53960
rect 57630 52790 57700 53940
rect 57630 52530 57650 52790
rect 57690 52530 57700 52790
rect 58710 53940 58720 54180
rect 58760 53940 58780 54180
rect 58710 52790 58780 53940
rect 58160 52760 58240 52770
rect 57850 52722 58050 52728
rect 57740 52690 57820 52710
rect 57740 52630 57750 52690
rect 57810 52678 57820 52690
rect 57850 52688 57862 52722
rect 58038 52720 58050 52722
rect 58160 52720 58170 52760
rect 58038 52700 58170 52720
rect 58230 52720 58240 52760
rect 58348 52722 58548 52728
rect 58348 52720 58360 52722
rect 58230 52700 58360 52720
rect 58038 52690 58360 52700
rect 58038 52688 58050 52690
rect 57850 52682 58050 52688
rect 58348 52688 58360 52690
rect 58536 52688 58548 52722
rect 58348 52682 58548 52688
rect 58580 52690 58660 52710
rect 57812 52644 57820 52678
rect 57810 52630 57820 52644
rect 57740 52610 57820 52630
rect 57850 52634 58050 52640
rect 57850 52600 57862 52634
rect 58038 52630 58050 52634
rect 58348 52634 58548 52640
rect 58348 52630 58360 52634
rect 58038 52600 58360 52630
rect 58536 52600 58548 52634
rect 58580 52630 58590 52690
rect 58650 52630 58660 52690
rect 58580 52610 58660 52630
rect 57850 52594 58050 52600
rect 57630 52470 57700 52530
rect 57630 52230 57650 52470
rect 57690 52230 57700 52470
rect 58160 52590 58240 52600
rect 58348 52594 58548 52600
rect 58160 52530 58170 52590
rect 58230 52530 58240 52590
rect 58160 52480 58240 52530
rect 58160 52420 58170 52480
rect 58230 52420 58240 52480
rect 57850 52412 58050 52418
rect 57740 52380 57820 52400
rect 57740 52320 57750 52380
rect 57810 52368 57820 52380
rect 57850 52378 57862 52412
rect 58038 52410 58050 52412
rect 58160 52410 58240 52420
rect 58710 52550 58720 52790
rect 58760 52550 58780 52790
rect 58710 52470 58780 52550
rect 58348 52412 58548 52418
rect 58348 52410 58360 52412
rect 58038 52380 58360 52410
rect 58038 52378 58050 52380
rect 57850 52372 58050 52378
rect 58348 52378 58360 52380
rect 58536 52378 58548 52412
rect 58348 52372 58548 52378
rect 58580 52380 58660 52400
rect 57812 52334 57820 52368
rect 57810 52320 57820 52334
rect 57740 52300 57820 52320
rect 57850 52324 58050 52330
rect 57850 52290 57862 52324
rect 58038 52320 58050 52324
rect 58348 52324 58548 52330
rect 58348 52320 58360 52324
rect 58038 52310 58360 52320
rect 58038 52290 58170 52310
rect 57850 52284 58050 52290
rect 58160 52250 58170 52290
rect 58230 52290 58360 52310
rect 58536 52290 58548 52324
rect 58580 52320 58590 52380
rect 58650 52320 58660 52380
rect 58580 52300 58660 52320
rect 58230 52250 58240 52290
rect 58348 52284 58548 52290
rect 58160 52240 58240 52250
rect 57630 51080 57700 52230
rect 57630 50820 57650 51080
rect 57690 50820 57700 51080
rect 58710 52230 58720 52470
rect 58760 52230 58780 52470
rect 58710 51080 58780 52230
rect 58160 51050 58240 51060
rect 57850 51012 58050 51018
rect 57740 50980 57820 51000
rect 57740 50920 57750 50980
rect 57810 50968 57820 50980
rect 57850 50978 57862 51012
rect 58038 51010 58050 51012
rect 58160 51010 58170 51050
rect 58038 50990 58170 51010
rect 58230 51010 58240 51050
rect 58348 51012 58548 51018
rect 58348 51010 58360 51012
rect 58230 50990 58360 51010
rect 58038 50980 58360 50990
rect 58038 50978 58050 50980
rect 57850 50972 58050 50978
rect 58348 50978 58360 50980
rect 58536 50978 58548 51012
rect 58348 50972 58548 50978
rect 58580 50980 58660 51000
rect 57812 50934 57820 50968
rect 57810 50920 57820 50934
rect 57740 50900 57820 50920
rect 57850 50924 58050 50930
rect 57850 50890 57862 50924
rect 58038 50920 58050 50924
rect 58348 50924 58548 50930
rect 58348 50920 58360 50924
rect 58038 50890 58360 50920
rect 58536 50890 58548 50924
rect 58580 50920 58590 50980
rect 58650 50920 58660 50980
rect 58580 50900 58660 50920
rect 57850 50884 58050 50890
rect 57630 50760 57700 50820
rect 57630 50520 57650 50760
rect 57690 50520 57700 50760
rect 58160 50880 58240 50890
rect 58348 50884 58548 50890
rect 58160 50820 58170 50880
rect 58230 50820 58240 50880
rect 58160 50770 58240 50820
rect 58160 50710 58170 50770
rect 58230 50710 58240 50770
rect 57850 50702 58050 50708
rect 57740 50670 57820 50690
rect 57740 50610 57750 50670
rect 57810 50658 57820 50670
rect 57850 50668 57862 50702
rect 58038 50700 58050 50702
rect 58160 50700 58240 50710
rect 58710 50840 58720 51080
rect 58760 50840 58780 51080
rect 58710 50760 58780 50840
rect 58348 50702 58548 50708
rect 58348 50700 58360 50702
rect 58038 50670 58360 50700
rect 58038 50668 58050 50670
rect 57850 50662 58050 50668
rect 58348 50668 58360 50670
rect 58536 50668 58548 50702
rect 58348 50662 58548 50668
rect 58580 50670 58660 50690
rect 57812 50624 57820 50658
rect 57810 50610 57820 50624
rect 57740 50590 57820 50610
rect 57850 50614 58050 50620
rect 57850 50580 57862 50614
rect 58038 50610 58050 50614
rect 58348 50614 58548 50620
rect 58348 50610 58360 50614
rect 58038 50600 58360 50610
rect 58038 50580 58170 50600
rect 57850 50574 58050 50580
rect 58160 50540 58170 50580
rect 58230 50580 58360 50600
rect 58536 50580 58548 50614
rect 58580 50610 58590 50670
rect 58650 50610 58660 50670
rect 58580 50590 58660 50610
rect 58230 50540 58240 50580
rect 58348 50574 58548 50580
rect 58160 50530 58240 50540
rect 57630 49370 57700 50520
rect 57630 49110 57650 49370
rect 57690 49110 57700 49370
rect 58710 50520 58720 50760
rect 58760 50520 58780 50760
rect 58710 49370 58780 50520
rect 58160 49340 58240 49350
rect 57850 49302 58050 49308
rect 57740 49270 57820 49290
rect 57740 49210 57750 49270
rect 57810 49258 57820 49270
rect 57850 49268 57862 49302
rect 58038 49300 58050 49302
rect 58160 49300 58170 49340
rect 58038 49280 58170 49300
rect 58230 49300 58240 49340
rect 58348 49302 58548 49308
rect 58348 49300 58360 49302
rect 58230 49280 58360 49300
rect 58038 49270 58360 49280
rect 58038 49268 58050 49270
rect 57850 49262 58050 49268
rect 58348 49268 58360 49270
rect 58536 49268 58548 49302
rect 58348 49262 58548 49268
rect 58580 49270 58660 49290
rect 57812 49224 57820 49258
rect 57810 49210 57820 49224
rect 57740 49190 57820 49210
rect 57850 49214 58050 49220
rect 57850 49180 57862 49214
rect 58038 49210 58050 49214
rect 58348 49214 58548 49220
rect 58348 49210 58360 49214
rect 58038 49180 58360 49210
rect 58536 49180 58548 49214
rect 58580 49210 58590 49270
rect 58650 49210 58660 49270
rect 58580 49190 58660 49210
rect 57850 49174 58050 49180
rect 57630 49050 57700 49110
rect 57630 48810 57650 49050
rect 57690 48810 57700 49050
rect 58160 49170 58240 49180
rect 58348 49174 58548 49180
rect 58160 49110 58170 49170
rect 58230 49110 58240 49170
rect 58160 49060 58240 49110
rect 58160 49000 58170 49060
rect 58230 49000 58240 49060
rect 57850 48992 58050 48998
rect 57740 48960 57820 48980
rect 57740 48900 57750 48960
rect 57810 48948 57820 48960
rect 57850 48958 57862 48992
rect 58038 48990 58050 48992
rect 58160 48990 58240 49000
rect 58710 49130 58720 49370
rect 58760 49130 58780 49370
rect 58710 49050 58780 49130
rect 58348 48992 58548 48998
rect 58348 48990 58360 48992
rect 58038 48960 58360 48990
rect 58038 48958 58050 48960
rect 57850 48952 58050 48958
rect 58348 48958 58360 48960
rect 58536 48958 58548 48992
rect 58348 48952 58548 48958
rect 58580 48960 58660 48980
rect 57812 48914 57820 48948
rect 57810 48900 57820 48914
rect 57740 48880 57820 48900
rect 57850 48904 58050 48910
rect 57850 48870 57862 48904
rect 58038 48900 58050 48904
rect 58348 48904 58548 48910
rect 58348 48900 58360 48904
rect 58038 48890 58360 48900
rect 58038 48870 58170 48890
rect 57850 48864 58050 48870
rect 58160 48830 58170 48870
rect 58230 48870 58360 48890
rect 58536 48870 58548 48904
rect 58580 48900 58590 48960
rect 58650 48900 58660 48960
rect 58580 48880 58660 48900
rect 58230 48830 58240 48870
rect 58348 48864 58548 48870
rect 58160 48820 58240 48830
rect 57630 47660 57700 48810
rect 57630 47400 57650 47660
rect 57690 47400 57700 47660
rect 58710 48810 58720 49050
rect 58760 48810 58780 49050
rect 58710 47660 58780 48810
rect 58160 47630 58240 47640
rect 57850 47592 58050 47598
rect 57740 47560 57820 47580
rect 57740 47500 57750 47560
rect 57810 47548 57820 47560
rect 57850 47558 57862 47592
rect 58038 47590 58050 47592
rect 58160 47590 58170 47630
rect 58038 47570 58170 47590
rect 58230 47590 58240 47630
rect 58348 47592 58548 47598
rect 58348 47590 58360 47592
rect 58230 47570 58360 47590
rect 58038 47560 58360 47570
rect 58038 47558 58050 47560
rect 57850 47552 58050 47558
rect 58348 47558 58360 47560
rect 58536 47558 58548 47592
rect 58348 47552 58548 47558
rect 58580 47560 58660 47580
rect 57812 47514 57820 47548
rect 57810 47500 57820 47514
rect 57740 47480 57820 47500
rect 57850 47504 58050 47510
rect 57850 47470 57862 47504
rect 58038 47500 58050 47504
rect 58348 47504 58548 47510
rect 58348 47500 58360 47504
rect 58038 47470 58360 47500
rect 58536 47470 58548 47504
rect 58580 47500 58590 47560
rect 58650 47500 58660 47560
rect 58580 47480 58660 47500
rect 57850 47464 58050 47470
rect 57630 47340 57700 47400
rect 57630 47100 57650 47340
rect 57690 47100 57700 47340
rect 58160 47460 58240 47470
rect 58348 47464 58548 47470
rect 58160 47400 58170 47460
rect 58230 47400 58240 47460
rect 58160 47350 58240 47400
rect 58160 47290 58170 47350
rect 58230 47290 58240 47350
rect 57850 47282 58050 47288
rect 57740 47250 57820 47270
rect 57740 47190 57750 47250
rect 57810 47238 57820 47250
rect 57850 47248 57862 47282
rect 58038 47280 58050 47282
rect 58160 47280 58240 47290
rect 58710 47420 58720 47660
rect 58760 47420 58780 47660
rect 58710 47340 58780 47420
rect 58348 47282 58548 47288
rect 58348 47280 58360 47282
rect 58038 47250 58360 47280
rect 58038 47248 58050 47250
rect 57850 47242 58050 47248
rect 58348 47248 58360 47250
rect 58536 47248 58548 47282
rect 58348 47242 58548 47248
rect 58580 47250 58660 47270
rect 57812 47204 57820 47238
rect 57810 47190 57820 47204
rect 57740 47170 57820 47190
rect 57850 47194 58050 47200
rect 57850 47160 57862 47194
rect 58038 47190 58050 47194
rect 58348 47194 58548 47200
rect 58348 47190 58360 47194
rect 58038 47180 58360 47190
rect 58038 47160 58170 47180
rect 57850 47154 58050 47160
rect 58160 47120 58170 47160
rect 58230 47160 58360 47180
rect 58536 47160 58548 47194
rect 58580 47190 58590 47250
rect 58650 47190 58660 47250
rect 58580 47170 58660 47190
rect 58230 47120 58240 47160
rect 58348 47154 58548 47160
rect 58160 47110 58240 47120
rect 57630 45950 57700 47100
rect 57630 45690 57650 45950
rect 57690 45690 57700 45950
rect 58710 47100 58720 47340
rect 58760 47100 58780 47340
rect 58710 45950 58780 47100
rect 58160 45920 58240 45930
rect 57850 45882 58050 45888
rect 57740 45850 57820 45870
rect 57740 45790 57750 45850
rect 57810 45838 57820 45850
rect 57850 45848 57862 45882
rect 58038 45880 58050 45882
rect 58160 45880 58170 45920
rect 58038 45860 58170 45880
rect 58230 45880 58240 45920
rect 58348 45882 58548 45888
rect 58348 45880 58360 45882
rect 58230 45860 58360 45880
rect 58038 45850 58360 45860
rect 58038 45848 58050 45850
rect 57850 45842 58050 45848
rect 58348 45848 58360 45850
rect 58536 45848 58548 45882
rect 58348 45842 58548 45848
rect 58580 45850 58660 45870
rect 57812 45804 57820 45838
rect 57810 45790 57820 45804
rect 57740 45770 57820 45790
rect 57850 45794 58050 45800
rect 57850 45760 57862 45794
rect 58038 45790 58050 45794
rect 58348 45794 58548 45800
rect 58348 45790 58360 45794
rect 58038 45760 58360 45790
rect 58536 45760 58548 45794
rect 58580 45790 58590 45850
rect 58650 45790 58660 45850
rect 58580 45770 58660 45790
rect 57850 45754 58050 45760
rect 57630 45630 57700 45690
rect 57630 45390 57650 45630
rect 57690 45390 57700 45630
rect 58160 45750 58240 45760
rect 58348 45754 58548 45760
rect 58160 45690 58170 45750
rect 58230 45690 58240 45750
rect 58160 45640 58240 45690
rect 58160 45580 58170 45640
rect 58230 45580 58240 45640
rect 57850 45572 58050 45578
rect 57740 45540 57820 45560
rect 57740 45480 57750 45540
rect 57810 45528 57820 45540
rect 57850 45538 57862 45572
rect 58038 45570 58050 45572
rect 58160 45570 58240 45580
rect 58710 45710 58720 45950
rect 58760 45710 58780 45950
rect 58710 45630 58780 45710
rect 58348 45572 58548 45578
rect 58348 45570 58360 45572
rect 58038 45540 58360 45570
rect 58038 45538 58050 45540
rect 57850 45532 58050 45538
rect 58348 45538 58360 45540
rect 58536 45538 58548 45572
rect 58348 45532 58548 45538
rect 58580 45540 58660 45560
rect 57812 45494 57820 45528
rect 57810 45480 57820 45494
rect 57740 45460 57820 45480
rect 57850 45484 58050 45490
rect 57850 45450 57862 45484
rect 58038 45480 58050 45484
rect 58348 45484 58548 45490
rect 58348 45480 58360 45484
rect 58038 45470 58360 45480
rect 58038 45450 58170 45470
rect 57850 45444 58050 45450
rect 58160 45410 58170 45450
rect 58230 45450 58360 45470
rect 58536 45450 58548 45484
rect 58580 45480 58590 45540
rect 58650 45480 58660 45540
rect 58580 45460 58660 45480
rect 58230 45410 58240 45450
rect 58348 45444 58548 45450
rect 58160 45400 58240 45410
rect 57630 44240 57700 45390
rect 57630 43980 57650 44240
rect 57690 43980 57700 44240
rect 58710 45390 58720 45630
rect 58760 45390 58780 45630
rect 58710 44240 58780 45390
rect 58160 44210 58240 44220
rect 57850 44172 58050 44178
rect 57740 44140 57820 44160
rect 57740 44080 57750 44140
rect 57810 44128 57820 44140
rect 57850 44138 57862 44172
rect 58038 44170 58050 44172
rect 58160 44170 58170 44210
rect 58038 44150 58170 44170
rect 58230 44170 58240 44210
rect 58348 44172 58548 44178
rect 58348 44170 58360 44172
rect 58230 44150 58360 44170
rect 58038 44140 58360 44150
rect 58038 44138 58050 44140
rect 57850 44132 58050 44138
rect 58348 44138 58360 44140
rect 58536 44138 58548 44172
rect 58348 44132 58548 44138
rect 58580 44140 58660 44160
rect 57812 44094 57820 44128
rect 57810 44080 57820 44094
rect 57740 44060 57820 44080
rect 57850 44084 58050 44090
rect 57850 44050 57862 44084
rect 58038 44080 58050 44084
rect 58348 44084 58548 44090
rect 58348 44080 58360 44084
rect 58038 44050 58360 44080
rect 58536 44050 58548 44084
rect 58580 44080 58590 44140
rect 58650 44080 58660 44140
rect 58580 44060 58660 44080
rect 57850 44044 58050 44050
rect 57630 43920 57700 43980
rect 57630 43680 57650 43920
rect 57690 43680 57700 43920
rect 58160 44040 58240 44050
rect 58348 44044 58548 44050
rect 58160 43980 58170 44040
rect 58230 43980 58240 44040
rect 58160 43930 58240 43980
rect 58160 43870 58170 43930
rect 58230 43870 58240 43930
rect 57850 43862 58050 43868
rect 57740 43830 57820 43850
rect 57740 43770 57750 43830
rect 57810 43818 57820 43830
rect 57850 43828 57862 43862
rect 58038 43860 58050 43862
rect 58160 43860 58240 43870
rect 58710 44000 58720 44240
rect 58760 44000 58780 44240
rect 58710 43920 58780 44000
rect 58348 43862 58548 43868
rect 58348 43860 58360 43862
rect 58038 43830 58360 43860
rect 58038 43828 58050 43830
rect 57850 43822 58050 43828
rect 58348 43828 58360 43830
rect 58536 43828 58548 43862
rect 58348 43822 58548 43828
rect 58580 43830 58660 43850
rect 57812 43784 57820 43818
rect 57810 43770 57820 43784
rect 57740 43750 57820 43770
rect 57850 43774 58050 43780
rect 57850 43740 57862 43774
rect 58038 43770 58050 43774
rect 58348 43774 58548 43780
rect 58348 43770 58360 43774
rect 58038 43760 58360 43770
rect 58038 43740 58170 43760
rect 57850 43734 58050 43740
rect 58160 43700 58170 43740
rect 58230 43740 58360 43760
rect 58536 43740 58548 43774
rect 58580 43770 58590 43830
rect 58650 43770 58660 43830
rect 58580 43750 58660 43770
rect 58230 43700 58240 43740
rect 58348 43734 58548 43740
rect 58160 43690 58240 43700
rect 57630 42530 57700 43680
rect 57630 42270 57650 42530
rect 57690 42270 57700 42530
rect 58710 43680 58720 43920
rect 58760 43680 58780 43920
rect 58710 42530 58780 43680
rect 58160 42500 58240 42510
rect 57850 42462 58050 42468
rect 57740 42430 57820 42450
rect 57740 42370 57750 42430
rect 57810 42418 57820 42430
rect 57850 42428 57862 42462
rect 58038 42460 58050 42462
rect 58160 42460 58170 42500
rect 58038 42440 58170 42460
rect 58230 42460 58240 42500
rect 58348 42462 58548 42468
rect 58348 42460 58360 42462
rect 58230 42440 58360 42460
rect 58038 42430 58360 42440
rect 58038 42428 58050 42430
rect 57850 42422 58050 42428
rect 58348 42428 58360 42430
rect 58536 42428 58548 42462
rect 58348 42422 58548 42428
rect 58580 42430 58660 42450
rect 57812 42384 57820 42418
rect 57810 42370 57820 42384
rect 57740 42350 57820 42370
rect 57850 42374 58050 42380
rect 57850 42340 57862 42374
rect 58038 42370 58050 42374
rect 58348 42374 58548 42380
rect 58348 42370 58360 42374
rect 58038 42340 58360 42370
rect 58536 42340 58548 42374
rect 58580 42370 58590 42430
rect 58650 42370 58660 42430
rect 58580 42350 58660 42370
rect 57850 42334 58050 42340
rect 57630 42210 57700 42270
rect 57630 41970 57650 42210
rect 57690 41970 57700 42210
rect 58160 42330 58240 42340
rect 58348 42334 58548 42340
rect 58160 42270 58170 42330
rect 58230 42270 58240 42330
rect 58160 42220 58240 42270
rect 58160 42160 58170 42220
rect 58230 42160 58240 42220
rect 57850 42152 58050 42158
rect 57740 42120 57820 42140
rect 57740 42060 57750 42120
rect 57810 42108 57820 42120
rect 57850 42118 57862 42152
rect 58038 42150 58050 42152
rect 58160 42150 58240 42160
rect 58710 42290 58720 42530
rect 58760 42290 58780 42530
rect 58710 42210 58780 42290
rect 58348 42152 58548 42158
rect 58348 42150 58360 42152
rect 58038 42120 58360 42150
rect 58038 42118 58050 42120
rect 57850 42112 58050 42118
rect 58348 42118 58360 42120
rect 58536 42118 58548 42152
rect 58348 42112 58548 42118
rect 58580 42120 58660 42140
rect 57812 42074 57820 42108
rect 57810 42060 57820 42074
rect 57740 42040 57820 42060
rect 57850 42064 58050 42070
rect 57850 42030 57862 42064
rect 58038 42060 58050 42064
rect 58348 42064 58548 42070
rect 58348 42060 58360 42064
rect 58038 42050 58360 42060
rect 58038 42030 58170 42050
rect 57850 42024 58050 42030
rect 58160 41990 58170 42030
rect 58230 42030 58360 42050
rect 58536 42030 58548 42064
rect 58580 42060 58590 42120
rect 58650 42060 58660 42120
rect 58580 42040 58660 42060
rect 58230 41990 58240 42030
rect 58348 42024 58548 42030
rect 58160 41980 58240 41990
rect 57630 40820 57700 41970
rect 57630 40560 57650 40820
rect 57690 40560 57700 40820
rect 58710 41970 58720 42210
rect 58760 41970 58780 42210
rect 58710 40820 58780 41970
rect 58160 40790 58240 40800
rect 57850 40752 58050 40758
rect 57740 40720 57820 40740
rect 57740 40660 57750 40720
rect 57810 40708 57820 40720
rect 57850 40718 57862 40752
rect 58038 40750 58050 40752
rect 58160 40750 58170 40790
rect 58038 40730 58170 40750
rect 58230 40750 58240 40790
rect 58348 40752 58548 40758
rect 58348 40750 58360 40752
rect 58230 40730 58360 40750
rect 58038 40720 58360 40730
rect 58038 40718 58050 40720
rect 57850 40712 58050 40718
rect 58348 40718 58360 40720
rect 58536 40718 58548 40752
rect 58348 40712 58548 40718
rect 58580 40720 58660 40740
rect 57812 40674 57820 40708
rect 57810 40660 57820 40674
rect 57740 40640 57820 40660
rect 57850 40664 58050 40670
rect 57850 40630 57862 40664
rect 58038 40660 58050 40664
rect 58348 40664 58548 40670
rect 58348 40660 58360 40664
rect 58038 40630 58360 40660
rect 58536 40630 58548 40664
rect 58580 40660 58590 40720
rect 58650 40660 58660 40720
rect 58580 40640 58660 40660
rect 57850 40624 58050 40630
rect 57630 40500 57700 40560
rect 57630 40260 57650 40500
rect 57690 40260 57700 40500
rect 58160 40620 58240 40630
rect 58348 40624 58548 40630
rect 58160 40560 58170 40620
rect 58230 40560 58240 40620
rect 58160 40510 58240 40560
rect 58160 40450 58170 40510
rect 58230 40450 58240 40510
rect 57850 40442 58050 40448
rect 57740 40410 57820 40430
rect 57740 40350 57750 40410
rect 57810 40398 57820 40410
rect 57850 40408 57862 40442
rect 58038 40440 58050 40442
rect 58160 40440 58240 40450
rect 58710 40580 58720 40820
rect 58760 40580 58780 40820
rect 58710 40500 58780 40580
rect 58348 40442 58548 40448
rect 58348 40440 58360 40442
rect 58038 40410 58360 40440
rect 58038 40408 58050 40410
rect 57850 40402 58050 40408
rect 58348 40408 58360 40410
rect 58536 40408 58548 40442
rect 58348 40402 58548 40408
rect 58580 40410 58660 40430
rect 57812 40364 57820 40398
rect 57810 40350 57820 40364
rect 57740 40330 57820 40350
rect 57850 40354 58050 40360
rect 57850 40320 57862 40354
rect 58038 40350 58050 40354
rect 58348 40354 58548 40360
rect 58348 40350 58360 40354
rect 58038 40340 58360 40350
rect 58038 40320 58170 40340
rect 57850 40314 58050 40320
rect 58160 40280 58170 40320
rect 58230 40320 58360 40340
rect 58536 40320 58548 40354
rect 58580 40350 58590 40410
rect 58650 40350 58660 40410
rect 58580 40330 58660 40350
rect 58230 40280 58240 40320
rect 58348 40314 58548 40320
rect 58160 40270 58240 40280
rect 57630 39690 57700 40260
rect 58710 40260 58720 40500
rect 58760 40260 58780 40500
rect 58710 39690 58780 40260
rect 57630 39680 57710 39690
rect 57630 39620 57640 39680
rect 57700 39620 57710 39680
rect 58700 39680 58780 39690
rect 58700 39620 58710 39680
rect 58770 39620 58780 39680
rect 58700 39610 58780 39620
rect 58810 66480 58840 67050
rect 58810 66470 58870 66480
rect 58810 66400 58870 66410
rect 58810 64770 58840 66400
rect 58900 65950 58930 67050
rect 58870 65940 58930 65950
rect 58870 65870 58930 65880
rect 58810 64760 58870 64770
rect 58810 64690 58870 64700
rect 58810 63060 58840 64690
rect 58900 64240 58930 65870
rect 58870 64230 58930 64240
rect 58870 64160 58930 64170
rect 58810 63050 58870 63060
rect 58810 62980 58870 62990
rect 58810 61350 58840 62980
rect 58900 62530 58930 64160
rect 58870 62520 58930 62530
rect 58870 62450 58930 62460
rect 58810 61340 58870 61350
rect 58810 61270 58870 61280
rect 58810 59640 58840 61270
rect 58900 60820 58930 62450
rect 58870 60810 58930 60820
rect 58870 60740 58930 60750
rect 58810 59630 58870 59640
rect 58810 59560 58870 59570
rect 58810 57930 58840 59560
rect 58900 59110 58930 60740
rect 58870 59100 58930 59110
rect 58870 59030 58930 59040
rect 58810 57920 58870 57930
rect 58810 57850 58870 57860
rect 58810 56220 58840 57850
rect 58900 57400 58930 59030
rect 58870 57390 58930 57400
rect 58870 57320 58930 57330
rect 58810 56210 58870 56220
rect 58810 56140 58870 56150
rect 58810 54510 58840 56140
rect 58900 55690 58930 57320
rect 58870 55680 58930 55690
rect 58870 55610 58930 55620
rect 58810 54500 58870 54510
rect 58810 54430 58870 54440
rect 58810 52800 58840 54430
rect 58900 53980 58930 55610
rect 58870 53970 58930 53980
rect 58870 53900 58930 53910
rect 58810 52790 58870 52800
rect 58810 52720 58870 52730
rect 58810 51090 58840 52720
rect 58900 52270 58930 53900
rect 58870 52260 58930 52270
rect 58870 52190 58930 52200
rect 58810 51080 58870 51090
rect 58810 51010 58870 51020
rect 58810 49380 58840 51010
rect 58900 50560 58930 52190
rect 58870 50550 58930 50560
rect 58870 50480 58930 50490
rect 58810 49370 58870 49380
rect 58810 49300 58870 49310
rect 58810 47670 58840 49300
rect 58900 48850 58930 50480
rect 58870 48840 58930 48850
rect 58870 48770 58930 48780
rect 58810 47660 58870 47670
rect 58810 47590 58870 47600
rect 58810 45960 58840 47590
rect 58900 47140 58930 48770
rect 58870 47130 58930 47140
rect 58870 47060 58930 47070
rect 58810 45950 58870 45960
rect 58810 45880 58870 45890
rect 58810 44250 58840 45880
rect 58900 45430 58930 47060
rect 58870 45420 58930 45430
rect 58870 45350 58930 45360
rect 58810 44240 58870 44250
rect 58810 44170 58870 44180
rect 58810 42540 58840 44170
rect 58900 43720 58930 45350
rect 58870 43710 58930 43720
rect 58870 43640 58930 43650
rect 58810 42530 58870 42540
rect 58810 42460 58870 42470
rect 58810 40830 58840 42460
rect 58900 42010 58930 43640
rect 58870 42000 58930 42010
rect 58870 41930 58930 41940
rect 58810 40820 58870 40830
rect 58810 40750 58870 40760
rect 57160 39220 57220 39230
rect 57340 39230 57600 39240
rect 54170 39160 54230 39170
rect 57400 39210 57600 39230
rect 57340 39160 57400 39170
rect 58810 38840 58840 40750
rect 58900 40300 58930 41930
rect 58870 40290 58930 40300
rect 58870 40220 58930 40230
rect 58900 39690 58930 40220
rect 58870 39680 58930 39690
rect 58870 39610 58930 39620
rect 58960 66390 58990 67050
rect 58960 66380 59020 66390
rect 58960 66310 59020 66320
rect 58960 64680 58990 66310
rect 58960 64670 59020 64680
rect 58960 64600 59020 64610
rect 58960 42450 58990 64600
rect 59080 62970 59110 67050
rect 59080 62960 59140 62970
rect 59080 62890 59140 62900
rect 59080 61250 59110 62890
rect 59080 61240 59140 61250
rect 59080 61170 59140 61180
rect 59080 45870 59110 61170
rect 59200 59550 59230 67050
rect 59200 59540 59260 59550
rect 59200 59470 59260 59480
rect 59200 47580 59230 59470
rect 59320 57840 59350 67050
rect 59320 57830 59380 57840
rect 59320 57760 59380 57770
rect 59320 56130 59350 57760
rect 59320 56120 59380 56130
rect 59320 56050 59380 56060
rect 59320 54420 59350 56050
rect 59320 54410 59380 54420
rect 59320 54340 59380 54350
rect 59320 52710 59350 54340
rect 59320 52700 59380 52710
rect 59320 52630 59380 52640
rect 59320 51000 59350 52630
rect 59320 50990 59380 51000
rect 59320 50920 59380 50930
rect 59320 49290 59350 50920
rect 59320 49280 59380 49290
rect 59320 49210 59380 49220
rect 59200 47570 59260 47580
rect 59200 47500 59260 47510
rect 59080 45860 59140 45870
rect 59080 45790 59140 45800
rect 59080 44160 59110 45790
rect 59080 44150 59140 44160
rect 59080 44080 59140 44090
rect 58960 42440 59020 42450
rect 58960 42370 59020 42380
rect 58960 40740 58990 42370
rect 58960 40730 59020 40740
rect 58960 40660 59020 40670
rect 58960 39240 58990 40660
rect 59080 39300 59110 44080
rect 59200 39360 59230 47500
rect 59320 39420 59350 49210
rect 59440 39690 59470 67050
rect 59560 39690 59590 67050
rect 59680 39690 59710 67050
rect 61840 39690 61870 67050
rect 61960 39690 61990 67050
rect 62080 39690 62110 67050
rect 62200 39690 62230 67050
rect 62320 39690 62350 67050
rect 62440 59550 62470 67050
rect 62560 66390 62590 67050
rect 62530 66380 62590 66390
rect 62530 66310 62590 66320
rect 62560 64680 62590 66310
rect 62530 64670 62590 64680
rect 62530 64600 62590 64610
rect 62560 62970 62590 64600
rect 62530 62960 62590 62970
rect 62530 62890 62590 62900
rect 62560 61260 62590 62890
rect 62530 61250 62590 61260
rect 62530 61180 62590 61190
rect 62410 59540 62470 59550
rect 62410 59470 62470 59480
rect 62440 57840 62470 59470
rect 62410 57830 62470 57840
rect 62410 57760 62470 57770
rect 62440 56130 62470 57760
rect 62410 56120 62470 56130
rect 62410 56050 62470 56060
rect 62440 54420 62470 56050
rect 62410 54410 62470 54420
rect 62410 54340 62470 54350
rect 62440 52710 62470 54340
rect 62410 52700 62470 52710
rect 62410 52630 62470 52640
rect 62440 51000 62470 52630
rect 62410 50990 62470 51000
rect 62410 50920 62470 50930
rect 62440 49290 62470 50920
rect 62410 49280 62470 49290
rect 62410 49210 62470 49220
rect 62440 47580 62470 49210
rect 62410 47570 62470 47580
rect 62410 47500 62470 47510
rect 59320 39410 59760 39420
rect 59320 39390 59700 39410
rect 59200 39350 59580 39360
rect 59200 39330 59520 39350
rect 59080 39290 59400 39300
rect 59080 39270 59340 39290
rect 58960 39230 59220 39240
rect 58960 39210 59160 39230
rect 59700 39340 59760 39350
rect 62440 39300 62470 47500
rect 62560 45870 62590 61180
rect 62530 45860 62590 45870
rect 62530 45790 62590 45800
rect 62560 44160 62590 45790
rect 62530 44150 62590 44160
rect 62530 44080 62590 44090
rect 62560 42450 62590 44080
rect 62530 42440 62590 42450
rect 62530 42370 62590 42380
rect 62560 40740 62590 42370
rect 62530 40730 62590 40740
rect 62530 40660 62590 40670
rect 59520 39280 59580 39290
rect 62150 39290 62470 39300
rect 59340 39220 59400 39230
rect 62210 39270 62470 39290
rect 62560 39240 62590 40660
rect 62620 66470 62690 67050
rect 62620 66210 62640 66470
rect 62680 66210 62690 66470
rect 63700 66470 63770 67050
rect 63150 66440 63230 66450
rect 62840 66402 63040 66408
rect 62730 66370 62810 66390
rect 62730 66310 62740 66370
rect 62800 66358 62810 66370
rect 62840 66368 62852 66402
rect 63028 66400 63040 66402
rect 63150 66400 63160 66440
rect 63028 66380 63160 66400
rect 63220 66400 63230 66440
rect 63338 66402 63538 66408
rect 63338 66400 63350 66402
rect 63220 66380 63350 66400
rect 63028 66370 63350 66380
rect 63028 66368 63040 66370
rect 62840 66362 63040 66368
rect 63338 66368 63350 66370
rect 63526 66368 63538 66402
rect 63338 66362 63538 66368
rect 63570 66370 63650 66390
rect 62802 66324 62810 66358
rect 62800 66310 62810 66324
rect 62730 66290 62810 66310
rect 62840 66314 63040 66320
rect 62840 66280 62852 66314
rect 63028 66310 63040 66314
rect 63338 66314 63538 66320
rect 63338 66310 63350 66314
rect 63028 66280 63350 66310
rect 63526 66280 63538 66314
rect 63570 66310 63580 66370
rect 63640 66310 63650 66370
rect 63570 66290 63650 66310
rect 62840 66274 63040 66280
rect 62620 66150 62690 66210
rect 62620 65910 62640 66150
rect 62680 65910 62690 66150
rect 63150 66270 63230 66280
rect 63338 66274 63538 66280
rect 63150 66210 63160 66270
rect 63220 66210 63230 66270
rect 63150 66160 63230 66210
rect 63150 66100 63160 66160
rect 63220 66100 63230 66160
rect 62840 66092 63040 66098
rect 62730 66060 62810 66080
rect 62730 66000 62740 66060
rect 62800 66048 62810 66060
rect 62840 66058 62852 66092
rect 63028 66090 63040 66092
rect 63150 66090 63230 66100
rect 63700 66230 63710 66470
rect 63750 66230 63770 66470
rect 63700 66150 63770 66230
rect 63338 66092 63538 66098
rect 63338 66090 63350 66092
rect 63028 66060 63350 66090
rect 63028 66058 63040 66060
rect 62840 66052 63040 66058
rect 63338 66058 63350 66060
rect 63526 66058 63538 66092
rect 63338 66052 63538 66058
rect 63570 66060 63650 66080
rect 62802 66014 62810 66048
rect 62800 66000 62810 66014
rect 62730 65980 62810 66000
rect 62840 66004 63040 66010
rect 62840 65970 62852 66004
rect 63028 66000 63040 66004
rect 63338 66004 63538 66010
rect 63338 66000 63350 66004
rect 63028 65990 63350 66000
rect 63028 65970 63160 65990
rect 62840 65964 63040 65970
rect 63150 65930 63160 65970
rect 63220 65970 63350 65990
rect 63526 65970 63538 66004
rect 63570 66000 63580 66060
rect 63640 66000 63650 66060
rect 63570 65980 63650 66000
rect 63220 65930 63230 65970
rect 63338 65964 63538 65970
rect 63150 65920 63230 65930
rect 62620 64760 62690 65910
rect 62620 64500 62640 64760
rect 62680 64500 62690 64760
rect 63700 65910 63710 66150
rect 63750 65910 63770 66150
rect 63700 64760 63770 65910
rect 63150 64730 63230 64740
rect 62840 64692 63040 64698
rect 62730 64660 62810 64680
rect 62730 64600 62740 64660
rect 62800 64648 62810 64660
rect 62840 64658 62852 64692
rect 63028 64690 63040 64692
rect 63150 64690 63160 64730
rect 63028 64670 63160 64690
rect 63220 64690 63230 64730
rect 63338 64692 63538 64698
rect 63338 64690 63350 64692
rect 63220 64670 63350 64690
rect 63028 64660 63350 64670
rect 63028 64658 63040 64660
rect 62840 64652 63040 64658
rect 63338 64658 63350 64660
rect 63526 64658 63538 64692
rect 63338 64652 63538 64658
rect 63570 64660 63650 64680
rect 62802 64614 62810 64648
rect 62800 64600 62810 64614
rect 62730 64580 62810 64600
rect 62840 64604 63040 64610
rect 62840 64570 62852 64604
rect 63028 64600 63040 64604
rect 63338 64604 63538 64610
rect 63338 64600 63350 64604
rect 63028 64570 63350 64600
rect 63526 64570 63538 64604
rect 63570 64600 63580 64660
rect 63640 64600 63650 64660
rect 63570 64580 63650 64600
rect 62840 64564 63040 64570
rect 62620 64440 62690 64500
rect 62620 64200 62640 64440
rect 62680 64200 62690 64440
rect 63150 64560 63230 64570
rect 63338 64564 63538 64570
rect 63150 64500 63160 64560
rect 63220 64500 63230 64560
rect 63150 64450 63230 64500
rect 63150 64390 63160 64450
rect 63220 64390 63230 64450
rect 62840 64382 63040 64388
rect 62730 64350 62810 64370
rect 62730 64290 62740 64350
rect 62800 64338 62810 64350
rect 62840 64348 62852 64382
rect 63028 64380 63040 64382
rect 63150 64380 63230 64390
rect 63700 64520 63710 64760
rect 63750 64520 63770 64760
rect 63700 64440 63770 64520
rect 63338 64382 63538 64388
rect 63338 64380 63350 64382
rect 63028 64350 63350 64380
rect 63028 64348 63040 64350
rect 62840 64342 63040 64348
rect 63338 64348 63350 64350
rect 63526 64348 63538 64382
rect 63338 64342 63538 64348
rect 63570 64350 63650 64370
rect 62802 64304 62810 64338
rect 62800 64290 62810 64304
rect 62730 64270 62810 64290
rect 62840 64294 63040 64300
rect 62840 64260 62852 64294
rect 63028 64290 63040 64294
rect 63338 64294 63538 64300
rect 63338 64290 63350 64294
rect 63028 64280 63350 64290
rect 63028 64260 63160 64280
rect 62840 64254 63040 64260
rect 63150 64220 63160 64260
rect 63220 64260 63350 64280
rect 63526 64260 63538 64294
rect 63570 64290 63580 64350
rect 63640 64290 63650 64350
rect 63570 64270 63650 64290
rect 63220 64220 63230 64260
rect 63338 64254 63538 64260
rect 63150 64210 63230 64220
rect 62620 63050 62690 64200
rect 62620 62790 62640 63050
rect 62680 62790 62690 63050
rect 63700 64200 63710 64440
rect 63750 64200 63770 64440
rect 63700 63050 63770 64200
rect 63150 63020 63230 63030
rect 62840 62982 63040 62988
rect 62730 62950 62810 62970
rect 62730 62890 62740 62950
rect 62800 62938 62810 62950
rect 62840 62948 62852 62982
rect 63028 62980 63040 62982
rect 63150 62980 63160 63020
rect 63028 62960 63160 62980
rect 63220 62980 63230 63020
rect 63338 62982 63538 62988
rect 63338 62980 63350 62982
rect 63220 62960 63350 62980
rect 63028 62950 63350 62960
rect 63028 62948 63040 62950
rect 62840 62942 63040 62948
rect 63338 62948 63350 62950
rect 63526 62948 63538 62982
rect 63338 62942 63538 62948
rect 63570 62950 63650 62970
rect 62802 62904 62810 62938
rect 62800 62890 62810 62904
rect 62730 62870 62810 62890
rect 62840 62894 63040 62900
rect 62840 62860 62852 62894
rect 63028 62890 63040 62894
rect 63338 62894 63538 62900
rect 63338 62890 63350 62894
rect 63028 62860 63350 62890
rect 63526 62860 63538 62894
rect 63570 62890 63580 62950
rect 63640 62890 63650 62950
rect 63570 62870 63650 62890
rect 62840 62854 63040 62860
rect 62620 62730 62690 62790
rect 62620 62490 62640 62730
rect 62680 62490 62690 62730
rect 63150 62850 63230 62860
rect 63338 62854 63538 62860
rect 63150 62790 63160 62850
rect 63220 62790 63230 62850
rect 63150 62740 63230 62790
rect 63150 62680 63160 62740
rect 63220 62680 63230 62740
rect 62840 62672 63040 62678
rect 62730 62640 62810 62660
rect 62730 62580 62740 62640
rect 62800 62628 62810 62640
rect 62840 62638 62852 62672
rect 63028 62670 63040 62672
rect 63150 62670 63230 62680
rect 63700 62810 63710 63050
rect 63750 62810 63770 63050
rect 63700 62730 63770 62810
rect 63338 62672 63538 62678
rect 63338 62670 63350 62672
rect 63028 62640 63350 62670
rect 63028 62638 63040 62640
rect 62840 62632 63040 62638
rect 63338 62638 63350 62640
rect 63526 62638 63538 62672
rect 63338 62632 63538 62638
rect 63570 62640 63650 62660
rect 62802 62594 62810 62628
rect 62800 62580 62810 62594
rect 62730 62560 62810 62580
rect 62840 62584 63040 62590
rect 62840 62550 62852 62584
rect 63028 62580 63040 62584
rect 63338 62584 63538 62590
rect 63338 62580 63350 62584
rect 63028 62570 63350 62580
rect 63028 62550 63160 62570
rect 62840 62544 63040 62550
rect 63150 62510 63160 62550
rect 63220 62550 63350 62570
rect 63526 62550 63538 62584
rect 63570 62580 63580 62640
rect 63640 62580 63650 62640
rect 63570 62560 63650 62580
rect 63220 62510 63230 62550
rect 63338 62544 63538 62550
rect 63150 62500 63230 62510
rect 62620 61340 62690 62490
rect 62620 61080 62640 61340
rect 62680 61080 62690 61340
rect 63700 62490 63710 62730
rect 63750 62490 63770 62730
rect 63700 61340 63770 62490
rect 63150 61310 63230 61320
rect 62840 61272 63040 61278
rect 62730 61240 62810 61260
rect 62730 61180 62740 61240
rect 62800 61228 62810 61240
rect 62840 61238 62852 61272
rect 63028 61270 63040 61272
rect 63150 61270 63160 61310
rect 63028 61250 63160 61270
rect 63220 61270 63230 61310
rect 63338 61272 63538 61278
rect 63338 61270 63350 61272
rect 63220 61250 63350 61270
rect 63028 61240 63350 61250
rect 63028 61238 63040 61240
rect 62840 61232 63040 61238
rect 63338 61238 63350 61240
rect 63526 61238 63538 61272
rect 63338 61232 63538 61238
rect 63570 61240 63650 61260
rect 62802 61194 62810 61228
rect 62800 61180 62810 61194
rect 62730 61160 62810 61180
rect 62840 61184 63040 61190
rect 62840 61150 62852 61184
rect 63028 61180 63040 61184
rect 63338 61184 63538 61190
rect 63338 61180 63350 61184
rect 63028 61150 63350 61180
rect 63526 61150 63538 61184
rect 63570 61180 63580 61240
rect 63640 61180 63650 61240
rect 63570 61160 63650 61180
rect 62840 61144 63040 61150
rect 62620 61020 62690 61080
rect 62620 60780 62640 61020
rect 62680 60780 62690 61020
rect 63150 61140 63230 61150
rect 63338 61144 63538 61150
rect 63150 61080 63160 61140
rect 63220 61080 63230 61140
rect 63150 61030 63230 61080
rect 63150 60970 63160 61030
rect 63220 60970 63230 61030
rect 62840 60962 63040 60968
rect 62730 60930 62810 60950
rect 62730 60870 62740 60930
rect 62800 60918 62810 60930
rect 62840 60928 62852 60962
rect 63028 60960 63040 60962
rect 63150 60960 63230 60970
rect 63700 61100 63710 61340
rect 63750 61100 63770 61340
rect 63700 61020 63770 61100
rect 63338 60962 63538 60968
rect 63338 60960 63350 60962
rect 63028 60930 63350 60960
rect 63028 60928 63040 60930
rect 62840 60922 63040 60928
rect 63338 60928 63350 60930
rect 63526 60928 63538 60962
rect 63338 60922 63538 60928
rect 63570 60930 63650 60950
rect 62802 60884 62810 60918
rect 62800 60870 62810 60884
rect 62730 60850 62810 60870
rect 62840 60874 63040 60880
rect 62840 60840 62852 60874
rect 63028 60870 63040 60874
rect 63338 60874 63538 60880
rect 63338 60870 63350 60874
rect 63028 60860 63350 60870
rect 63028 60840 63160 60860
rect 62840 60834 63040 60840
rect 63150 60800 63160 60840
rect 63220 60840 63350 60860
rect 63526 60840 63538 60874
rect 63570 60870 63580 60930
rect 63640 60870 63650 60930
rect 63570 60850 63650 60870
rect 63220 60800 63230 60840
rect 63338 60834 63538 60840
rect 63150 60790 63230 60800
rect 62620 59630 62690 60780
rect 62620 59370 62640 59630
rect 62680 59370 62690 59630
rect 63700 60780 63710 61020
rect 63750 60780 63770 61020
rect 63700 59630 63770 60780
rect 63150 59600 63230 59610
rect 62840 59562 63040 59568
rect 62730 59530 62810 59550
rect 62730 59470 62740 59530
rect 62800 59518 62810 59530
rect 62840 59528 62852 59562
rect 63028 59560 63040 59562
rect 63150 59560 63160 59600
rect 63028 59540 63160 59560
rect 63220 59560 63230 59600
rect 63338 59562 63538 59568
rect 63338 59560 63350 59562
rect 63220 59540 63350 59560
rect 63028 59530 63350 59540
rect 63028 59528 63040 59530
rect 62840 59522 63040 59528
rect 63338 59528 63350 59530
rect 63526 59528 63538 59562
rect 63338 59522 63538 59528
rect 63570 59530 63650 59550
rect 62802 59484 62810 59518
rect 62800 59470 62810 59484
rect 62730 59450 62810 59470
rect 62840 59474 63040 59480
rect 62840 59440 62852 59474
rect 63028 59470 63040 59474
rect 63338 59474 63538 59480
rect 63338 59470 63350 59474
rect 63028 59440 63350 59470
rect 63526 59440 63538 59474
rect 63570 59470 63580 59530
rect 63640 59470 63650 59530
rect 63570 59450 63650 59470
rect 62840 59434 63040 59440
rect 62620 59310 62690 59370
rect 62620 59070 62640 59310
rect 62680 59070 62690 59310
rect 63150 59430 63230 59440
rect 63338 59434 63538 59440
rect 63150 59370 63160 59430
rect 63220 59370 63230 59430
rect 63150 59320 63230 59370
rect 63150 59260 63160 59320
rect 63220 59260 63230 59320
rect 62840 59252 63040 59258
rect 62730 59220 62810 59240
rect 62730 59160 62740 59220
rect 62800 59208 62810 59220
rect 62840 59218 62852 59252
rect 63028 59250 63040 59252
rect 63150 59250 63230 59260
rect 63700 59390 63710 59630
rect 63750 59390 63770 59630
rect 63700 59310 63770 59390
rect 63338 59252 63538 59258
rect 63338 59250 63350 59252
rect 63028 59220 63350 59250
rect 63028 59218 63040 59220
rect 62840 59212 63040 59218
rect 63338 59218 63350 59220
rect 63526 59218 63538 59252
rect 63338 59212 63538 59218
rect 63570 59220 63650 59240
rect 62802 59174 62810 59208
rect 62800 59160 62810 59174
rect 62730 59140 62810 59160
rect 62840 59164 63040 59170
rect 62840 59130 62852 59164
rect 63028 59160 63040 59164
rect 63338 59164 63538 59170
rect 63338 59160 63350 59164
rect 63028 59150 63350 59160
rect 63028 59130 63160 59150
rect 62840 59124 63040 59130
rect 63150 59090 63160 59130
rect 63220 59130 63350 59150
rect 63526 59130 63538 59164
rect 63570 59160 63580 59220
rect 63640 59160 63650 59220
rect 63570 59140 63650 59160
rect 63220 59090 63230 59130
rect 63338 59124 63538 59130
rect 63150 59080 63230 59090
rect 62620 57920 62690 59070
rect 62620 57660 62640 57920
rect 62680 57660 62690 57920
rect 63700 59070 63710 59310
rect 63750 59070 63770 59310
rect 63700 57920 63770 59070
rect 63150 57890 63230 57900
rect 62840 57852 63040 57858
rect 62730 57820 62810 57840
rect 62730 57760 62740 57820
rect 62800 57808 62810 57820
rect 62840 57818 62852 57852
rect 63028 57850 63040 57852
rect 63150 57850 63160 57890
rect 63028 57830 63160 57850
rect 63220 57850 63230 57890
rect 63338 57852 63538 57858
rect 63338 57850 63350 57852
rect 63220 57830 63350 57850
rect 63028 57820 63350 57830
rect 63028 57818 63040 57820
rect 62840 57812 63040 57818
rect 63338 57818 63350 57820
rect 63526 57818 63538 57852
rect 63338 57812 63538 57818
rect 63570 57820 63650 57840
rect 62802 57774 62810 57808
rect 62800 57760 62810 57774
rect 62730 57740 62810 57760
rect 62840 57764 63040 57770
rect 62840 57730 62852 57764
rect 63028 57760 63040 57764
rect 63338 57764 63538 57770
rect 63338 57760 63350 57764
rect 63028 57730 63350 57760
rect 63526 57730 63538 57764
rect 63570 57760 63580 57820
rect 63640 57760 63650 57820
rect 63570 57740 63650 57760
rect 62840 57724 63040 57730
rect 62620 57600 62690 57660
rect 62620 57360 62640 57600
rect 62680 57360 62690 57600
rect 63150 57720 63230 57730
rect 63338 57724 63538 57730
rect 63150 57660 63160 57720
rect 63220 57660 63230 57720
rect 63150 57610 63230 57660
rect 63150 57550 63160 57610
rect 63220 57550 63230 57610
rect 62840 57542 63040 57548
rect 62730 57510 62810 57530
rect 62730 57450 62740 57510
rect 62800 57498 62810 57510
rect 62840 57508 62852 57542
rect 63028 57540 63040 57542
rect 63150 57540 63230 57550
rect 63700 57680 63710 57920
rect 63750 57680 63770 57920
rect 63700 57600 63770 57680
rect 63338 57542 63538 57548
rect 63338 57540 63350 57542
rect 63028 57510 63350 57540
rect 63028 57508 63040 57510
rect 62840 57502 63040 57508
rect 63338 57508 63350 57510
rect 63526 57508 63538 57542
rect 63338 57502 63538 57508
rect 63570 57510 63650 57530
rect 62802 57464 62810 57498
rect 62800 57450 62810 57464
rect 62730 57430 62810 57450
rect 62840 57454 63040 57460
rect 62840 57420 62852 57454
rect 63028 57450 63040 57454
rect 63338 57454 63538 57460
rect 63338 57450 63350 57454
rect 63028 57440 63350 57450
rect 63028 57420 63160 57440
rect 62840 57414 63040 57420
rect 63150 57380 63160 57420
rect 63220 57420 63350 57440
rect 63526 57420 63538 57454
rect 63570 57450 63580 57510
rect 63640 57450 63650 57510
rect 63570 57430 63650 57450
rect 63220 57380 63230 57420
rect 63338 57414 63538 57420
rect 63150 57370 63230 57380
rect 62620 56210 62690 57360
rect 62620 55950 62640 56210
rect 62680 55950 62690 56210
rect 63700 57360 63710 57600
rect 63750 57360 63770 57600
rect 63700 56210 63770 57360
rect 63150 56180 63230 56190
rect 62840 56142 63040 56148
rect 62730 56110 62810 56130
rect 62730 56050 62740 56110
rect 62800 56098 62810 56110
rect 62840 56108 62852 56142
rect 63028 56140 63040 56142
rect 63150 56140 63160 56180
rect 63028 56120 63160 56140
rect 63220 56140 63230 56180
rect 63338 56142 63538 56148
rect 63338 56140 63350 56142
rect 63220 56120 63350 56140
rect 63028 56110 63350 56120
rect 63028 56108 63040 56110
rect 62840 56102 63040 56108
rect 63338 56108 63350 56110
rect 63526 56108 63538 56142
rect 63338 56102 63538 56108
rect 63570 56110 63650 56130
rect 62802 56064 62810 56098
rect 62800 56050 62810 56064
rect 62730 56030 62810 56050
rect 62840 56054 63040 56060
rect 62840 56020 62852 56054
rect 63028 56050 63040 56054
rect 63338 56054 63538 56060
rect 63338 56050 63350 56054
rect 63028 56020 63350 56050
rect 63526 56020 63538 56054
rect 63570 56050 63580 56110
rect 63640 56050 63650 56110
rect 63570 56030 63650 56050
rect 62840 56014 63040 56020
rect 62620 55890 62690 55950
rect 62620 55650 62640 55890
rect 62680 55650 62690 55890
rect 63150 56010 63230 56020
rect 63338 56014 63538 56020
rect 63150 55950 63160 56010
rect 63220 55950 63230 56010
rect 63150 55900 63230 55950
rect 63150 55840 63160 55900
rect 63220 55840 63230 55900
rect 62840 55832 63040 55838
rect 62730 55800 62810 55820
rect 62730 55740 62740 55800
rect 62800 55788 62810 55800
rect 62840 55798 62852 55832
rect 63028 55830 63040 55832
rect 63150 55830 63230 55840
rect 63700 55970 63710 56210
rect 63750 55970 63770 56210
rect 63700 55890 63770 55970
rect 63338 55832 63538 55838
rect 63338 55830 63350 55832
rect 63028 55800 63350 55830
rect 63028 55798 63040 55800
rect 62840 55792 63040 55798
rect 63338 55798 63350 55800
rect 63526 55798 63538 55832
rect 63338 55792 63538 55798
rect 63570 55800 63650 55820
rect 62802 55754 62810 55788
rect 62800 55740 62810 55754
rect 62730 55720 62810 55740
rect 62840 55744 63040 55750
rect 62840 55710 62852 55744
rect 63028 55740 63040 55744
rect 63338 55744 63538 55750
rect 63338 55740 63350 55744
rect 63028 55730 63350 55740
rect 63028 55710 63160 55730
rect 62840 55704 63040 55710
rect 63150 55670 63160 55710
rect 63220 55710 63350 55730
rect 63526 55710 63538 55744
rect 63570 55740 63580 55800
rect 63640 55740 63650 55800
rect 63570 55720 63650 55740
rect 63220 55670 63230 55710
rect 63338 55704 63538 55710
rect 63150 55660 63230 55670
rect 62620 54500 62690 55650
rect 62620 54240 62640 54500
rect 62680 54240 62690 54500
rect 63700 55650 63710 55890
rect 63750 55650 63770 55890
rect 63700 54500 63770 55650
rect 63150 54470 63230 54480
rect 62840 54432 63040 54438
rect 62730 54400 62810 54420
rect 62730 54340 62740 54400
rect 62800 54388 62810 54400
rect 62840 54398 62852 54432
rect 63028 54430 63040 54432
rect 63150 54430 63160 54470
rect 63028 54410 63160 54430
rect 63220 54430 63230 54470
rect 63338 54432 63538 54438
rect 63338 54430 63350 54432
rect 63220 54410 63350 54430
rect 63028 54400 63350 54410
rect 63028 54398 63040 54400
rect 62840 54392 63040 54398
rect 63338 54398 63350 54400
rect 63526 54398 63538 54432
rect 63338 54392 63538 54398
rect 63570 54400 63650 54420
rect 62802 54354 62810 54388
rect 62800 54340 62810 54354
rect 62730 54320 62810 54340
rect 62840 54344 63040 54350
rect 62840 54310 62852 54344
rect 63028 54340 63040 54344
rect 63338 54344 63538 54350
rect 63338 54340 63350 54344
rect 63028 54310 63350 54340
rect 63526 54310 63538 54344
rect 63570 54340 63580 54400
rect 63640 54340 63650 54400
rect 63570 54320 63650 54340
rect 62840 54304 63040 54310
rect 62620 54180 62690 54240
rect 62620 53940 62640 54180
rect 62680 53940 62690 54180
rect 63150 54300 63230 54310
rect 63338 54304 63538 54310
rect 63150 54240 63160 54300
rect 63220 54240 63230 54300
rect 63150 54190 63230 54240
rect 63150 54130 63160 54190
rect 63220 54130 63230 54190
rect 62840 54122 63040 54128
rect 62730 54090 62810 54110
rect 62730 54030 62740 54090
rect 62800 54078 62810 54090
rect 62840 54088 62852 54122
rect 63028 54120 63040 54122
rect 63150 54120 63230 54130
rect 63700 54260 63710 54500
rect 63750 54260 63770 54500
rect 63700 54180 63770 54260
rect 63338 54122 63538 54128
rect 63338 54120 63350 54122
rect 63028 54090 63350 54120
rect 63028 54088 63040 54090
rect 62840 54082 63040 54088
rect 63338 54088 63350 54090
rect 63526 54088 63538 54122
rect 63338 54082 63538 54088
rect 63570 54090 63650 54110
rect 62802 54044 62810 54078
rect 62800 54030 62810 54044
rect 62730 54010 62810 54030
rect 62840 54034 63040 54040
rect 62840 54000 62852 54034
rect 63028 54030 63040 54034
rect 63338 54034 63538 54040
rect 63338 54030 63350 54034
rect 63028 54020 63350 54030
rect 63028 54000 63160 54020
rect 62840 53994 63040 54000
rect 63150 53960 63160 54000
rect 63220 54000 63350 54020
rect 63526 54000 63538 54034
rect 63570 54030 63580 54090
rect 63640 54030 63650 54090
rect 63570 54010 63650 54030
rect 63220 53960 63230 54000
rect 63338 53994 63538 54000
rect 63150 53950 63230 53960
rect 62620 52790 62690 53940
rect 62620 52530 62640 52790
rect 62680 52530 62690 52790
rect 63700 53940 63710 54180
rect 63750 53940 63770 54180
rect 63700 52790 63770 53940
rect 63150 52760 63230 52770
rect 62840 52722 63040 52728
rect 62730 52690 62810 52710
rect 62730 52630 62740 52690
rect 62800 52678 62810 52690
rect 62840 52688 62852 52722
rect 63028 52720 63040 52722
rect 63150 52720 63160 52760
rect 63028 52700 63160 52720
rect 63220 52720 63230 52760
rect 63338 52722 63538 52728
rect 63338 52720 63350 52722
rect 63220 52700 63350 52720
rect 63028 52690 63350 52700
rect 63028 52688 63040 52690
rect 62840 52682 63040 52688
rect 63338 52688 63350 52690
rect 63526 52688 63538 52722
rect 63338 52682 63538 52688
rect 63570 52690 63650 52710
rect 62802 52644 62810 52678
rect 62800 52630 62810 52644
rect 62730 52610 62810 52630
rect 62840 52634 63040 52640
rect 62840 52600 62852 52634
rect 63028 52630 63040 52634
rect 63338 52634 63538 52640
rect 63338 52630 63350 52634
rect 63028 52600 63350 52630
rect 63526 52600 63538 52634
rect 63570 52630 63580 52690
rect 63640 52630 63650 52690
rect 63570 52610 63650 52630
rect 62840 52594 63040 52600
rect 62620 52470 62690 52530
rect 62620 52230 62640 52470
rect 62680 52230 62690 52470
rect 63150 52590 63230 52600
rect 63338 52594 63538 52600
rect 63150 52530 63160 52590
rect 63220 52530 63230 52590
rect 63150 52480 63230 52530
rect 63150 52420 63160 52480
rect 63220 52420 63230 52480
rect 62840 52412 63040 52418
rect 62730 52380 62810 52400
rect 62730 52320 62740 52380
rect 62800 52368 62810 52380
rect 62840 52378 62852 52412
rect 63028 52410 63040 52412
rect 63150 52410 63230 52420
rect 63700 52550 63710 52790
rect 63750 52550 63770 52790
rect 63700 52470 63770 52550
rect 63338 52412 63538 52418
rect 63338 52410 63350 52412
rect 63028 52380 63350 52410
rect 63028 52378 63040 52380
rect 62840 52372 63040 52378
rect 63338 52378 63350 52380
rect 63526 52378 63538 52412
rect 63338 52372 63538 52378
rect 63570 52380 63650 52400
rect 62802 52334 62810 52368
rect 62800 52320 62810 52334
rect 62730 52300 62810 52320
rect 62840 52324 63040 52330
rect 62840 52290 62852 52324
rect 63028 52320 63040 52324
rect 63338 52324 63538 52330
rect 63338 52320 63350 52324
rect 63028 52310 63350 52320
rect 63028 52290 63160 52310
rect 62840 52284 63040 52290
rect 63150 52250 63160 52290
rect 63220 52290 63350 52310
rect 63526 52290 63538 52324
rect 63570 52320 63580 52380
rect 63640 52320 63650 52380
rect 63570 52300 63650 52320
rect 63220 52250 63230 52290
rect 63338 52284 63538 52290
rect 63150 52240 63230 52250
rect 62620 51080 62690 52230
rect 62620 50820 62640 51080
rect 62680 50820 62690 51080
rect 63700 52230 63710 52470
rect 63750 52230 63770 52470
rect 63700 51080 63770 52230
rect 63150 51050 63230 51060
rect 62840 51012 63040 51018
rect 62730 50980 62810 51000
rect 62730 50920 62740 50980
rect 62800 50968 62810 50980
rect 62840 50978 62852 51012
rect 63028 51010 63040 51012
rect 63150 51010 63160 51050
rect 63028 50990 63160 51010
rect 63220 51010 63230 51050
rect 63338 51012 63538 51018
rect 63338 51010 63350 51012
rect 63220 50990 63350 51010
rect 63028 50980 63350 50990
rect 63028 50978 63040 50980
rect 62840 50972 63040 50978
rect 63338 50978 63350 50980
rect 63526 50978 63538 51012
rect 63338 50972 63538 50978
rect 63570 50980 63650 51000
rect 62802 50934 62810 50968
rect 62800 50920 62810 50934
rect 62730 50900 62810 50920
rect 62840 50924 63040 50930
rect 62840 50890 62852 50924
rect 63028 50920 63040 50924
rect 63338 50924 63538 50930
rect 63338 50920 63350 50924
rect 63028 50890 63350 50920
rect 63526 50890 63538 50924
rect 63570 50920 63580 50980
rect 63640 50920 63650 50980
rect 63570 50900 63650 50920
rect 62840 50884 63040 50890
rect 62620 50760 62690 50820
rect 62620 50520 62640 50760
rect 62680 50520 62690 50760
rect 63150 50880 63230 50890
rect 63338 50884 63538 50890
rect 63150 50820 63160 50880
rect 63220 50820 63230 50880
rect 63150 50770 63230 50820
rect 63150 50710 63160 50770
rect 63220 50710 63230 50770
rect 62840 50702 63040 50708
rect 62730 50670 62810 50690
rect 62730 50610 62740 50670
rect 62800 50658 62810 50670
rect 62840 50668 62852 50702
rect 63028 50700 63040 50702
rect 63150 50700 63230 50710
rect 63700 50840 63710 51080
rect 63750 50840 63770 51080
rect 63700 50760 63770 50840
rect 63338 50702 63538 50708
rect 63338 50700 63350 50702
rect 63028 50670 63350 50700
rect 63028 50668 63040 50670
rect 62840 50662 63040 50668
rect 63338 50668 63350 50670
rect 63526 50668 63538 50702
rect 63338 50662 63538 50668
rect 63570 50670 63650 50690
rect 62802 50624 62810 50658
rect 62800 50610 62810 50624
rect 62730 50590 62810 50610
rect 62840 50614 63040 50620
rect 62840 50580 62852 50614
rect 63028 50610 63040 50614
rect 63338 50614 63538 50620
rect 63338 50610 63350 50614
rect 63028 50600 63350 50610
rect 63028 50580 63160 50600
rect 62840 50574 63040 50580
rect 63150 50540 63160 50580
rect 63220 50580 63350 50600
rect 63526 50580 63538 50614
rect 63570 50610 63580 50670
rect 63640 50610 63650 50670
rect 63570 50590 63650 50610
rect 63220 50540 63230 50580
rect 63338 50574 63538 50580
rect 63150 50530 63230 50540
rect 62620 49370 62690 50520
rect 62620 49110 62640 49370
rect 62680 49110 62690 49370
rect 63700 50520 63710 50760
rect 63750 50520 63770 50760
rect 63700 49370 63770 50520
rect 63150 49340 63230 49350
rect 62840 49302 63040 49308
rect 62730 49270 62810 49290
rect 62730 49210 62740 49270
rect 62800 49258 62810 49270
rect 62840 49268 62852 49302
rect 63028 49300 63040 49302
rect 63150 49300 63160 49340
rect 63028 49280 63160 49300
rect 63220 49300 63230 49340
rect 63338 49302 63538 49308
rect 63338 49300 63350 49302
rect 63220 49280 63350 49300
rect 63028 49270 63350 49280
rect 63028 49268 63040 49270
rect 62840 49262 63040 49268
rect 63338 49268 63350 49270
rect 63526 49268 63538 49302
rect 63338 49262 63538 49268
rect 63570 49270 63650 49290
rect 62802 49224 62810 49258
rect 62800 49210 62810 49224
rect 62730 49190 62810 49210
rect 62840 49214 63040 49220
rect 62840 49180 62852 49214
rect 63028 49210 63040 49214
rect 63338 49214 63538 49220
rect 63338 49210 63350 49214
rect 63028 49180 63350 49210
rect 63526 49180 63538 49214
rect 63570 49210 63580 49270
rect 63640 49210 63650 49270
rect 63570 49190 63650 49210
rect 62840 49174 63040 49180
rect 62620 49050 62690 49110
rect 62620 48810 62640 49050
rect 62680 48810 62690 49050
rect 63150 49170 63230 49180
rect 63338 49174 63538 49180
rect 63150 49110 63160 49170
rect 63220 49110 63230 49170
rect 63150 49060 63230 49110
rect 63150 49000 63160 49060
rect 63220 49000 63230 49060
rect 62840 48992 63040 48998
rect 62730 48960 62810 48980
rect 62730 48900 62740 48960
rect 62800 48948 62810 48960
rect 62840 48958 62852 48992
rect 63028 48990 63040 48992
rect 63150 48990 63230 49000
rect 63700 49130 63710 49370
rect 63750 49130 63770 49370
rect 63700 49050 63770 49130
rect 63338 48992 63538 48998
rect 63338 48990 63350 48992
rect 63028 48960 63350 48990
rect 63028 48958 63040 48960
rect 62840 48952 63040 48958
rect 63338 48958 63350 48960
rect 63526 48958 63538 48992
rect 63338 48952 63538 48958
rect 63570 48960 63650 48980
rect 62802 48914 62810 48948
rect 62800 48900 62810 48914
rect 62730 48880 62810 48900
rect 62840 48904 63040 48910
rect 62840 48870 62852 48904
rect 63028 48900 63040 48904
rect 63338 48904 63538 48910
rect 63338 48900 63350 48904
rect 63028 48890 63350 48900
rect 63028 48870 63160 48890
rect 62840 48864 63040 48870
rect 63150 48830 63160 48870
rect 63220 48870 63350 48890
rect 63526 48870 63538 48904
rect 63570 48900 63580 48960
rect 63640 48900 63650 48960
rect 63570 48880 63650 48900
rect 63220 48830 63230 48870
rect 63338 48864 63538 48870
rect 63150 48820 63230 48830
rect 62620 47660 62690 48810
rect 62620 47400 62640 47660
rect 62680 47400 62690 47660
rect 63700 48810 63710 49050
rect 63750 48810 63770 49050
rect 63700 47660 63770 48810
rect 63150 47630 63230 47640
rect 62840 47592 63040 47598
rect 62730 47560 62810 47580
rect 62730 47500 62740 47560
rect 62800 47548 62810 47560
rect 62840 47558 62852 47592
rect 63028 47590 63040 47592
rect 63150 47590 63160 47630
rect 63028 47570 63160 47590
rect 63220 47590 63230 47630
rect 63338 47592 63538 47598
rect 63338 47590 63350 47592
rect 63220 47570 63350 47590
rect 63028 47560 63350 47570
rect 63028 47558 63040 47560
rect 62840 47552 63040 47558
rect 63338 47558 63350 47560
rect 63526 47558 63538 47592
rect 63338 47552 63538 47558
rect 63570 47560 63650 47580
rect 62802 47514 62810 47548
rect 62800 47500 62810 47514
rect 62730 47480 62810 47500
rect 62840 47504 63040 47510
rect 62840 47470 62852 47504
rect 63028 47500 63040 47504
rect 63338 47504 63538 47510
rect 63338 47500 63350 47504
rect 63028 47470 63350 47500
rect 63526 47470 63538 47504
rect 63570 47500 63580 47560
rect 63640 47500 63650 47560
rect 63570 47480 63650 47500
rect 62840 47464 63040 47470
rect 62620 47340 62690 47400
rect 62620 47100 62640 47340
rect 62680 47100 62690 47340
rect 63150 47460 63230 47470
rect 63338 47464 63538 47470
rect 63150 47400 63160 47460
rect 63220 47400 63230 47460
rect 63150 47350 63230 47400
rect 63150 47290 63160 47350
rect 63220 47290 63230 47350
rect 62840 47282 63040 47288
rect 62730 47250 62810 47270
rect 62730 47190 62740 47250
rect 62800 47238 62810 47250
rect 62840 47248 62852 47282
rect 63028 47280 63040 47282
rect 63150 47280 63230 47290
rect 63700 47420 63710 47660
rect 63750 47420 63770 47660
rect 63700 47340 63770 47420
rect 63338 47282 63538 47288
rect 63338 47280 63350 47282
rect 63028 47250 63350 47280
rect 63028 47248 63040 47250
rect 62840 47242 63040 47248
rect 63338 47248 63350 47250
rect 63526 47248 63538 47282
rect 63338 47242 63538 47248
rect 63570 47250 63650 47270
rect 62802 47204 62810 47238
rect 62800 47190 62810 47204
rect 62730 47170 62810 47190
rect 62840 47194 63040 47200
rect 62840 47160 62852 47194
rect 63028 47190 63040 47194
rect 63338 47194 63538 47200
rect 63338 47190 63350 47194
rect 63028 47180 63350 47190
rect 63028 47160 63160 47180
rect 62840 47154 63040 47160
rect 63150 47120 63160 47160
rect 63220 47160 63350 47180
rect 63526 47160 63538 47194
rect 63570 47190 63580 47250
rect 63640 47190 63650 47250
rect 63570 47170 63650 47190
rect 63220 47120 63230 47160
rect 63338 47154 63538 47160
rect 63150 47110 63230 47120
rect 62620 45950 62690 47100
rect 62620 45690 62640 45950
rect 62680 45690 62690 45950
rect 63700 47100 63710 47340
rect 63750 47100 63770 47340
rect 63700 45950 63770 47100
rect 63150 45920 63230 45930
rect 62840 45882 63040 45888
rect 62730 45850 62810 45870
rect 62730 45790 62740 45850
rect 62800 45838 62810 45850
rect 62840 45848 62852 45882
rect 63028 45880 63040 45882
rect 63150 45880 63160 45920
rect 63028 45860 63160 45880
rect 63220 45880 63230 45920
rect 63338 45882 63538 45888
rect 63338 45880 63350 45882
rect 63220 45860 63350 45880
rect 63028 45850 63350 45860
rect 63028 45848 63040 45850
rect 62840 45842 63040 45848
rect 63338 45848 63350 45850
rect 63526 45848 63538 45882
rect 63338 45842 63538 45848
rect 63570 45850 63650 45870
rect 62802 45804 62810 45838
rect 62800 45790 62810 45804
rect 62730 45770 62810 45790
rect 62840 45794 63040 45800
rect 62840 45760 62852 45794
rect 63028 45790 63040 45794
rect 63338 45794 63538 45800
rect 63338 45790 63350 45794
rect 63028 45760 63350 45790
rect 63526 45760 63538 45794
rect 63570 45790 63580 45850
rect 63640 45790 63650 45850
rect 63570 45770 63650 45790
rect 62840 45754 63040 45760
rect 62620 45630 62690 45690
rect 62620 45390 62640 45630
rect 62680 45390 62690 45630
rect 63150 45750 63230 45760
rect 63338 45754 63538 45760
rect 63150 45690 63160 45750
rect 63220 45690 63230 45750
rect 63150 45640 63230 45690
rect 63150 45580 63160 45640
rect 63220 45580 63230 45640
rect 62840 45572 63040 45578
rect 62730 45540 62810 45560
rect 62730 45480 62740 45540
rect 62800 45528 62810 45540
rect 62840 45538 62852 45572
rect 63028 45570 63040 45572
rect 63150 45570 63230 45580
rect 63700 45710 63710 45950
rect 63750 45710 63770 45950
rect 63700 45630 63770 45710
rect 63338 45572 63538 45578
rect 63338 45570 63350 45572
rect 63028 45540 63350 45570
rect 63028 45538 63040 45540
rect 62840 45532 63040 45538
rect 63338 45538 63350 45540
rect 63526 45538 63538 45572
rect 63338 45532 63538 45538
rect 63570 45540 63650 45560
rect 62802 45494 62810 45528
rect 62800 45480 62810 45494
rect 62730 45460 62810 45480
rect 62840 45484 63040 45490
rect 62840 45450 62852 45484
rect 63028 45480 63040 45484
rect 63338 45484 63538 45490
rect 63338 45480 63350 45484
rect 63028 45470 63350 45480
rect 63028 45450 63160 45470
rect 62840 45444 63040 45450
rect 63150 45410 63160 45450
rect 63220 45450 63350 45470
rect 63526 45450 63538 45484
rect 63570 45480 63580 45540
rect 63640 45480 63650 45540
rect 63570 45460 63650 45480
rect 63220 45410 63230 45450
rect 63338 45444 63538 45450
rect 63150 45400 63230 45410
rect 62620 44240 62690 45390
rect 62620 43980 62640 44240
rect 62680 43980 62690 44240
rect 63700 45390 63710 45630
rect 63750 45390 63770 45630
rect 63700 44240 63770 45390
rect 63150 44210 63230 44220
rect 62840 44172 63040 44178
rect 62730 44140 62810 44160
rect 62730 44080 62740 44140
rect 62800 44128 62810 44140
rect 62840 44138 62852 44172
rect 63028 44170 63040 44172
rect 63150 44170 63160 44210
rect 63028 44150 63160 44170
rect 63220 44170 63230 44210
rect 63338 44172 63538 44178
rect 63338 44170 63350 44172
rect 63220 44150 63350 44170
rect 63028 44140 63350 44150
rect 63028 44138 63040 44140
rect 62840 44132 63040 44138
rect 63338 44138 63350 44140
rect 63526 44138 63538 44172
rect 63338 44132 63538 44138
rect 63570 44140 63650 44160
rect 62802 44094 62810 44128
rect 62800 44080 62810 44094
rect 62730 44060 62810 44080
rect 62840 44084 63040 44090
rect 62840 44050 62852 44084
rect 63028 44080 63040 44084
rect 63338 44084 63538 44090
rect 63338 44080 63350 44084
rect 63028 44050 63350 44080
rect 63526 44050 63538 44084
rect 63570 44080 63580 44140
rect 63640 44080 63650 44140
rect 63570 44060 63650 44080
rect 62840 44044 63040 44050
rect 62620 43920 62690 43980
rect 62620 43680 62640 43920
rect 62680 43680 62690 43920
rect 63150 44040 63230 44050
rect 63338 44044 63538 44050
rect 63150 43980 63160 44040
rect 63220 43980 63230 44040
rect 63150 43930 63230 43980
rect 63150 43870 63160 43930
rect 63220 43870 63230 43930
rect 62840 43862 63040 43868
rect 62730 43830 62810 43850
rect 62730 43770 62740 43830
rect 62800 43818 62810 43830
rect 62840 43828 62852 43862
rect 63028 43860 63040 43862
rect 63150 43860 63230 43870
rect 63700 44000 63710 44240
rect 63750 44000 63770 44240
rect 63700 43920 63770 44000
rect 63338 43862 63538 43868
rect 63338 43860 63350 43862
rect 63028 43830 63350 43860
rect 63028 43828 63040 43830
rect 62840 43822 63040 43828
rect 63338 43828 63350 43830
rect 63526 43828 63538 43862
rect 63338 43822 63538 43828
rect 63570 43830 63650 43850
rect 62802 43784 62810 43818
rect 62800 43770 62810 43784
rect 62730 43750 62810 43770
rect 62840 43774 63040 43780
rect 62840 43740 62852 43774
rect 63028 43770 63040 43774
rect 63338 43774 63538 43780
rect 63338 43770 63350 43774
rect 63028 43760 63350 43770
rect 63028 43740 63160 43760
rect 62840 43734 63040 43740
rect 63150 43700 63160 43740
rect 63220 43740 63350 43760
rect 63526 43740 63538 43774
rect 63570 43770 63580 43830
rect 63640 43770 63650 43830
rect 63570 43750 63650 43770
rect 63220 43700 63230 43740
rect 63338 43734 63538 43740
rect 63150 43690 63230 43700
rect 62620 42530 62690 43680
rect 62620 42270 62640 42530
rect 62680 42270 62690 42530
rect 63700 43680 63710 43920
rect 63750 43680 63770 43920
rect 63700 42530 63770 43680
rect 63150 42500 63230 42510
rect 62840 42462 63040 42468
rect 62730 42430 62810 42450
rect 62730 42370 62740 42430
rect 62800 42418 62810 42430
rect 62840 42428 62852 42462
rect 63028 42460 63040 42462
rect 63150 42460 63160 42500
rect 63028 42440 63160 42460
rect 63220 42460 63230 42500
rect 63338 42462 63538 42468
rect 63338 42460 63350 42462
rect 63220 42440 63350 42460
rect 63028 42430 63350 42440
rect 63028 42428 63040 42430
rect 62840 42422 63040 42428
rect 63338 42428 63350 42430
rect 63526 42428 63538 42462
rect 63338 42422 63538 42428
rect 63570 42430 63650 42450
rect 62802 42384 62810 42418
rect 62800 42370 62810 42384
rect 62730 42350 62810 42370
rect 62840 42374 63040 42380
rect 62840 42340 62852 42374
rect 63028 42370 63040 42374
rect 63338 42374 63538 42380
rect 63338 42370 63350 42374
rect 63028 42340 63350 42370
rect 63526 42340 63538 42374
rect 63570 42370 63580 42430
rect 63640 42370 63650 42430
rect 63570 42350 63650 42370
rect 62840 42334 63040 42340
rect 62620 42210 62690 42270
rect 62620 41970 62640 42210
rect 62680 41970 62690 42210
rect 63150 42330 63230 42340
rect 63338 42334 63538 42340
rect 63150 42270 63160 42330
rect 63220 42270 63230 42330
rect 63150 42220 63230 42270
rect 63150 42160 63160 42220
rect 63220 42160 63230 42220
rect 62840 42152 63040 42158
rect 62730 42120 62810 42140
rect 62730 42060 62740 42120
rect 62800 42108 62810 42120
rect 62840 42118 62852 42152
rect 63028 42150 63040 42152
rect 63150 42150 63230 42160
rect 63700 42290 63710 42530
rect 63750 42290 63770 42530
rect 63700 42210 63770 42290
rect 63338 42152 63538 42158
rect 63338 42150 63350 42152
rect 63028 42120 63350 42150
rect 63028 42118 63040 42120
rect 62840 42112 63040 42118
rect 63338 42118 63350 42120
rect 63526 42118 63538 42152
rect 63338 42112 63538 42118
rect 63570 42120 63650 42140
rect 62802 42074 62810 42108
rect 62800 42060 62810 42074
rect 62730 42040 62810 42060
rect 62840 42064 63040 42070
rect 62840 42030 62852 42064
rect 63028 42060 63040 42064
rect 63338 42064 63538 42070
rect 63338 42060 63350 42064
rect 63028 42050 63350 42060
rect 63028 42030 63160 42050
rect 62840 42024 63040 42030
rect 63150 41990 63160 42030
rect 63220 42030 63350 42050
rect 63526 42030 63538 42064
rect 63570 42060 63580 42120
rect 63640 42060 63650 42120
rect 63570 42040 63650 42060
rect 63220 41990 63230 42030
rect 63338 42024 63538 42030
rect 63150 41980 63230 41990
rect 62620 40820 62690 41970
rect 62620 40560 62640 40820
rect 62680 40560 62690 40820
rect 63700 41970 63710 42210
rect 63750 41970 63770 42210
rect 63700 40820 63770 41970
rect 63150 40790 63230 40800
rect 62840 40752 63040 40758
rect 62730 40720 62810 40740
rect 62730 40660 62740 40720
rect 62800 40708 62810 40720
rect 62840 40718 62852 40752
rect 63028 40750 63040 40752
rect 63150 40750 63160 40790
rect 63028 40730 63160 40750
rect 63220 40750 63230 40790
rect 63338 40752 63538 40758
rect 63338 40750 63350 40752
rect 63220 40730 63350 40750
rect 63028 40720 63350 40730
rect 63028 40718 63040 40720
rect 62840 40712 63040 40718
rect 63338 40718 63350 40720
rect 63526 40718 63538 40752
rect 63338 40712 63538 40718
rect 63570 40720 63650 40740
rect 62802 40674 62810 40708
rect 62800 40660 62810 40674
rect 62730 40640 62810 40660
rect 62840 40664 63040 40670
rect 62840 40630 62852 40664
rect 63028 40660 63040 40664
rect 63338 40664 63538 40670
rect 63338 40660 63350 40664
rect 63028 40630 63350 40660
rect 63526 40630 63538 40664
rect 63570 40660 63580 40720
rect 63640 40660 63650 40720
rect 63570 40640 63650 40660
rect 62840 40624 63040 40630
rect 62620 40500 62690 40560
rect 62620 40260 62640 40500
rect 62680 40260 62690 40500
rect 63150 40620 63230 40630
rect 63338 40624 63538 40630
rect 63150 40560 63160 40620
rect 63220 40560 63230 40620
rect 63150 40510 63230 40560
rect 63150 40450 63160 40510
rect 63220 40450 63230 40510
rect 62840 40442 63040 40448
rect 62730 40410 62810 40430
rect 62730 40350 62740 40410
rect 62800 40398 62810 40410
rect 62840 40408 62852 40442
rect 63028 40440 63040 40442
rect 63150 40440 63230 40450
rect 63700 40580 63710 40820
rect 63750 40580 63770 40820
rect 63700 40500 63770 40580
rect 63338 40442 63538 40448
rect 63338 40440 63350 40442
rect 63028 40410 63350 40440
rect 63028 40408 63040 40410
rect 62840 40402 63040 40408
rect 63338 40408 63350 40410
rect 63526 40408 63538 40442
rect 63338 40402 63538 40408
rect 63570 40410 63650 40430
rect 62802 40364 62810 40398
rect 62800 40350 62810 40364
rect 62730 40330 62810 40350
rect 62840 40354 63040 40360
rect 62840 40320 62852 40354
rect 63028 40350 63040 40354
rect 63338 40354 63538 40360
rect 63338 40350 63350 40354
rect 63028 40340 63350 40350
rect 63028 40320 63160 40340
rect 62840 40314 63040 40320
rect 63150 40280 63160 40320
rect 63220 40320 63350 40340
rect 63526 40320 63538 40354
rect 63570 40350 63580 40410
rect 63640 40350 63650 40410
rect 63570 40330 63650 40350
rect 63220 40280 63230 40320
rect 63338 40314 63538 40320
rect 63150 40270 63230 40280
rect 62620 39690 62690 40260
rect 63700 40260 63710 40500
rect 63750 40260 63770 40500
rect 63700 39690 63770 40260
rect 62620 39680 62700 39690
rect 62620 39620 62630 39680
rect 62690 39620 62700 39680
rect 63690 39680 63770 39690
rect 63690 39620 63700 39680
rect 63760 39620 63770 39680
rect 63690 39610 63770 39620
rect 63800 66480 63830 67050
rect 63800 66470 63860 66480
rect 63800 66400 63860 66410
rect 63800 64770 63830 66400
rect 63890 65950 63920 67050
rect 63860 65940 63920 65950
rect 63860 65870 63920 65880
rect 63800 64760 63860 64770
rect 63800 64690 63860 64700
rect 63800 63060 63830 64690
rect 63890 64240 63920 65870
rect 63860 64230 63920 64240
rect 63860 64160 63920 64170
rect 63800 63050 63860 63060
rect 63800 62980 63860 62990
rect 63800 61350 63830 62980
rect 63890 62530 63920 64160
rect 63860 62520 63920 62530
rect 63860 62450 63920 62460
rect 63800 61340 63860 61350
rect 63800 61270 63860 61280
rect 63800 59640 63830 61270
rect 63890 60820 63920 62450
rect 63860 60810 63920 60820
rect 63860 60740 63920 60750
rect 63800 59630 63860 59640
rect 63800 59560 63860 59570
rect 63800 57930 63830 59560
rect 63890 59110 63920 60740
rect 63860 59100 63920 59110
rect 63860 59030 63920 59040
rect 63800 57920 63860 57930
rect 63800 57850 63860 57860
rect 63800 56220 63830 57850
rect 63890 57400 63920 59030
rect 63860 57390 63920 57400
rect 63860 57320 63920 57330
rect 63800 56210 63860 56220
rect 63800 56140 63860 56150
rect 63800 54510 63830 56140
rect 63890 55690 63920 57320
rect 63860 55680 63920 55690
rect 63860 55610 63920 55620
rect 63800 54500 63860 54510
rect 63800 54430 63860 54440
rect 63800 52800 63830 54430
rect 63890 53980 63920 55610
rect 63860 53970 63920 53980
rect 63860 53900 63920 53910
rect 63800 52790 63860 52800
rect 63800 52720 63860 52730
rect 63800 51090 63830 52720
rect 63890 52270 63920 53900
rect 63860 52260 63920 52270
rect 63860 52190 63920 52200
rect 63800 51080 63860 51090
rect 63800 51010 63860 51020
rect 63800 49380 63830 51010
rect 63890 50560 63920 52190
rect 63860 50550 63920 50560
rect 63860 50480 63920 50490
rect 63800 49370 63860 49380
rect 63800 49300 63860 49310
rect 63800 47670 63830 49300
rect 63890 48850 63920 50480
rect 63860 48840 63920 48850
rect 63860 48770 63920 48780
rect 63800 47660 63860 47670
rect 63800 47590 63860 47600
rect 63800 45960 63830 47590
rect 63890 47140 63920 48770
rect 63860 47130 63920 47140
rect 63860 47060 63920 47070
rect 63800 45950 63860 45960
rect 63800 45880 63860 45890
rect 63800 44250 63830 45880
rect 63890 45430 63920 47060
rect 63860 45420 63920 45430
rect 63860 45350 63920 45360
rect 63800 44240 63860 44250
rect 63800 44170 63860 44180
rect 63800 42540 63830 44170
rect 63890 43720 63920 45350
rect 63860 43710 63920 43720
rect 63860 43640 63920 43650
rect 63800 42530 63860 42540
rect 63800 42460 63860 42470
rect 63800 40830 63830 42460
rect 63890 42010 63920 43640
rect 63860 42000 63920 42010
rect 63860 41930 63920 41940
rect 63800 40820 63860 40830
rect 63800 40750 63860 40760
rect 62150 39220 62210 39230
rect 62330 39230 62590 39240
rect 59160 39160 59220 39170
rect 62390 39210 62590 39230
rect 62330 39160 62390 39170
rect 63800 38840 63830 40750
rect 63890 40300 63920 41930
rect 63860 40290 63920 40300
rect 63860 40220 63920 40230
rect 63890 39690 63920 40220
rect 63860 39680 63920 39690
rect 63860 39610 63920 39620
rect 63950 66390 63980 67050
rect 63950 66380 64010 66390
rect 63950 66310 64010 66320
rect 63950 64680 63980 66310
rect 63950 64670 64010 64680
rect 63950 64600 64010 64610
rect 63950 62970 63980 64600
rect 63950 62960 64010 62970
rect 63950 62890 64010 62900
rect 63950 61260 63980 62890
rect 63950 61250 64010 61260
rect 63950 61180 64010 61190
rect 63950 45870 63980 61180
rect 64070 59550 64100 67050
rect 64070 59540 64130 59550
rect 64070 59470 64130 59480
rect 64070 57840 64100 59470
rect 64070 57830 64130 57840
rect 64070 57760 64130 57770
rect 64070 56130 64100 57760
rect 64070 56120 64130 56130
rect 64070 56050 64130 56060
rect 64070 54420 64100 56050
rect 64070 54410 64130 54420
rect 64070 54340 64130 54350
rect 64070 52710 64100 54340
rect 64070 52700 64130 52710
rect 64070 52630 64130 52640
rect 64070 51000 64100 52630
rect 64070 50990 64130 51000
rect 64070 50920 64130 50930
rect 64070 49290 64100 50920
rect 64070 49280 64130 49290
rect 64070 49210 64130 49220
rect 64070 47580 64100 49210
rect 64070 47570 64130 47580
rect 64070 47500 64130 47510
rect 63950 45860 64010 45870
rect 63950 45790 64010 45800
rect 63950 44160 63980 45790
rect 63950 44150 64010 44160
rect 63950 44080 64010 44090
rect 63950 42450 63980 44080
rect 63950 42440 64010 42450
rect 63950 42370 64010 42380
rect 63950 40740 63980 42370
rect 63950 40730 64010 40740
rect 63950 40660 64010 40670
rect 63950 39240 63980 40660
rect 64070 39300 64100 47500
rect 64190 39690 64220 67050
rect 64310 39690 64340 67050
rect 64430 39690 64460 67050
rect 64550 39690 64580 67050
rect 64670 39690 64700 67050
rect 66830 39690 66860 67050
rect 66950 39690 66980 67050
rect 67070 39690 67100 67050
rect 67190 39690 67220 67050
rect 67310 39690 67340 67050
rect 67430 59550 67460 67050
rect 67550 66390 67580 67050
rect 67520 66380 67580 66390
rect 67520 66310 67580 66320
rect 67550 64680 67580 66310
rect 67520 64670 67580 64680
rect 67520 64600 67580 64610
rect 67550 62970 67580 64600
rect 67520 62960 67580 62970
rect 67520 62890 67580 62900
rect 67550 61260 67580 62890
rect 67520 61250 67580 61260
rect 67520 61180 67580 61190
rect 67400 59540 67460 59550
rect 67400 59470 67460 59480
rect 67430 57840 67460 59470
rect 67400 57830 67460 57840
rect 67400 57760 67460 57770
rect 67430 56130 67460 57760
rect 67400 56120 67460 56130
rect 67400 56050 67460 56060
rect 67430 54420 67460 56050
rect 67400 54410 67460 54420
rect 67400 54340 67460 54350
rect 67430 52710 67460 54340
rect 67400 52700 67460 52710
rect 67400 52630 67460 52640
rect 67430 51000 67460 52630
rect 67400 50990 67460 51000
rect 67400 50920 67460 50930
rect 67430 49290 67460 50920
rect 67400 49280 67460 49290
rect 67400 49210 67460 49220
rect 67430 47580 67460 49210
rect 67400 47570 67460 47580
rect 67400 47500 67460 47510
rect 67430 39300 67460 47500
rect 67550 45870 67580 61180
rect 67520 45860 67580 45870
rect 67520 45790 67580 45800
rect 67550 44160 67580 45790
rect 67520 44150 67580 44160
rect 67520 44080 67580 44090
rect 67550 42450 67580 44080
rect 67520 42440 67580 42450
rect 67520 42370 67580 42380
rect 67550 40740 67580 42370
rect 67520 40730 67580 40740
rect 67520 40660 67580 40670
rect 64070 39290 64390 39300
rect 64070 39270 64330 39290
rect 63950 39230 64210 39240
rect 63950 39210 64150 39230
rect 64330 39220 64390 39230
rect 67140 39290 67460 39300
rect 67200 39270 67460 39290
rect 67550 39240 67580 40660
rect 67610 66470 67680 67050
rect 67610 66210 67630 66470
rect 67670 66210 67680 66470
rect 68690 66470 68760 67050
rect 68140 66440 68220 66450
rect 67830 66402 68030 66408
rect 67720 66370 67800 66390
rect 67720 66310 67730 66370
rect 67790 66358 67800 66370
rect 67830 66368 67842 66402
rect 68018 66400 68030 66402
rect 68140 66400 68150 66440
rect 68018 66380 68150 66400
rect 68210 66400 68220 66440
rect 68328 66402 68528 66408
rect 68328 66400 68340 66402
rect 68210 66380 68340 66400
rect 68018 66370 68340 66380
rect 68018 66368 68030 66370
rect 67830 66362 68030 66368
rect 68328 66368 68340 66370
rect 68516 66368 68528 66402
rect 68328 66362 68528 66368
rect 68560 66370 68640 66390
rect 67792 66324 67800 66358
rect 67790 66310 67800 66324
rect 67720 66290 67800 66310
rect 67830 66314 68030 66320
rect 67830 66280 67842 66314
rect 68018 66310 68030 66314
rect 68328 66314 68528 66320
rect 68328 66310 68340 66314
rect 68018 66280 68340 66310
rect 68516 66280 68528 66314
rect 68560 66310 68570 66370
rect 68630 66310 68640 66370
rect 68560 66290 68640 66310
rect 67830 66274 68030 66280
rect 67610 66150 67680 66210
rect 67610 65910 67630 66150
rect 67670 65910 67680 66150
rect 68140 66270 68220 66280
rect 68328 66274 68528 66280
rect 68140 66210 68150 66270
rect 68210 66210 68220 66270
rect 68140 66160 68220 66210
rect 68140 66100 68150 66160
rect 68210 66100 68220 66160
rect 67830 66092 68030 66098
rect 67720 66060 67800 66080
rect 67720 66000 67730 66060
rect 67790 66048 67800 66060
rect 67830 66058 67842 66092
rect 68018 66090 68030 66092
rect 68140 66090 68220 66100
rect 68690 66230 68700 66470
rect 68740 66230 68760 66470
rect 68690 66150 68760 66230
rect 68328 66092 68528 66098
rect 68328 66090 68340 66092
rect 68018 66060 68340 66090
rect 68018 66058 68030 66060
rect 67830 66052 68030 66058
rect 68328 66058 68340 66060
rect 68516 66058 68528 66092
rect 68328 66052 68528 66058
rect 68560 66060 68640 66080
rect 67792 66014 67800 66048
rect 67790 66000 67800 66014
rect 67720 65980 67800 66000
rect 67830 66004 68030 66010
rect 67830 65970 67842 66004
rect 68018 66000 68030 66004
rect 68328 66004 68528 66010
rect 68328 66000 68340 66004
rect 68018 65990 68340 66000
rect 68018 65970 68150 65990
rect 67830 65964 68030 65970
rect 68140 65930 68150 65970
rect 68210 65970 68340 65990
rect 68516 65970 68528 66004
rect 68560 66000 68570 66060
rect 68630 66000 68640 66060
rect 68560 65980 68640 66000
rect 68210 65930 68220 65970
rect 68328 65964 68528 65970
rect 68140 65920 68220 65930
rect 67610 64760 67680 65910
rect 67610 64500 67630 64760
rect 67670 64500 67680 64760
rect 68690 65910 68700 66150
rect 68740 65910 68760 66150
rect 68690 64760 68760 65910
rect 68140 64730 68220 64740
rect 67830 64692 68030 64698
rect 67720 64660 67800 64680
rect 67720 64600 67730 64660
rect 67790 64648 67800 64660
rect 67830 64658 67842 64692
rect 68018 64690 68030 64692
rect 68140 64690 68150 64730
rect 68018 64670 68150 64690
rect 68210 64690 68220 64730
rect 68328 64692 68528 64698
rect 68328 64690 68340 64692
rect 68210 64670 68340 64690
rect 68018 64660 68340 64670
rect 68018 64658 68030 64660
rect 67830 64652 68030 64658
rect 68328 64658 68340 64660
rect 68516 64658 68528 64692
rect 68328 64652 68528 64658
rect 68560 64660 68640 64680
rect 67792 64614 67800 64648
rect 67790 64600 67800 64614
rect 67720 64580 67800 64600
rect 67830 64604 68030 64610
rect 67830 64570 67842 64604
rect 68018 64600 68030 64604
rect 68328 64604 68528 64610
rect 68328 64600 68340 64604
rect 68018 64570 68340 64600
rect 68516 64570 68528 64604
rect 68560 64600 68570 64660
rect 68630 64600 68640 64660
rect 68560 64580 68640 64600
rect 67830 64564 68030 64570
rect 67610 64440 67680 64500
rect 67610 64200 67630 64440
rect 67670 64200 67680 64440
rect 68140 64560 68220 64570
rect 68328 64564 68528 64570
rect 68140 64500 68150 64560
rect 68210 64500 68220 64560
rect 68140 64450 68220 64500
rect 68140 64390 68150 64450
rect 68210 64390 68220 64450
rect 67830 64382 68030 64388
rect 67720 64350 67800 64370
rect 67720 64290 67730 64350
rect 67790 64338 67800 64350
rect 67830 64348 67842 64382
rect 68018 64380 68030 64382
rect 68140 64380 68220 64390
rect 68690 64520 68700 64760
rect 68740 64520 68760 64760
rect 68690 64440 68760 64520
rect 68328 64382 68528 64388
rect 68328 64380 68340 64382
rect 68018 64350 68340 64380
rect 68018 64348 68030 64350
rect 67830 64342 68030 64348
rect 68328 64348 68340 64350
rect 68516 64348 68528 64382
rect 68328 64342 68528 64348
rect 68560 64350 68640 64370
rect 67792 64304 67800 64338
rect 67790 64290 67800 64304
rect 67720 64270 67800 64290
rect 67830 64294 68030 64300
rect 67830 64260 67842 64294
rect 68018 64290 68030 64294
rect 68328 64294 68528 64300
rect 68328 64290 68340 64294
rect 68018 64280 68340 64290
rect 68018 64260 68150 64280
rect 67830 64254 68030 64260
rect 68140 64220 68150 64260
rect 68210 64260 68340 64280
rect 68516 64260 68528 64294
rect 68560 64290 68570 64350
rect 68630 64290 68640 64350
rect 68560 64270 68640 64290
rect 68210 64220 68220 64260
rect 68328 64254 68528 64260
rect 68140 64210 68220 64220
rect 67610 63050 67680 64200
rect 67610 62790 67630 63050
rect 67670 62790 67680 63050
rect 68690 64200 68700 64440
rect 68740 64200 68760 64440
rect 68690 63050 68760 64200
rect 68140 63020 68220 63030
rect 67830 62982 68030 62988
rect 67720 62950 67800 62970
rect 67720 62890 67730 62950
rect 67790 62938 67800 62950
rect 67830 62948 67842 62982
rect 68018 62980 68030 62982
rect 68140 62980 68150 63020
rect 68018 62960 68150 62980
rect 68210 62980 68220 63020
rect 68328 62982 68528 62988
rect 68328 62980 68340 62982
rect 68210 62960 68340 62980
rect 68018 62950 68340 62960
rect 68018 62948 68030 62950
rect 67830 62942 68030 62948
rect 68328 62948 68340 62950
rect 68516 62948 68528 62982
rect 68328 62942 68528 62948
rect 68560 62950 68640 62970
rect 67792 62904 67800 62938
rect 67790 62890 67800 62904
rect 67720 62870 67800 62890
rect 67830 62894 68030 62900
rect 67830 62860 67842 62894
rect 68018 62890 68030 62894
rect 68328 62894 68528 62900
rect 68328 62890 68340 62894
rect 68018 62860 68340 62890
rect 68516 62860 68528 62894
rect 68560 62890 68570 62950
rect 68630 62890 68640 62950
rect 68560 62870 68640 62890
rect 67830 62854 68030 62860
rect 67610 62730 67680 62790
rect 67610 62490 67630 62730
rect 67670 62490 67680 62730
rect 68140 62850 68220 62860
rect 68328 62854 68528 62860
rect 68140 62790 68150 62850
rect 68210 62790 68220 62850
rect 68140 62740 68220 62790
rect 68140 62680 68150 62740
rect 68210 62680 68220 62740
rect 67830 62672 68030 62678
rect 67720 62640 67800 62660
rect 67720 62580 67730 62640
rect 67790 62628 67800 62640
rect 67830 62638 67842 62672
rect 68018 62670 68030 62672
rect 68140 62670 68220 62680
rect 68690 62810 68700 63050
rect 68740 62810 68760 63050
rect 68690 62730 68760 62810
rect 68328 62672 68528 62678
rect 68328 62670 68340 62672
rect 68018 62640 68340 62670
rect 68018 62638 68030 62640
rect 67830 62632 68030 62638
rect 68328 62638 68340 62640
rect 68516 62638 68528 62672
rect 68328 62632 68528 62638
rect 68560 62640 68640 62660
rect 67792 62594 67800 62628
rect 67790 62580 67800 62594
rect 67720 62560 67800 62580
rect 67830 62584 68030 62590
rect 67830 62550 67842 62584
rect 68018 62580 68030 62584
rect 68328 62584 68528 62590
rect 68328 62580 68340 62584
rect 68018 62570 68340 62580
rect 68018 62550 68150 62570
rect 67830 62544 68030 62550
rect 68140 62510 68150 62550
rect 68210 62550 68340 62570
rect 68516 62550 68528 62584
rect 68560 62580 68570 62640
rect 68630 62580 68640 62640
rect 68560 62560 68640 62580
rect 68210 62510 68220 62550
rect 68328 62544 68528 62550
rect 68140 62500 68220 62510
rect 67610 61340 67680 62490
rect 67610 61080 67630 61340
rect 67670 61080 67680 61340
rect 68690 62490 68700 62730
rect 68740 62490 68760 62730
rect 68690 61340 68760 62490
rect 68140 61310 68220 61320
rect 67830 61272 68030 61278
rect 67720 61240 67800 61260
rect 67720 61180 67730 61240
rect 67790 61228 67800 61240
rect 67830 61238 67842 61272
rect 68018 61270 68030 61272
rect 68140 61270 68150 61310
rect 68018 61250 68150 61270
rect 68210 61270 68220 61310
rect 68328 61272 68528 61278
rect 68328 61270 68340 61272
rect 68210 61250 68340 61270
rect 68018 61240 68340 61250
rect 68018 61238 68030 61240
rect 67830 61232 68030 61238
rect 68328 61238 68340 61240
rect 68516 61238 68528 61272
rect 68328 61232 68528 61238
rect 68560 61240 68640 61260
rect 67792 61194 67800 61228
rect 67790 61180 67800 61194
rect 67720 61160 67800 61180
rect 67830 61184 68030 61190
rect 67830 61150 67842 61184
rect 68018 61180 68030 61184
rect 68328 61184 68528 61190
rect 68328 61180 68340 61184
rect 68018 61150 68340 61180
rect 68516 61150 68528 61184
rect 68560 61180 68570 61240
rect 68630 61180 68640 61240
rect 68560 61160 68640 61180
rect 67830 61144 68030 61150
rect 67610 61020 67680 61080
rect 67610 60780 67630 61020
rect 67670 60780 67680 61020
rect 68140 61140 68220 61150
rect 68328 61144 68528 61150
rect 68140 61080 68150 61140
rect 68210 61080 68220 61140
rect 68140 61030 68220 61080
rect 68140 60970 68150 61030
rect 68210 60970 68220 61030
rect 67830 60962 68030 60968
rect 67720 60930 67800 60950
rect 67720 60870 67730 60930
rect 67790 60918 67800 60930
rect 67830 60928 67842 60962
rect 68018 60960 68030 60962
rect 68140 60960 68220 60970
rect 68690 61100 68700 61340
rect 68740 61100 68760 61340
rect 68690 61020 68760 61100
rect 68328 60962 68528 60968
rect 68328 60960 68340 60962
rect 68018 60930 68340 60960
rect 68018 60928 68030 60930
rect 67830 60922 68030 60928
rect 68328 60928 68340 60930
rect 68516 60928 68528 60962
rect 68328 60922 68528 60928
rect 68560 60930 68640 60950
rect 67792 60884 67800 60918
rect 67790 60870 67800 60884
rect 67720 60850 67800 60870
rect 67830 60874 68030 60880
rect 67830 60840 67842 60874
rect 68018 60870 68030 60874
rect 68328 60874 68528 60880
rect 68328 60870 68340 60874
rect 68018 60860 68340 60870
rect 68018 60840 68150 60860
rect 67830 60834 68030 60840
rect 68140 60800 68150 60840
rect 68210 60840 68340 60860
rect 68516 60840 68528 60874
rect 68560 60870 68570 60930
rect 68630 60870 68640 60930
rect 68560 60850 68640 60870
rect 68210 60800 68220 60840
rect 68328 60834 68528 60840
rect 68140 60790 68220 60800
rect 67610 59630 67680 60780
rect 67610 59370 67630 59630
rect 67670 59370 67680 59630
rect 68690 60780 68700 61020
rect 68740 60780 68760 61020
rect 68690 59630 68760 60780
rect 68140 59600 68220 59610
rect 67830 59562 68030 59568
rect 67720 59530 67800 59550
rect 67720 59470 67730 59530
rect 67790 59518 67800 59530
rect 67830 59528 67842 59562
rect 68018 59560 68030 59562
rect 68140 59560 68150 59600
rect 68018 59540 68150 59560
rect 68210 59560 68220 59600
rect 68328 59562 68528 59568
rect 68328 59560 68340 59562
rect 68210 59540 68340 59560
rect 68018 59530 68340 59540
rect 68018 59528 68030 59530
rect 67830 59522 68030 59528
rect 68328 59528 68340 59530
rect 68516 59528 68528 59562
rect 68328 59522 68528 59528
rect 68560 59530 68640 59550
rect 67792 59484 67800 59518
rect 67790 59470 67800 59484
rect 67720 59450 67800 59470
rect 67830 59474 68030 59480
rect 67830 59440 67842 59474
rect 68018 59470 68030 59474
rect 68328 59474 68528 59480
rect 68328 59470 68340 59474
rect 68018 59440 68340 59470
rect 68516 59440 68528 59474
rect 68560 59470 68570 59530
rect 68630 59470 68640 59530
rect 68560 59450 68640 59470
rect 67830 59434 68030 59440
rect 67610 59310 67680 59370
rect 67610 59070 67630 59310
rect 67670 59070 67680 59310
rect 68140 59430 68220 59440
rect 68328 59434 68528 59440
rect 68140 59370 68150 59430
rect 68210 59370 68220 59430
rect 68140 59320 68220 59370
rect 68140 59260 68150 59320
rect 68210 59260 68220 59320
rect 67830 59252 68030 59258
rect 67720 59220 67800 59240
rect 67720 59160 67730 59220
rect 67790 59208 67800 59220
rect 67830 59218 67842 59252
rect 68018 59250 68030 59252
rect 68140 59250 68220 59260
rect 68690 59390 68700 59630
rect 68740 59390 68760 59630
rect 68690 59310 68760 59390
rect 68328 59252 68528 59258
rect 68328 59250 68340 59252
rect 68018 59220 68340 59250
rect 68018 59218 68030 59220
rect 67830 59212 68030 59218
rect 68328 59218 68340 59220
rect 68516 59218 68528 59252
rect 68328 59212 68528 59218
rect 68560 59220 68640 59240
rect 67792 59174 67800 59208
rect 67790 59160 67800 59174
rect 67720 59140 67800 59160
rect 67830 59164 68030 59170
rect 67830 59130 67842 59164
rect 68018 59160 68030 59164
rect 68328 59164 68528 59170
rect 68328 59160 68340 59164
rect 68018 59150 68340 59160
rect 68018 59130 68150 59150
rect 67830 59124 68030 59130
rect 68140 59090 68150 59130
rect 68210 59130 68340 59150
rect 68516 59130 68528 59164
rect 68560 59160 68570 59220
rect 68630 59160 68640 59220
rect 68560 59140 68640 59160
rect 68210 59090 68220 59130
rect 68328 59124 68528 59130
rect 68140 59080 68220 59090
rect 67610 57920 67680 59070
rect 67610 57660 67630 57920
rect 67670 57660 67680 57920
rect 68690 59070 68700 59310
rect 68740 59070 68760 59310
rect 68690 57920 68760 59070
rect 68140 57890 68220 57900
rect 67830 57852 68030 57858
rect 67720 57820 67800 57840
rect 67720 57760 67730 57820
rect 67790 57808 67800 57820
rect 67830 57818 67842 57852
rect 68018 57850 68030 57852
rect 68140 57850 68150 57890
rect 68018 57830 68150 57850
rect 68210 57850 68220 57890
rect 68328 57852 68528 57858
rect 68328 57850 68340 57852
rect 68210 57830 68340 57850
rect 68018 57820 68340 57830
rect 68018 57818 68030 57820
rect 67830 57812 68030 57818
rect 68328 57818 68340 57820
rect 68516 57818 68528 57852
rect 68328 57812 68528 57818
rect 68560 57820 68640 57840
rect 67792 57774 67800 57808
rect 67790 57760 67800 57774
rect 67720 57740 67800 57760
rect 67830 57764 68030 57770
rect 67830 57730 67842 57764
rect 68018 57760 68030 57764
rect 68328 57764 68528 57770
rect 68328 57760 68340 57764
rect 68018 57730 68340 57760
rect 68516 57730 68528 57764
rect 68560 57760 68570 57820
rect 68630 57760 68640 57820
rect 68560 57740 68640 57760
rect 67830 57724 68030 57730
rect 67610 57600 67680 57660
rect 67610 57360 67630 57600
rect 67670 57360 67680 57600
rect 68140 57720 68220 57730
rect 68328 57724 68528 57730
rect 68140 57660 68150 57720
rect 68210 57660 68220 57720
rect 68140 57610 68220 57660
rect 68140 57550 68150 57610
rect 68210 57550 68220 57610
rect 67830 57542 68030 57548
rect 67720 57510 67800 57530
rect 67720 57450 67730 57510
rect 67790 57498 67800 57510
rect 67830 57508 67842 57542
rect 68018 57540 68030 57542
rect 68140 57540 68220 57550
rect 68690 57680 68700 57920
rect 68740 57680 68760 57920
rect 68690 57600 68760 57680
rect 68328 57542 68528 57548
rect 68328 57540 68340 57542
rect 68018 57510 68340 57540
rect 68018 57508 68030 57510
rect 67830 57502 68030 57508
rect 68328 57508 68340 57510
rect 68516 57508 68528 57542
rect 68328 57502 68528 57508
rect 68560 57510 68640 57530
rect 67792 57464 67800 57498
rect 67790 57450 67800 57464
rect 67720 57430 67800 57450
rect 67830 57454 68030 57460
rect 67830 57420 67842 57454
rect 68018 57450 68030 57454
rect 68328 57454 68528 57460
rect 68328 57450 68340 57454
rect 68018 57440 68340 57450
rect 68018 57420 68150 57440
rect 67830 57414 68030 57420
rect 68140 57380 68150 57420
rect 68210 57420 68340 57440
rect 68516 57420 68528 57454
rect 68560 57450 68570 57510
rect 68630 57450 68640 57510
rect 68560 57430 68640 57450
rect 68210 57380 68220 57420
rect 68328 57414 68528 57420
rect 68140 57370 68220 57380
rect 67610 56210 67680 57360
rect 67610 55950 67630 56210
rect 67670 55950 67680 56210
rect 68690 57360 68700 57600
rect 68740 57360 68760 57600
rect 68690 56210 68760 57360
rect 68140 56180 68220 56190
rect 67830 56142 68030 56148
rect 67720 56110 67800 56130
rect 67720 56050 67730 56110
rect 67790 56098 67800 56110
rect 67830 56108 67842 56142
rect 68018 56140 68030 56142
rect 68140 56140 68150 56180
rect 68018 56120 68150 56140
rect 68210 56140 68220 56180
rect 68328 56142 68528 56148
rect 68328 56140 68340 56142
rect 68210 56120 68340 56140
rect 68018 56110 68340 56120
rect 68018 56108 68030 56110
rect 67830 56102 68030 56108
rect 68328 56108 68340 56110
rect 68516 56108 68528 56142
rect 68328 56102 68528 56108
rect 68560 56110 68640 56130
rect 67792 56064 67800 56098
rect 67790 56050 67800 56064
rect 67720 56030 67800 56050
rect 67830 56054 68030 56060
rect 67830 56020 67842 56054
rect 68018 56050 68030 56054
rect 68328 56054 68528 56060
rect 68328 56050 68340 56054
rect 68018 56020 68340 56050
rect 68516 56020 68528 56054
rect 68560 56050 68570 56110
rect 68630 56050 68640 56110
rect 68560 56030 68640 56050
rect 67830 56014 68030 56020
rect 67610 55890 67680 55950
rect 67610 55650 67630 55890
rect 67670 55650 67680 55890
rect 68140 56010 68220 56020
rect 68328 56014 68528 56020
rect 68140 55950 68150 56010
rect 68210 55950 68220 56010
rect 68140 55900 68220 55950
rect 68140 55840 68150 55900
rect 68210 55840 68220 55900
rect 67830 55832 68030 55838
rect 67720 55800 67800 55820
rect 67720 55740 67730 55800
rect 67790 55788 67800 55800
rect 67830 55798 67842 55832
rect 68018 55830 68030 55832
rect 68140 55830 68220 55840
rect 68690 55970 68700 56210
rect 68740 55970 68760 56210
rect 68690 55890 68760 55970
rect 68328 55832 68528 55838
rect 68328 55830 68340 55832
rect 68018 55800 68340 55830
rect 68018 55798 68030 55800
rect 67830 55792 68030 55798
rect 68328 55798 68340 55800
rect 68516 55798 68528 55832
rect 68328 55792 68528 55798
rect 68560 55800 68640 55820
rect 67792 55754 67800 55788
rect 67790 55740 67800 55754
rect 67720 55720 67800 55740
rect 67830 55744 68030 55750
rect 67830 55710 67842 55744
rect 68018 55740 68030 55744
rect 68328 55744 68528 55750
rect 68328 55740 68340 55744
rect 68018 55730 68340 55740
rect 68018 55710 68150 55730
rect 67830 55704 68030 55710
rect 68140 55670 68150 55710
rect 68210 55710 68340 55730
rect 68516 55710 68528 55744
rect 68560 55740 68570 55800
rect 68630 55740 68640 55800
rect 68560 55720 68640 55740
rect 68210 55670 68220 55710
rect 68328 55704 68528 55710
rect 68140 55660 68220 55670
rect 67610 54500 67680 55650
rect 67610 54240 67630 54500
rect 67670 54240 67680 54500
rect 68690 55650 68700 55890
rect 68740 55650 68760 55890
rect 68690 54500 68760 55650
rect 68140 54470 68220 54480
rect 67830 54432 68030 54438
rect 67720 54400 67800 54420
rect 67720 54340 67730 54400
rect 67790 54388 67800 54400
rect 67830 54398 67842 54432
rect 68018 54430 68030 54432
rect 68140 54430 68150 54470
rect 68018 54410 68150 54430
rect 68210 54430 68220 54470
rect 68328 54432 68528 54438
rect 68328 54430 68340 54432
rect 68210 54410 68340 54430
rect 68018 54400 68340 54410
rect 68018 54398 68030 54400
rect 67830 54392 68030 54398
rect 68328 54398 68340 54400
rect 68516 54398 68528 54432
rect 68328 54392 68528 54398
rect 68560 54400 68640 54420
rect 67792 54354 67800 54388
rect 67790 54340 67800 54354
rect 67720 54320 67800 54340
rect 67830 54344 68030 54350
rect 67830 54310 67842 54344
rect 68018 54340 68030 54344
rect 68328 54344 68528 54350
rect 68328 54340 68340 54344
rect 68018 54310 68340 54340
rect 68516 54310 68528 54344
rect 68560 54340 68570 54400
rect 68630 54340 68640 54400
rect 68560 54320 68640 54340
rect 67830 54304 68030 54310
rect 67610 54180 67680 54240
rect 67610 53940 67630 54180
rect 67670 53940 67680 54180
rect 68140 54300 68220 54310
rect 68328 54304 68528 54310
rect 68140 54240 68150 54300
rect 68210 54240 68220 54300
rect 68140 54190 68220 54240
rect 68140 54130 68150 54190
rect 68210 54130 68220 54190
rect 67830 54122 68030 54128
rect 67720 54090 67800 54110
rect 67720 54030 67730 54090
rect 67790 54078 67800 54090
rect 67830 54088 67842 54122
rect 68018 54120 68030 54122
rect 68140 54120 68220 54130
rect 68690 54260 68700 54500
rect 68740 54260 68760 54500
rect 68690 54180 68760 54260
rect 68328 54122 68528 54128
rect 68328 54120 68340 54122
rect 68018 54090 68340 54120
rect 68018 54088 68030 54090
rect 67830 54082 68030 54088
rect 68328 54088 68340 54090
rect 68516 54088 68528 54122
rect 68328 54082 68528 54088
rect 68560 54090 68640 54110
rect 67792 54044 67800 54078
rect 67790 54030 67800 54044
rect 67720 54010 67800 54030
rect 67830 54034 68030 54040
rect 67830 54000 67842 54034
rect 68018 54030 68030 54034
rect 68328 54034 68528 54040
rect 68328 54030 68340 54034
rect 68018 54020 68340 54030
rect 68018 54000 68150 54020
rect 67830 53994 68030 54000
rect 68140 53960 68150 54000
rect 68210 54000 68340 54020
rect 68516 54000 68528 54034
rect 68560 54030 68570 54090
rect 68630 54030 68640 54090
rect 68560 54010 68640 54030
rect 68210 53960 68220 54000
rect 68328 53994 68528 54000
rect 68140 53950 68220 53960
rect 67610 52790 67680 53940
rect 67610 52530 67630 52790
rect 67670 52530 67680 52790
rect 68690 53940 68700 54180
rect 68740 53940 68760 54180
rect 68690 52790 68760 53940
rect 68140 52760 68220 52770
rect 67830 52722 68030 52728
rect 67720 52690 67800 52710
rect 67720 52630 67730 52690
rect 67790 52678 67800 52690
rect 67830 52688 67842 52722
rect 68018 52720 68030 52722
rect 68140 52720 68150 52760
rect 68018 52700 68150 52720
rect 68210 52720 68220 52760
rect 68328 52722 68528 52728
rect 68328 52720 68340 52722
rect 68210 52700 68340 52720
rect 68018 52690 68340 52700
rect 68018 52688 68030 52690
rect 67830 52682 68030 52688
rect 68328 52688 68340 52690
rect 68516 52688 68528 52722
rect 68328 52682 68528 52688
rect 68560 52690 68640 52710
rect 67792 52644 67800 52678
rect 67790 52630 67800 52644
rect 67720 52610 67800 52630
rect 67830 52634 68030 52640
rect 67830 52600 67842 52634
rect 68018 52630 68030 52634
rect 68328 52634 68528 52640
rect 68328 52630 68340 52634
rect 68018 52600 68340 52630
rect 68516 52600 68528 52634
rect 68560 52630 68570 52690
rect 68630 52630 68640 52690
rect 68560 52610 68640 52630
rect 67830 52594 68030 52600
rect 67610 52470 67680 52530
rect 67610 52230 67630 52470
rect 67670 52230 67680 52470
rect 68140 52590 68220 52600
rect 68328 52594 68528 52600
rect 68140 52530 68150 52590
rect 68210 52530 68220 52590
rect 68140 52480 68220 52530
rect 68140 52420 68150 52480
rect 68210 52420 68220 52480
rect 67830 52412 68030 52418
rect 67720 52380 67800 52400
rect 67720 52320 67730 52380
rect 67790 52368 67800 52380
rect 67830 52378 67842 52412
rect 68018 52410 68030 52412
rect 68140 52410 68220 52420
rect 68690 52550 68700 52790
rect 68740 52550 68760 52790
rect 68690 52470 68760 52550
rect 68328 52412 68528 52418
rect 68328 52410 68340 52412
rect 68018 52380 68340 52410
rect 68018 52378 68030 52380
rect 67830 52372 68030 52378
rect 68328 52378 68340 52380
rect 68516 52378 68528 52412
rect 68328 52372 68528 52378
rect 68560 52380 68640 52400
rect 67792 52334 67800 52368
rect 67790 52320 67800 52334
rect 67720 52300 67800 52320
rect 67830 52324 68030 52330
rect 67830 52290 67842 52324
rect 68018 52320 68030 52324
rect 68328 52324 68528 52330
rect 68328 52320 68340 52324
rect 68018 52310 68340 52320
rect 68018 52290 68150 52310
rect 67830 52284 68030 52290
rect 68140 52250 68150 52290
rect 68210 52290 68340 52310
rect 68516 52290 68528 52324
rect 68560 52320 68570 52380
rect 68630 52320 68640 52380
rect 68560 52300 68640 52320
rect 68210 52250 68220 52290
rect 68328 52284 68528 52290
rect 68140 52240 68220 52250
rect 67610 51080 67680 52230
rect 67610 50820 67630 51080
rect 67670 50820 67680 51080
rect 68690 52230 68700 52470
rect 68740 52230 68760 52470
rect 68690 51080 68760 52230
rect 68140 51050 68220 51060
rect 67830 51012 68030 51018
rect 67720 50980 67800 51000
rect 67720 50920 67730 50980
rect 67790 50968 67800 50980
rect 67830 50978 67842 51012
rect 68018 51010 68030 51012
rect 68140 51010 68150 51050
rect 68018 50990 68150 51010
rect 68210 51010 68220 51050
rect 68328 51012 68528 51018
rect 68328 51010 68340 51012
rect 68210 50990 68340 51010
rect 68018 50980 68340 50990
rect 68018 50978 68030 50980
rect 67830 50972 68030 50978
rect 68328 50978 68340 50980
rect 68516 50978 68528 51012
rect 68328 50972 68528 50978
rect 68560 50980 68640 51000
rect 67792 50934 67800 50968
rect 67790 50920 67800 50934
rect 67720 50900 67800 50920
rect 67830 50924 68030 50930
rect 67830 50890 67842 50924
rect 68018 50920 68030 50924
rect 68328 50924 68528 50930
rect 68328 50920 68340 50924
rect 68018 50890 68340 50920
rect 68516 50890 68528 50924
rect 68560 50920 68570 50980
rect 68630 50920 68640 50980
rect 68560 50900 68640 50920
rect 67830 50884 68030 50890
rect 67610 50760 67680 50820
rect 67610 50520 67630 50760
rect 67670 50520 67680 50760
rect 68140 50880 68220 50890
rect 68328 50884 68528 50890
rect 68140 50820 68150 50880
rect 68210 50820 68220 50880
rect 68140 50770 68220 50820
rect 68140 50710 68150 50770
rect 68210 50710 68220 50770
rect 67830 50702 68030 50708
rect 67720 50670 67800 50690
rect 67720 50610 67730 50670
rect 67790 50658 67800 50670
rect 67830 50668 67842 50702
rect 68018 50700 68030 50702
rect 68140 50700 68220 50710
rect 68690 50840 68700 51080
rect 68740 50840 68760 51080
rect 68690 50760 68760 50840
rect 68328 50702 68528 50708
rect 68328 50700 68340 50702
rect 68018 50670 68340 50700
rect 68018 50668 68030 50670
rect 67830 50662 68030 50668
rect 68328 50668 68340 50670
rect 68516 50668 68528 50702
rect 68328 50662 68528 50668
rect 68560 50670 68640 50690
rect 67792 50624 67800 50658
rect 67790 50610 67800 50624
rect 67720 50590 67800 50610
rect 67830 50614 68030 50620
rect 67830 50580 67842 50614
rect 68018 50610 68030 50614
rect 68328 50614 68528 50620
rect 68328 50610 68340 50614
rect 68018 50600 68340 50610
rect 68018 50580 68150 50600
rect 67830 50574 68030 50580
rect 68140 50540 68150 50580
rect 68210 50580 68340 50600
rect 68516 50580 68528 50614
rect 68560 50610 68570 50670
rect 68630 50610 68640 50670
rect 68560 50590 68640 50610
rect 68210 50540 68220 50580
rect 68328 50574 68528 50580
rect 68140 50530 68220 50540
rect 67610 49370 67680 50520
rect 67610 49110 67630 49370
rect 67670 49110 67680 49370
rect 68690 50520 68700 50760
rect 68740 50520 68760 50760
rect 68690 49370 68760 50520
rect 68140 49340 68220 49350
rect 67830 49302 68030 49308
rect 67720 49270 67800 49290
rect 67720 49210 67730 49270
rect 67790 49258 67800 49270
rect 67830 49268 67842 49302
rect 68018 49300 68030 49302
rect 68140 49300 68150 49340
rect 68018 49280 68150 49300
rect 68210 49300 68220 49340
rect 68328 49302 68528 49308
rect 68328 49300 68340 49302
rect 68210 49280 68340 49300
rect 68018 49270 68340 49280
rect 68018 49268 68030 49270
rect 67830 49262 68030 49268
rect 68328 49268 68340 49270
rect 68516 49268 68528 49302
rect 68328 49262 68528 49268
rect 68560 49270 68640 49290
rect 67792 49224 67800 49258
rect 67790 49210 67800 49224
rect 67720 49190 67800 49210
rect 67830 49214 68030 49220
rect 67830 49180 67842 49214
rect 68018 49210 68030 49214
rect 68328 49214 68528 49220
rect 68328 49210 68340 49214
rect 68018 49180 68340 49210
rect 68516 49180 68528 49214
rect 68560 49210 68570 49270
rect 68630 49210 68640 49270
rect 68560 49190 68640 49210
rect 67830 49174 68030 49180
rect 67610 49050 67680 49110
rect 67610 48810 67630 49050
rect 67670 48810 67680 49050
rect 68140 49170 68220 49180
rect 68328 49174 68528 49180
rect 68140 49110 68150 49170
rect 68210 49110 68220 49170
rect 68140 49060 68220 49110
rect 68140 49000 68150 49060
rect 68210 49000 68220 49060
rect 67830 48992 68030 48998
rect 67720 48960 67800 48980
rect 67720 48900 67730 48960
rect 67790 48948 67800 48960
rect 67830 48958 67842 48992
rect 68018 48990 68030 48992
rect 68140 48990 68220 49000
rect 68690 49130 68700 49370
rect 68740 49130 68760 49370
rect 68690 49050 68760 49130
rect 68328 48992 68528 48998
rect 68328 48990 68340 48992
rect 68018 48960 68340 48990
rect 68018 48958 68030 48960
rect 67830 48952 68030 48958
rect 68328 48958 68340 48960
rect 68516 48958 68528 48992
rect 68328 48952 68528 48958
rect 68560 48960 68640 48980
rect 67792 48914 67800 48948
rect 67790 48900 67800 48914
rect 67720 48880 67800 48900
rect 67830 48904 68030 48910
rect 67830 48870 67842 48904
rect 68018 48900 68030 48904
rect 68328 48904 68528 48910
rect 68328 48900 68340 48904
rect 68018 48890 68340 48900
rect 68018 48870 68150 48890
rect 67830 48864 68030 48870
rect 68140 48830 68150 48870
rect 68210 48870 68340 48890
rect 68516 48870 68528 48904
rect 68560 48900 68570 48960
rect 68630 48900 68640 48960
rect 68560 48880 68640 48900
rect 68210 48830 68220 48870
rect 68328 48864 68528 48870
rect 68140 48820 68220 48830
rect 67610 47660 67680 48810
rect 67610 47400 67630 47660
rect 67670 47400 67680 47660
rect 68690 48810 68700 49050
rect 68740 48810 68760 49050
rect 68690 47660 68760 48810
rect 68140 47630 68220 47640
rect 67830 47592 68030 47598
rect 67720 47560 67800 47580
rect 67720 47500 67730 47560
rect 67790 47548 67800 47560
rect 67830 47558 67842 47592
rect 68018 47590 68030 47592
rect 68140 47590 68150 47630
rect 68018 47570 68150 47590
rect 68210 47590 68220 47630
rect 68328 47592 68528 47598
rect 68328 47590 68340 47592
rect 68210 47570 68340 47590
rect 68018 47560 68340 47570
rect 68018 47558 68030 47560
rect 67830 47552 68030 47558
rect 68328 47558 68340 47560
rect 68516 47558 68528 47592
rect 68328 47552 68528 47558
rect 68560 47560 68640 47580
rect 67792 47514 67800 47548
rect 67790 47500 67800 47514
rect 67720 47480 67800 47500
rect 67830 47504 68030 47510
rect 67830 47470 67842 47504
rect 68018 47500 68030 47504
rect 68328 47504 68528 47510
rect 68328 47500 68340 47504
rect 68018 47470 68340 47500
rect 68516 47470 68528 47504
rect 68560 47500 68570 47560
rect 68630 47500 68640 47560
rect 68560 47480 68640 47500
rect 67830 47464 68030 47470
rect 67610 47340 67680 47400
rect 67610 47100 67630 47340
rect 67670 47100 67680 47340
rect 68140 47460 68220 47470
rect 68328 47464 68528 47470
rect 68140 47400 68150 47460
rect 68210 47400 68220 47460
rect 68140 47350 68220 47400
rect 68140 47290 68150 47350
rect 68210 47290 68220 47350
rect 67830 47282 68030 47288
rect 67720 47250 67800 47270
rect 67720 47190 67730 47250
rect 67790 47238 67800 47250
rect 67830 47248 67842 47282
rect 68018 47280 68030 47282
rect 68140 47280 68220 47290
rect 68690 47420 68700 47660
rect 68740 47420 68760 47660
rect 68690 47340 68760 47420
rect 68328 47282 68528 47288
rect 68328 47280 68340 47282
rect 68018 47250 68340 47280
rect 68018 47248 68030 47250
rect 67830 47242 68030 47248
rect 68328 47248 68340 47250
rect 68516 47248 68528 47282
rect 68328 47242 68528 47248
rect 68560 47250 68640 47270
rect 67792 47204 67800 47238
rect 67790 47190 67800 47204
rect 67720 47170 67800 47190
rect 67830 47194 68030 47200
rect 67830 47160 67842 47194
rect 68018 47190 68030 47194
rect 68328 47194 68528 47200
rect 68328 47190 68340 47194
rect 68018 47180 68340 47190
rect 68018 47160 68150 47180
rect 67830 47154 68030 47160
rect 68140 47120 68150 47160
rect 68210 47160 68340 47180
rect 68516 47160 68528 47194
rect 68560 47190 68570 47250
rect 68630 47190 68640 47250
rect 68560 47170 68640 47190
rect 68210 47120 68220 47160
rect 68328 47154 68528 47160
rect 68140 47110 68220 47120
rect 67610 45950 67680 47100
rect 67610 45690 67630 45950
rect 67670 45690 67680 45950
rect 68690 47100 68700 47340
rect 68740 47100 68760 47340
rect 68690 45950 68760 47100
rect 68140 45920 68220 45930
rect 67830 45882 68030 45888
rect 67720 45850 67800 45870
rect 67720 45790 67730 45850
rect 67790 45838 67800 45850
rect 67830 45848 67842 45882
rect 68018 45880 68030 45882
rect 68140 45880 68150 45920
rect 68018 45860 68150 45880
rect 68210 45880 68220 45920
rect 68328 45882 68528 45888
rect 68328 45880 68340 45882
rect 68210 45860 68340 45880
rect 68018 45850 68340 45860
rect 68018 45848 68030 45850
rect 67830 45842 68030 45848
rect 68328 45848 68340 45850
rect 68516 45848 68528 45882
rect 68328 45842 68528 45848
rect 68560 45850 68640 45870
rect 67792 45804 67800 45838
rect 67790 45790 67800 45804
rect 67720 45770 67800 45790
rect 67830 45794 68030 45800
rect 67830 45760 67842 45794
rect 68018 45790 68030 45794
rect 68328 45794 68528 45800
rect 68328 45790 68340 45794
rect 68018 45760 68340 45790
rect 68516 45760 68528 45794
rect 68560 45790 68570 45850
rect 68630 45790 68640 45850
rect 68560 45770 68640 45790
rect 67830 45754 68030 45760
rect 67610 45630 67680 45690
rect 67610 45390 67630 45630
rect 67670 45390 67680 45630
rect 68140 45750 68220 45760
rect 68328 45754 68528 45760
rect 68140 45690 68150 45750
rect 68210 45690 68220 45750
rect 68140 45640 68220 45690
rect 68140 45580 68150 45640
rect 68210 45580 68220 45640
rect 67830 45572 68030 45578
rect 67720 45540 67800 45560
rect 67720 45480 67730 45540
rect 67790 45528 67800 45540
rect 67830 45538 67842 45572
rect 68018 45570 68030 45572
rect 68140 45570 68220 45580
rect 68690 45710 68700 45950
rect 68740 45710 68760 45950
rect 68690 45630 68760 45710
rect 68328 45572 68528 45578
rect 68328 45570 68340 45572
rect 68018 45540 68340 45570
rect 68018 45538 68030 45540
rect 67830 45532 68030 45538
rect 68328 45538 68340 45540
rect 68516 45538 68528 45572
rect 68328 45532 68528 45538
rect 68560 45540 68640 45560
rect 67792 45494 67800 45528
rect 67790 45480 67800 45494
rect 67720 45460 67800 45480
rect 67830 45484 68030 45490
rect 67830 45450 67842 45484
rect 68018 45480 68030 45484
rect 68328 45484 68528 45490
rect 68328 45480 68340 45484
rect 68018 45470 68340 45480
rect 68018 45450 68150 45470
rect 67830 45444 68030 45450
rect 68140 45410 68150 45450
rect 68210 45450 68340 45470
rect 68516 45450 68528 45484
rect 68560 45480 68570 45540
rect 68630 45480 68640 45540
rect 68560 45460 68640 45480
rect 68210 45410 68220 45450
rect 68328 45444 68528 45450
rect 68140 45400 68220 45410
rect 67610 44240 67680 45390
rect 67610 43980 67630 44240
rect 67670 43980 67680 44240
rect 68690 45390 68700 45630
rect 68740 45390 68760 45630
rect 68690 44240 68760 45390
rect 68140 44210 68220 44220
rect 67830 44172 68030 44178
rect 67720 44140 67800 44160
rect 67720 44080 67730 44140
rect 67790 44128 67800 44140
rect 67830 44138 67842 44172
rect 68018 44170 68030 44172
rect 68140 44170 68150 44210
rect 68018 44150 68150 44170
rect 68210 44170 68220 44210
rect 68328 44172 68528 44178
rect 68328 44170 68340 44172
rect 68210 44150 68340 44170
rect 68018 44140 68340 44150
rect 68018 44138 68030 44140
rect 67830 44132 68030 44138
rect 68328 44138 68340 44140
rect 68516 44138 68528 44172
rect 68328 44132 68528 44138
rect 68560 44140 68640 44160
rect 67792 44094 67800 44128
rect 67790 44080 67800 44094
rect 67720 44060 67800 44080
rect 67830 44084 68030 44090
rect 67830 44050 67842 44084
rect 68018 44080 68030 44084
rect 68328 44084 68528 44090
rect 68328 44080 68340 44084
rect 68018 44050 68340 44080
rect 68516 44050 68528 44084
rect 68560 44080 68570 44140
rect 68630 44080 68640 44140
rect 68560 44060 68640 44080
rect 67830 44044 68030 44050
rect 67610 43920 67680 43980
rect 67610 43680 67630 43920
rect 67670 43680 67680 43920
rect 68140 44040 68220 44050
rect 68328 44044 68528 44050
rect 68140 43980 68150 44040
rect 68210 43980 68220 44040
rect 68140 43930 68220 43980
rect 68140 43870 68150 43930
rect 68210 43870 68220 43930
rect 67830 43862 68030 43868
rect 67720 43830 67800 43850
rect 67720 43770 67730 43830
rect 67790 43818 67800 43830
rect 67830 43828 67842 43862
rect 68018 43860 68030 43862
rect 68140 43860 68220 43870
rect 68690 44000 68700 44240
rect 68740 44000 68760 44240
rect 68690 43920 68760 44000
rect 68328 43862 68528 43868
rect 68328 43860 68340 43862
rect 68018 43830 68340 43860
rect 68018 43828 68030 43830
rect 67830 43822 68030 43828
rect 68328 43828 68340 43830
rect 68516 43828 68528 43862
rect 68328 43822 68528 43828
rect 68560 43830 68640 43850
rect 67792 43784 67800 43818
rect 67790 43770 67800 43784
rect 67720 43750 67800 43770
rect 67830 43774 68030 43780
rect 67830 43740 67842 43774
rect 68018 43770 68030 43774
rect 68328 43774 68528 43780
rect 68328 43770 68340 43774
rect 68018 43760 68340 43770
rect 68018 43740 68150 43760
rect 67830 43734 68030 43740
rect 68140 43700 68150 43740
rect 68210 43740 68340 43760
rect 68516 43740 68528 43774
rect 68560 43770 68570 43830
rect 68630 43770 68640 43830
rect 68560 43750 68640 43770
rect 68210 43700 68220 43740
rect 68328 43734 68528 43740
rect 68140 43690 68220 43700
rect 67610 42530 67680 43680
rect 67610 42270 67630 42530
rect 67670 42270 67680 42530
rect 68690 43680 68700 43920
rect 68740 43680 68760 43920
rect 68690 42530 68760 43680
rect 68140 42500 68220 42510
rect 67830 42462 68030 42468
rect 67720 42430 67800 42450
rect 67720 42370 67730 42430
rect 67790 42418 67800 42430
rect 67830 42428 67842 42462
rect 68018 42460 68030 42462
rect 68140 42460 68150 42500
rect 68018 42440 68150 42460
rect 68210 42460 68220 42500
rect 68328 42462 68528 42468
rect 68328 42460 68340 42462
rect 68210 42440 68340 42460
rect 68018 42430 68340 42440
rect 68018 42428 68030 42430
rect 67830 42422 68030 42428
rect 68328 42428 68340 42430
rect 68516 42428 68528 42462
rect 68328 42422 68528 42428
rect 68560 42430 68640 42450
rect 67792 42384 67800 42418
rect 67790 42370 67800 42384
rect 67720 42350 67800 42370
rect 67830 42374 68030 42380
rect 67830 42340 67842 42374
rect 68018 42370 68030 42374
rect 68328 42374 68528 42380
rect 68328 42370 68340 42374
rect 68018 42340 68340 42370
rect 68516 42340 68528 42374
rect 68560 42370 68570 42430
rect 68630 42370 68640 42430
rect 68560 42350 68640 42370
rect 67830 42334 68030 42340
rect 67610 42210 67680 42270
rect 67610 41970 67630 42210
rect 67670 41970 67680 42210
rect 68140 42330 68220 42340
rect 68328 42334 68528 42340
rect 68140 42270 68150 42330
rect 68210 42270 68220 42330
rect 68140 42220 68220 42270
rect 68140 42160 68150 42220
rect 68210 42160 68220 42220
rect 67830 42152 68030 42158
rect 67720 42120 67800 42140
rect 67720 42060 67730 42120
rect 67790 42108 67800 42120
rect 67830 42118 67842 42152
rect 68018 42150 68030 42152
rect 68140 42150 68220 42160
rect 68690 42290 68700 42530
rect 68740 42290 68760 42530
rect 68690 42210 68760 42290
rect 68328 42152 68528 42158
rect 68328 42150 68340 42152
rect 68018 42120 68340 42150
rect 68018 42118 68030 42120
rect 67830 42112 68030 42118
rect 68328 42118 68340 42120
rect 68516 42118 68528 42152
rect 68328 42112 68528 42118
rect 68560 42120 68640 42140
rect 67792 42074 67800 42108
rect 67790 42060 67800 42074
rect 67720 42040 67800 42060
rect 67830 42064 68030 42070
rect 67830 42030 67842 42064
rect 68018 42060 68030 42064
rect 68328 42064 68528 42070
rect 68328 42060 68340 42064
rect 68018 42050 68340 42060
rect 68018 42030 68150 42050
rect 67830 42024 68030 42030
rect 68140 41990 68150 42030
rect 68210 42030 68340 42050
rect 68516 42030 68528 42064
rect 68560 42060 68570 42120
rect 68630 42060 68640 42120
rect 68560 42040 68640 42060
rect 68210 41990 68220 42030
rect 68328 42024 68528 42030
rect 68140 41980 68220 41990
rect 67610 40820 67680 41970
rect 67610 40560 67630 40820
rect 67670 40560 67680 40820
rect 68690 41970 68700 42210
rect 68740 41970 68760 42210
rect 68690 40820 68760 41970
rect 68140 40790 68220 40800
rect 67830 40752 68030 40758
rect 67720 40720 67800 40740
rect 67720 40660 67730 40720
rect 67790 40708 67800 40720
rect 67830 40718 67842 40752
rect 68018 40750 68030 40752
rect 68140 40750 68150 40790
rect 68018 40730 68150 40750
rect 68210 40750 68220 40790
rect 68328 40752 68528 40758
rect 68328 40750 68340 40752
rect 68210 40730 68340 40750
rect 68018 40720 68340 40730
rect 68018 40718 68030 40720
rect 67830 40712 68030 40718
rect 68328 40718 68340 40720
rect 68516 40718 68528 40752
rect 68328 40712 68528 40718
rect 68560 40720 68640 40740
rect 67792 40674 67800 40708
rect 67790 40660 67800 40674
rect 67720 40640 67800 40660
rect 67830 40664 68030 40670
rect 67830 40630 67842 40664
rect 68018 40660 68030 40664
rect 68328 40664 68528 40670
rect 68328 40660 68340 40664
rect 68018 40630 68340 40660
rect 68516 40630 68528 40664
rect 68560 40660 68570 40720
rect 68630 40660 68640 40720
rect 68560 40640 68640 40660
rect 67830 40624 68030 40630
rect 67610 40500 67680 40560
rect 67610 40260 67630 40500
rect 67670 40260 67680 40500
rect 68140 40620 68220 40630
rect 68328 40624 68528 40630
rect 68140 40560 68150 40620
rect 68210 40560 68220 40620
rect 68140 40510 68220 40560
rect 68140 40450 68150 40510
rect 68210 40450 68220 40510
rect 67830 40442 68030 40448
rect 67720 40410 67800 40430
rect 67720 40350 67730 40410
rect 67790 40398 67800 40410
rect 67830 40408 67842 40442
rect 68018 40440 68030 40442
rect 68140 40440 68220 40450
rect 68690 40580 68700 40820
rect 68740 40580 68760 40820
rect 68690 40500 68760 40580
rect 68328 40442 68528 40448
rect 68328 40440 68340 40442
rect 68018 40410 68340 40440
rect 68018 40408 68030 40410
rect 67830 40402 68030 40408
rect 68328 40408 68340 40410
rect 68516 40408 68528 40442
rect 68328 40402 68528 40408
rect 68560 40410 68640 40430
rect 67792 40364 67800 40398
rect 67790 40350 67800 40364
rect 67720 40330 67800 40350
rect 67830 40354 68030 40360
rect 67830 40320 67842 40354
rect 68018 40350 68030 40354
rect 68328 40354 68528 40360
rect 68328 40350 68340 40354
rect 68018 40340 68340 40350
rect 68018 40320 68150 40340
rect 67830 40314 68030 40320
rect 68140 40280 68150 40320
rect 68210 40320 68340 40340
rect 68516 40320 68528 40354
rect 68560 40350 68570 40410
rect 68630 40350 68640 40410
rect 68560 40330 68640 40350
rect 68210 40280 68220 40320
rect 68328 40314 68528 40320
rect 68140 40270 68220 40280
rect 67610 39690 67680 40260
rect 68690 40260 68700 40500
rect 68740 40260 68760 40500
rect 68690 39690 68760 40260
rect 67610 39680 67690 39690
rect 67610 39620 67620 39680
rect 67680 39620 67690 39680
rect 68680 39680 68760 39690
rect 68680 39620 68690 39680
rect 68750 39620 68760 39680
rect 68680 39610 68760 39620
rect 68790 66480 68820 67050
rect 68790 66470 68850 66480
rect 68790 66400 68850 66410
rect 68790 64770 68820 66400
rect 68880 65950 68910 67050
rect 68850 65940 68910 65950
rect 68850 65870 68910 65880
rect 68790 64760 68850 64770
rect 68790 64690 68850 64700
rect 68790 63060 68820 64690
rect 68880 64240 68910 65870
rect 68850 64230 68910 64240
rect 68850 64160 68910 64170
rect 68790 63050 68850 63060
rect 68790 62980 68850 62990
rect 68790 61350 68820 62980
rect 68880 62530 68910 64160
rect 68850 62520 68910 62530
rect 68850 62450 68910 62460
rect 68790 61340 68850 61350
rect 68790 61270 68850 61280
rect 68790 59640 68820 61270
rect 68880 60820 68910 62450
rect 68850 60810 68910 60820
rect 68850 60740 68910 60750
rect 68790 59630 68850 59640
rect 68790 59560 68850 59570
rect 68790 57930 68820 59560
rect 68880 59110 68910 60740
rect 68850 59100 68910 59110
rect 68850 59030 68910 59040
rect 68790 57920 68850 57930
rect 68790 57850 68850 57860
rect 68790 56220 68820 57850
rect 68880 57400 68910 59030
rect 68850 57390 68910 57400
rect 68850 57320 68910 57330
rect 68790 56210 68850 56220
rect 68790 56140 68850 56150
rect 68790 54510 68820 56140
rect 68880 55690 68910 57320
rect 68850 55680 68910 55690
rect 68850 55610 68910 55620
rect 68790 54500 68850 54510
rect 68790 54430 68850 54440
rect 68790 52800 68820 54430
rect 68880 53980 68910 55610
rect 68850 53970 68910 53980
rect 68850 53900 68910 53910
rect 68790 52790 68850 52800
rect 68790 52720 68850 52730
rect 68790 51090 68820 52720
rect 68880 52270 68910 53900
rect 68850 52260 68910 52270
rect 68850 52190 68910 52200
rect 68790 51080 68850 51090
rect 68790 51010 68850 51020
rect 68790 49380 68820 51010
rect 68880 50560 68910 52190
rect 68850 50550 68910 50560
rect 68850 50480 68910 50490
rect 68790 49370 68850 49380
rect 68790 49300 68850 49310
rect 68790 47670 68820 49300
rect 68880 48850 68910 50480
rect 68850 48840 68910 48850
rect 68850 48770 68910 48780
rect 68790 47660 68850 47670
rect 68790 47590 68850 47600
rect 68790 45960 68820 47590
rect 68880 47140 68910 48770
rect 68850 47130 68910 47140
rect 68850 47060 68910 47070
rect 68790 45950 68850 45960
rect 68790 45880 68850 45890
rect 68790 44250 68820 45880
rect 68880 45430 68910 47060
rect 68850 45420 68910 45430
rect 68850 45350 68910 45360
rect 68790 44240 68850 44250
rect 68790 44170 68850 44180
rect 68790 42540 68820 44170
rect 68880 43720 68910 45350
rect 68850 43710 68910 43720
rect 68850 43640 68910 43650
rect 68790 42530 68850 42540
rect 68790 42460 68850 42470
rect 68790 40830 68820 42460
rect 68880 42010 68910 43640
rect 68850 42000 68910 42010
rect 68850 41930 68910 41940
rect 68790 40820 68850 40830
rect 68790 40750 68850 40760
rect 67140 39220 67200 39230
rect 67320 39230 67580 39240
rect 64150 39160 64210 39170
rect 67380 39210 67580 39230
rect 67320 39160 67380 39170
rect 68790 38840 68820 40750
rect 68880 40300 68910 41930
rect 68850 40290 68910 40300
rect 68850 40220 68910 40230
rect 68880 39690 68910 40220
rect 68850 39680 68910 39690
rect 68850 39610 68910 39620
rect 68940 66390 68970 67050
rect 68940 66380 69000 66390
rect 68940 66310 69000 66320
rect 68940 64680 68970 66310
rect 68940 64670 69000 64680
rect 68940 64600 69000 64610
rect 68940 62970 68970 64600
rect 68940 62960 69000 62970
rect 68940 62890 69000 62900
rect 68940 61260 68970 62890
rect 68940 61250 69000 61260
rect 68940 61180 69000 61190
rect 68940 45870 68970 61180
rect 69060 59550 69090 67050
rect 69060 59540 69120 59550
rect 69060 59470 69120 59480
rect 69060 57840 69090 59470
rect 69060 57830 69120 57840
rect 69060 57760 69120 57770
rect 69060 56130 69090 57760
rect 69060 56120 69120 56130
rect 69060 56050 69120 56060
rect 69060 54420 69090 56050
rect 69060 54410 69120 54420
rect 69060 54340 69120 54350
rect 69060 52710 69090 54340
rect 69060 52700 69120 52710
rect 69060 52630 69120 52640
rect 69060 51000 69090 52630
rect 69060 50990 69120 51000
rect 69060 50920 69120 50930
rect 69060 49290 69090 50920
rect 69060 49280 69120 49290
rect 69060 49210 69120 49220
rect 69060 47580 69090 49210
rect 69060 47570 69120 47580
rect 69060 47500 69120 47510
rect 68940 45860 69000 45870
rect 68940 45790 69000 45800
rect 68940 44160 68970 45790
rect 68940 44150 69000 44160
rect 68940 44080 69000 44090
rect 68940 42450 68970 44080
rect 68940 42440 69000 42450
rect 68940 42370 69000 42380
rect 68940 40740 68970 42370
rect 68940 40730 69000 40740
rect 68940 40660 69000 40670
rect 68940 39240 68970 40660
rect 69060 39300 69090 47500
rect 69180 39690 69210 67050
rect 69300 39690 69330 67050
rect 69420 39690 69450 67050
rect 69540 39690 69570 67050
rect 69660 39690 69690 67050
rect 71820 39690 71850 67050
rect 71940 39690 71970 67050
rect 72060 39690 72090 67050
rect 72180 39690 72210 67050
rect 72300 39690 72330 67050
rect 72420 39690 72450 67050
rect 72540 66390 72570 67050
rect 72510 66380 72570 66390
rect 72510 66310 72570 66320
rect 72540 64680 72570 66310
rect 72510 64670 72570 64680
rect 72510 64600 72570 64610
rect 72540 62970 72570 64600
rect 72510 62960 72570 62970
rect 72510 62890 72570 62900
rect 72540 61260 72570 62890
rect 72510 61250 72570 61260
rect 72510 61180 72570 61190
rect 72540 59550 72570 61180
rect 72510 59540 72570 59550
rect 72510 59470 72570 59480
rect 72540 57840 72570 59470
rect 72510 57830 72570 57840
rect 72510 57760 72570 57770
rect 72540 56130 72570 57760
rect 72510 56120 72570 56130
rect 72510 56050 72570 56060
rect 72540 54420 72570 56050
rect 72510 54410 72570 54420
rect 72510 54340 72570 54350
rect 72540 52710 72570 54340
rect 72510 52700 72570 52710
rect 72510 52630 72570 52640
rect 72540 51000 72570 52630
rect 72510 50990 72570 51000
rect 72510 50920 72570 50930
rect 72540 49290 72570 50920
rect 72510 49280 72570 49290
rect 72510 49210 72570 49220
rect 72540 47580 72570 49210
rect 72510 47570 72570 47580
rect 72510 47500 72570 47510
rect 72540 45870 72570 47500
rect 72510 45860 72570 45870
rect 72510 45790 72570 45800
rect 72540 44160 72570 45790
rect 72510 44150 72570 44160
rect 72510 44080 72570 44090
rect 72540 42450 72570 44080
rect 72510 42440 72570 42450
rect 72510 42370 72570 42380
rect 72540 40740 72570 42370
rect 72510 40730 72570 40740
rect 72510 40660 72570 40670
rect 69060 39290 69380 39300
rect 69060 39270 69320 39290
rect 68940 39230 69200 39240
rect 68940 39210 69140 39230
rect 72540 39240 72570 40660
rect 72600 66470 72670 67050
rect 72600 66210 72620 66470
rect 72660 66210 72670 66470
rect 73680 66470 73750 67050
rect 73130 66440 73210 66450
rect 72820 66402 73020 66408
rect 72710 66370 72790 66390
rect 72710 66310 72720 66370
rect 72780 66358 72790 66370
rect 72820 66368 72832 66402
rect 73008 66400 73020 66402
rect 73130 66400 73140 66440
rect 73008 66380 73140 66400
rect 73200 66400 73210 66440
rect 73318 66402 73518 66408
rect 73318 66400 73330 66402
rect 73200 66380 73330 66400
rect 73008 66370 73330 66380
rect 73008 66368 73020 66370
rect 72820 66362 73020 66368
rect 73318 66368 73330 66370
rect 73506 66368 73518 66402
rect 73318 66362 73518 66368
rect 73550 66370 73630 66390
rect 72782 66324 72790 66358
rect 72780 66310 72790 66324
rect 72710 66290 72790 66310
rect 72820 66314 73020 66320
rect 72820 66280 72832 66314
rect 73008 66310 73020 66314
rect 73318 66314 73518 66320
rect 73318 66310 73330 66314
rect 73008 66280 73330 66310
rect 73506 66280 73518 66314
rect 73550 66310 73560 66370
rect 73620 66310 73630 66370
rect 73550 66290 73630 66310
rect 72820 66274 73020 66280
rect 72600 66150 72670 66210
rect 72600 65910 72620 66150
rect 72660 65910 72670 66150
rect 73130 66270 73210 66280
rect 73318 66274 73518 66280
rect 73130 66210 73140 66270
rect 73200 66210 73210 66270
rect 73130 66160 73210 66210
rect 73130 66100 73140 66160
rect 73200 66100 73210 66160
rect 72820 66092 73020 66098
rect 72710 66060 72790 66080
rect 72710 66000 72720 66060
rect 72780 66048 72790 66060
rect 72820 66058 72832 66092
rect 73008 66090 73020 66092
rect 73130 66090 73210 66100
rect 73680 66230 73690 66470
rect 73730 66230 73750 66470
rect 73680 66150 73750 66230
rect 73318 66092 73518 66098
rect 73318 66090 73330 66092
rect 73008 66060 73330 66090
rect 73008 66058 73020 66060
rect 72820 66052 73020 66058
rect 73318 66058 73330 66060
rect 73506 66058 73518 66092
rect 73318 66052 73518 66058
rect 73550 66060 73630 66080
rect 72782 66014 72790 66048
rect 72780 66000 72790 66014
rect 72710 65980 72790 66000
rect 72820 66004 73020 66010
rect 72820 65970 72832 66004
rect 73008 66000 73020 66004
rect 73318 66004 73518 66010
rect 73318 66000 73330 66004
rect 73008 65990 73330 66000
rect 73008 65970 73140 65990
rect 72820 65964 73020 65970
rect 73130 65930 73140 65970
rect 73200 65970 73330 65990
rect 73506 65970 73518 66004
rect 73550 66000 73560 66060
rect 73620 66000 73630 66060
rect 73550 65980 73630 66000
rect 73200 65930 73210 65970
rect 73318 65964 73518 65970
rect 73130 65920 73210 65930
rect 72600 64760 72670 65910
rect 72600 64500 72620 64760
rect 72660 64500 72670 64760
rect 73680 65910 73690 66150
rect 73730 65910 73750 66150
rect 73680 64760 73750 65910
rect 73130 64730 73210 64740
rect 72820 64692 73020 64698
rect 72710 64660 72790 64680
rect 72710 64600 72720 64660
rect 72780 64648 72790 64660
rect 72820 64658 72832 64692
rect 73008 64690 73020 64692
rect 73130 64690 73140 64730
rect 73008 64670 73140 64690
rect 73200 64690 73210 64730
rect 73318 64692 73518 64698
rect 73318 64690 73330 64692
rect 73200 64670 73330 64690
rect 73008 64660 73330 64670
rect 73008 64658 73020 64660
rect 72820 64652 73020 64658
rect 73318 64658 73330 64660
rect 73506 64658 73518 64692
rect 73318 64652 73518 64658
rect 73550 64660 73630 64680
rect 72782 64614 72790 64648
rect 72780 64600 72790 64614
rect 72710 64580 72790 64600
rect 72820 64604 73020 64610
rect 72820 64570 72832 64604
rect 73008 64600 73020 64604
rect 73318 64604 73518 64610
rect 73318 64600 73330 64604
rect 73008 64570 73330 64600
rect 73506 64570 73518 64604
rect 73550 64600 73560 64660
rect 73620 64600 73630 64660
rect 73550 64580 73630 64600
rect 72820 64564 73020 64570
rect 72600 64440 72670 64500
rect 72600 64200 72620 64440
rect 72660 64200 72670 64440
rect 73130 64560 73210 64570
rect 73318 64564 73518 64570
rect 73130 64500 73140 64560
rect 73200 64500 73210 64560
rect 73130 64450 73210 64500
rect 73130 64390 73140 64450
rect 73200 64390 73210 64450
rect 72820 64382 73020 64388
rect 72710 64350 72790 64370
rect 72710 64290 72720 64350
rect 72780 64338 72790 64350
rect 72820 64348 72832 64382
rect 73008 64380 73020 64382
rect 73130 64380 73210 64390
rect 73680 64520 73690 64760
rect 73730 64520 73750 64760
rect 73680 64440 73750 64520
rect 73318 64382 73518 64388
rect 73318 64380 73330 64382
rect 73008 64350 73330 64380
rect 73008 64348 73020 64350
rect 72820 64342 73020 64348
rect 73318 64348 73330 64350
rect 73506 64348 73518 64382
rect 73318 64342 73518 64348
rect 73550 64350 73630 64370
rect 72782 64304 72790 64338
rect 72780 64290 72790 64304
rect 72710 64270 72790 64290
rect 72820 64294 73020 64300
rect 72820 64260 72832 64294
rect 73008 64290 73020 64294
rect 73318 64294 73518 64300
rect 73318 64290 73330 64294
rect 73008 64280 73330 64290
rect 73008 64260 73140 64280
rect 72820 64254 73020 64260
rect 73130 64220 73140 64260
rect 73200 64260 73330 64280
rect 73506 64260 73518 64294
rect 73550 64290 73560 64350
rect 73620 64290 73630 64350
rect 73550 64270 73630 64290
rect 73200 64220 73210 64260
rect 73318 64254 73518 64260
rect 73130 64210 73210 64220
rect 72600 63050 72670 64200
rect 72600 62790 72620 63050
rect 72660 62790 72670 63050
rect 73680 64200 73690 64440
rect 73730 64200 73750 64440
rect 73680 63050 73750 64200
rect 73130 63020 73210 63030
rect 72820 62982 73020 62988
rect 72710 62950 72790 62970
rect 72710 62890 72720 62950
rect 72780 62938 72790 62950
rect 72820 62948 72832 62982
rect 73008 62980 73020 62982
rect 73130 62980 73140 63020
rect 73008 62960 73140 62980
rect 73200 62980 73210 63020
rect 73318 62982 73518 62988
rect 73318 62980 73330 62982
rect 73200 62960 73330 62980
rect 73008 62950 73330 62960
rect 73008 62948 73020 62950
rect 72820 62942 73020 62948
rect 73318 62948 73330 62950
rect 73506 62948 73518 62982
rect 73318 62942 73518 62948
rect 73550 62950 73630 62970
rect 72782 62904 72790 62938
rect 72780 62890 72790 62904
rect 72710 62870 72790 62890
rect 72820 62894 73020 62900
rect 72820 62860 72832 62894
rect 73008 62890 73020 62894
rect 73318 62894 73518 62900
rect 73318 62890 73330 62894
rect 73008 62860 73330 62890
rect 73506 62860 73518 62894
rect 73550 62890 73560 62950
rect 73620 62890 73630 62950
rect 73550 62870 73630 62890
rect 72820 62854 73020 62860
rect 72600 62730 72670 62790
rect 72600 62490 72620 62730
rect 72660 62490 72670 62730
rect 73130 62850 73210 62860
rect 73318 62854 73518 62860
rect 73130 62790 73140 62850
rect 73200 62790 73210 62850
rect 73130 62740 73210 62790
rect 73130 62680 73140 62740
rect 73200 62680 73210 62740
rect 72820 62672 73020 62678
rect 72710 62640 72790 62660
rect 72710 62580 72720 62640
rect 72780 62628 72790 62640
rect 72820 62638 72832 62672
rect 73008 62670 73020 62672
rect 73130 62670 73210 62680
rect 73680 62810 73690 63050
rect 73730 62810 73750 63050
rect 73680 62730 73750 62810
rect 73318 62672 73518 62678
rect 73318 62670 73330 62672
rect 73008 62640 73330 62670
rect 73008 62638 73020 62640
rect 72820 62632 73020 62638
rect 73318 62638 73330 62640
rect 73506 62638 73518 62672
rect 73318 62632 73518 62638
rect 73550 62640 73630 62660
rect 72782 62594 72790 62628
rect 72780 62580 72790 62594
rect 72710 62560 72790 62580
rect 72820 62584 73020 62590
rect 72820 62550 72832 62584
rect 73008 62580 73020 62584
rect 73318 62584 73518 62590
rect 73318 62580 73330 62584
rect 73008 62570 73330 62580
rect 73008 62550 73140 62570
rect 72820 62544 73020 62550
rect 73130 62510 73140 62550
rect 73200 62550 73330 62570
rect 73506 62550 73518 62584
rect 73550 62580 73560 62640
rect 73620 62580 73630 62640
rect 73550 62560 73630 62580
rect 73200 62510 73210 62550
rect 73318 62544 73518 62550
rect 73130 62500 73210 62510
rect 72600 61340 72670 62490
rect 72600 61080 72620 61340
rect 72660 61080 72670 61340
rect 73680 62490 73690 62730
rect 73730 62490 73750 62730
rect 73680 61340 73750 62490
rect 73130 61310 73210 61320
rect 72820 61272 73020 61278
rect 72710 61240 72790 61260
rect 72710 61180 72720 61240
rect 72780 61228 72790 61240
rect 72820 61238 72832 61272
rect 73008 61270 73020 61272
rect 73130 61270 73140 61310
rect 73008 61250 73140 61270
rect 73200 61270 73210 61310
rect 73318 61272 73518 61278
rect 73318 61270 73330 61272
rect 73200 61250 73330 61270
rect 73008 61240 73330 61250
rect 73008 61238 73020 61240
rect 72820 61232 73020 61238
rect 73318 61238 73330 61240
rect 73506 61238 73518 61272
rect 73318 61232 73518 61238
rect 73550 61240 73630 61260
rect 72782 61194 72790 61228
rect 72780 61180 72790 61194
rect 72710 61160 72790 61180
rect 72820 61184 73020 61190
rect 72820 61150 72832 61184
rect 73008 61180 73020 61184
rect 73318 61184 73518 61190
rect 73318 61180 73330 61184
rect 73008 61150 73330 61180
rect 73506 61150 73518 61184
rect 73550 61180 73560 61240
rect 73620 61180 73630 61240
rect 73550 61160 73630 61180
rect 72820 61144 73020 61150
rect 72600 61020 72670 61080
rect 72600 60780 72620 61020
rect 72660 60780 72670 61020
rect 73130 61140 73210 61150
rect 73318 61144 73518 61150
rect 73130 61080 73140 61140
rect 73200 61080 73210 61140
rect 73130 61030 73210 61080
rect 73130 60970 73140 61030
rect 73200 60970 73210 61030
rect 72820 60962 73020 60968
rect 72710 60930 72790 60950
rect 72710 60870 72720 60930
rect 72780 60918 72790 60930
rect 72820 60928 72832 60962
rect 73008 60960 73020 60962
rect 73130 60960 73210 60970
rect 73680 61100 73690 61340
rect 73730 61100 73750 61340
rect 73680 61020 73750 61100
rect 73318 60962 73518 60968
rect 73318 60960 73330 60962
rect 73008 60930 73330 60960
rect 73008 60928 73020 60930
rect 72820 60922 73020 60928
rect 73318 60928 73330 60930
rect 73506 60928 73518 60962
rect 73318 60922 73518 60928
rect 73550 60930 73630 60950
rect 72782 60884 72790 60918
rect 72780 60870 72790 60884
rect 72710 60850 72790 60870
rect 72820 60874 73020 60880
rect 72820 60840 72832 60874
rect 73008 60870 73020 60874
rect 73318 60874 73518 60880
rect 73318 60870 73330 60874
rect 73008 60860 73330 60870
rect 73008 60840 73140 60860
rect 72820 60834 73020 60840
rect 73130 60800 73140 60840
rect 73200 60840 73330 60860
rect 73506 60840 73518 60874
rect 73550 60870 73560 60930
rect 73620 60870 73630 60930
rect 73550 60850 73630 60870
rect 73200 60800 73210 60840
rect 73318 60834 73518 60840
rect 73130 60790 73210 60800
rect 72600 59630 72670 60780
rect 72600 59370 72620 59630
rect 72660 59370 72670 59630
rect 73680 60780 73690 61020
rect 73730 60780 73750 61020
rect 73680 59630 73750 60780
rect 73130 59600 73210 59610
rect 72820 59562 73020 59568
rect 72710 59530 72790 59550
rect 72710 59470 72720 59530
rect 72780 59518 72790 59530
rect 72820 59528 72832 59562
rect 73008 59560 73020 59562
rect 73130 59560 73140 59600
rect 73008 59540 73140 59560
rect 73200 59560 73210 59600
rect 73318 59562 73518 59568
rect 73318 59560 73330 59562
rect 73200 59540 73330 59560
rect 73008 59530 73330 59540
rect 73008 59528 73020 59530
rect 72820 59522 73020 59528
rect 73318 59528 73330 59530
rect 73506 59528 73518 59562
rect 73318 59522 73518 59528
rect 73550 59530 73630 59550
rect 72782 59484 72790 59518
rect 72780 59470 72790 59484
rect 72710 59450 72790 59470
rect 72820 59474 73020 59480
rect 72820 59440 72832 59474
rect 73008 59470 73020 59474
rect 73318 59474 73518 59480
rect 73318 59470 73330 59474
rect 73008 59440 73330 59470
rect 73506 59440 73518 59474
rect 73550 59470 73560 59530
rect 73620 59470 73630 59530
rect 73550 59450 73630 59470
rect 72820 59434 73020 59440
rect 72600 59310 72670 59370
rect 72600 59070 72620 59310
rect 72660 59070 72670 59310
rect 73130 59430 73210 59440
rect 73318 59434 73518 59440
rect 73130 59370 73140 59430
rect 73200 59370 73210 59430
rect 73130 59320 73210 59370
rect 73130 59260 73140 59320
rect 73200 59260 73210 59320
rect 72820 59252 73020 59258
rect 72710 59220 72790 59240
rect 72710 59160 72720 59220
rect 72780 59208 72790 59220
rect 72820 59218 72832 59252
rect 73008 59250 73020 59252
rect 73130 59250 73210 59260
rect 73680 59390 73690 59630
rect 73730 59390 73750 59630
rect 73680 59310 73750 59390
rect 73318 59252 73518 59258
rect 73318 59250 73330 59252
rect 73008 59220 73330 59250
rect 73008 59218 73020 59220
rect 72820 59212 73020 59218
rect 73318 59218 73330 59220
rect 73506 59218 73518 59252
rect 73318 59212 73518 59218
rect 73550 59220 73630 59240
rect 72782 59174 72790 59208
rect 72780 59160 72790 59174
rect 72710 59140 72790 59160
rect 72820 59164 73020 59170
rect 72820 59130 72832 59164
rect 73008 59160 73020 59164
rect 73318 59164 73518 59170
rect 73318 59160 73330 59164
rect 73008 59150 73330 59160
rect 73008 59130 73140 59150
rect 72820 59124 73020 59130
rect 73130 59090 73140 59130
rect 73200 59130 73330 59150
rect 73506 59130 73518 59164
rect 73550 59160 73560 59220
rect 73620 59160 73630 59220
rect 73550 59140 73630 59160
rect 73200 59090 73210 59130
rect 73318 59124 73518 59130
rect 73130 59080 73210 59090
rect 72600 57920 72670 59070
rect 72600 57660 72620 57920
rect 72660 57660 72670 57920
rect 73680 59070 73690 59310
rect 73730 59070 73750 59310
rect 73680 57920 73750 59070
rect 73130 57890 73210 57900
rect 72820 57852 73020 57858
rect 72710 57820 72790 57840
rect 72710 57760 72720 57820
rect 72780 57808 72790 57820
rect 72820 57818 72832 57852
rect 73008 57850 73020 57852
rect 73130 57850 73140 57890
rect 73008 57830 73140 57850
rect 73200 57850 73210 57890
rect 73318 57852 73518 57858
rect 73318 57850 73330 57852
rect 73200 57830 73330 57850
rect 73008 57820 73330 57830
rect 73008 57818 73020 57820
rect 72820 57812 73020 57818
rect 73318 57818 73330 57820
rect 73506 57818 73518 57852
rect 73318 57812 73518 57818
rect 73550 57820 73630 57840
rect 72782 57774 72790 57808
rect 72780 57760 72790 57774
rect 72710 57740 72790 57760
rect 72820 57764 73020 57770
rect 72820 57730 72832 57764
rect 73008 57760 73020 57764
rect 73318 57764 73518 57770
rect 73318 57760 73330 57764
rect 73008 57730 73330 57760
rect 73506 57730 73518 57764
rect 73550 57760 73560 57820
rect 73620 57760 73630 57820
rect 73550 57740 73630 57760
rect 72820 57724 73020 57730
rect 72600 57600 72670 57660
rect 72600 57360 72620 57600
rect 72660 57360 72670 57600
rect 73130 57720 73210 57730
rect 73318 57724 73518 57730
rect 73130 57660 73140 57720
rect 73200 57660 73210 57720
rect 73130 57610 73210 57660
rect 73130 57550 73140 57610
rect 73200 57550 73210 57610
rect 72820 57542 73020 57548
rect 72710 57510 72790 57530
rect 72710 57450 72720 57510
rect 72780 57498 72790 57510
rect 72820 57508 72832 57542
rect 73008 57540 73020 57542
rect 73130 57540 73210 57550
rect 73680 57680 73690 57920
rect 73730 57680 73750 57920
rect 73680 57600 73750 57680
rect 73318 57542 73518 57548
rect 73318 57540 73330 57542
rect 73008 57510 73330 57540
rect 73008 57508 73020 57510
rect 72820 57502 73020 57508
rect 73318 57508 73330 57510
rect 73506 57508 73518 57542
rect 73318 57502 73518 57508
rect 73550 57510 73630 57530
rect 72782 57464 72790 57498
rect 72780 57450 72790 57464
rect 72710 57430 72790 57450
rect 72820 57454 73020 57460
rect 72820 57420 72832 57454
rect 73008 57450 73020 57454
rect 73318 57454 73518 57460
rect 73318 57450 73330 57454
rect 73008 57440 73330 57450
rect 73008 57420 73140 57440
rect 72820 57414 73020 57420
rect 73130 57380 73140 57420
rect 73200 57420 73330 57440
rect 73506 57420 73518 57454
rect 73550 57450 73560 57510
rect 73620 57450 73630 57510
rect 73550 57430 73630 57450
rect 73200 57380 73210 57420
rect 73318 57414 73518 57420
rect 73130 57370 73210 57380
rect 72600 56210 72670 57360
rect 72600 55950 72620 56210
rect 72660 55950 72670 56210
rect 73680 57360 73690 57600
rect 73730 57360 73750 57600
rect 73680 56210 73750 57360
rect 73130 56180 73210 56190
rect 72820 56142 73020 56148
rect 72710 56110 72790 56130
rect 72710 56050 72720 56110
rect 72780 56098 72790 56110
rect 72820 56108 72832 56142
rect 73008 56140 73020 56142
rect 73130 56140 73140 56180
rect 73008 56120 73140 56140
rect 73200 56140 73210 56180
rect 73318 56142 73518 56148
rect 73318 56140 73330 56142
rect 73200 56120 73330 56140
rect 73008 56110 73330 56120
rect 73008 56108 73020 56110
rect 72820 56102 73020 56108
rect 73318 56108 73330 56110
rect 73506 56108 73518 56142
rect 73318 56102 73518 56108
rect 73550 56110 73630 56130
rect 72782 56064 72790 56098
rect 72780 56050 72790 56064
rect 72710 56030 72790 56050
rect 72820 56054 73020 56060
rect 72820 56020 72832 56054
rect 73008 56050 73020 56054
rect 73318 56054 73518 56060
rect 73318 56050 73330 56054
rect 73008 56020 73330 56050
rect 73506 56020 73518 56054
rect 73550 56050 73560 56110
rect 73620 56050 73630 56110
rect 73550 56030 73630 56050
rect 72820 56014 73020 56020
rect 72600 55890 72670 55950
rect 72600 55650 72620 55890
rect 72660 55650 72670 55890
rect 73130 56010 73210 56020
rect 73318 56014 73518 56020
rect 73130 55950 73140 56010
rect 73200 55950 73210 56010
rect 73130 55900 73210 55950
rect 73130 55840 73140 55900
rect 73200 55840 73210 55900
rect 72820 55832 73020 55838
rect 72710 55800 72790 55820
rect 72710 55740 72720 55800
rect 72780 55788 72790 55800
rect 72820 55798 72832 55832
rect 73008 55830 73020 55832
rect 73130 55830 73210 55840
rect 73680 55970 73690 56210
rect 73730 55970 73750 56210
rect 73680 55890 73750 55970
rect 73318 55832 73518 55838
rect 73318 55830 73330 55832
rect 73008 55800 73330 55830
rect 73008 55798 73020 55800
rect 72820 55792 73020 55798
rect 73318 55798 73330 55800
rect 73506 55798 73518 55832
rect 73318 55792 73518 55798
rect 73550 55800 73630 55820
rect 72782 55754 72790 55788
rect 72780 55740 72790 55754
rect 72710 55720 72790 55740
rect 72820 55744 73020 55750
rect 72820 55710 72832 55744
rect 73008 55740 73020 55744
rect 73318 55744 73518 55750
rect 73318 55740 73330 55744
rect 73008 55730 73330 55740
rect 73008 55710 73140 55730
rect 72820 55704 73020 55710
rect 73130 55670 73140 55710
rect 73200 55710 73330 55730
rect 73506 55710 73518 55744
rect 73550 55740 73560 55800
rect 73620 55740 73630 55800
rect 73550 55720 73630 55740
rect 73200 55670 73210 55710
rect 73318 55704 73518 55710
rect 73130 55660 73210 55670
rect 72600 54500 72670 55650
rect 72600 54240 72620 54500
rect 72660 54240 72670 54500
rect 73680 55650 73690 55890
rect 73730 55650 73750 55890
rect 73680 54500 73750 55650
rect 73130 54470 73210 54480
rect 72820 54432 73020 54438
rect 72710 54400 72790 54420
rect 72710 54340 72720 54400
rect 72780 54388 72790 54400
rect 72820 54398 72832 54432
rect 73008 54430 73020 54432
rect 73130 54430 73140 54470
rect 73008 54410 73140 54430
rect 73200 54430 73210 54470
rect 73318 54432 73518 54438
rect 73318 54430 73330 54432
rect 73200 54410 73330 54430
rect 73008 54400 73330 54410
rect 73008 54398 73020 54400
rect 72820 54392 73020 54398
rect 73318 54398 73330 54400
rect 73506 54398 73518 54432
rect 73318 54392 73518 54398
rect 73550 54400 73630 54420
rect 72782 54354 72790 54388
rect 72780 54340 72790 54354
rect 72710 54320 72790 54340
rect 72820 54344 73020 54350
rect 72820 54310 72832 54344
rect 73008 54340 73020 54344
rect 73318 54344 73518 54350
rect 73318 54340 73330 54344
rect 73008 54310 73330 54340
rect 73506 54310 73518 54344
rect 73550 54340 73560 54400
rect 73620 54340 73630 54400
rect 73550 54320 73630 54340
rect 72820 54304 73020 54310
rect 72600 54180 72670 54240
rect 72600 53940 72620 54180
rect 72660 53940 72670 54180
rect 73130 54300 73210 54310
rect 73318 54304 73518 54310
rect 73130 54240 73140 54300
rect 73200 54240 73210 54300
rect 73130 54190 73210 54240
rect 73130 54130 73140 54190
rect 73200 54130 73210 54190
rect 72820 54122 73020 54128
rect 72710 54090 72790 54110
rect 72710 54030 72720 54090
rect 72780 54078 72790 54090
rect 72820 54088 72832 54122
rect 73008 54120 73020 54122
rect 73130 54120 73210 54130
rect 73680 54260 73690 54500
rect 73730 54260 73750 54500
rect 73680 54180 73750 54260
rect 73318 54122 73518 54128
rect 73318 54120 73330 54122
rect 73008 54090 73330 54120
rect 73008 54088 73020 54090
rect 72820 54082 73020 54088
rect 73318 54088 73330 54090
rect 73506 54088 73518 54122
rect 73318 54082 73518 54088
rect 73550 54090 73630 54110
rect 72782 54044 72790 54078
rect 72780 54030 72790 54044
rect 72710 54010 72790 54030
rect 72820 54034 73020 54040
rect 72820 54000 72832 54034
rect 73008 54030 73020 54034
rect 73318 54034 73518 54040
rect 73318 54030 73330 54034
rect 73008 54020 73330 54030
rect 73008 54000 73140 54020
rect 72820 53994 73020 54000
rect 73130 53960 73140 54000
rect 73200 54000 73330 54020
rect 73506 54000 73518 54034
rect 73550 54030 73560 54090
rect 73620 54030 73630 54090
rect 73550 54010 73630 54030
rect 73200 53960 73210 54000
rect 73318 53994 73518 54000
rect 73130 53950 73210 53960
rect 72600 52790 72670 53940
rect 72600 52530 72620 52790
rect 72660 52530 72670 52790
rect 73680 53940 73690 54180
rect 73730 53940 73750 54180
rect 73680 52790 73750 53940
rect 73130 52760 73210 52770
rect 72820 52722 73020 52728
rect 72710 52690 72790 52710
rect 72710 52630 72720 52690
rect 72780 52678 72790 52690
rect 72820 52688 72832 52722
rect 73008 52720 73020 52722
rect 73130 52720 73140 52760
rect 73008 52700 73140 52720
rect 73200 52720 73210 52760
rect 73318 52722 73518 52728
rect 73318 52720 73330 52722
rect 73200 52700 73330 52720
rect 73008 52690 73330 52700
rect 73008 52688 73020 52690
rect 72820 52682 73020 52688
rect 73318 52688 73330 52690
rect 73506 52688 73518 52722
rect 73318 52682 73518 52688
rect 73550 52690 73630 52710
rect 72782 52644 72790 52678
rect 72780 52630 72790 52644
rect 72710 52610 72790 52630
rect 72820 52634 73020 52640
rect 72820 52600 72832 52634
rect 73008 52630 73020 52634
rect 73318 52634 73518 52640
rect 73318 52630 73330 52634
rect 73008 52600 73330 52630
rect 73506 52600 73518 52634
rect 73550 52630 73560 52690
rect 73620 52630 73630 52690
rect 73550 52610 73630 52630
rect 72820 52594 73020 52600
rect 72600 52470 72670 52530
rect 72600 52230 72620 52470
rect 72660 52230 72670 52470
rect 73130 52590 73210 52600
rect 73318 52594 73518 52600
rect 73130 52530 73140 52590
rect 73200 52530 73210 52590
rect 73130 52480 73210 52530
rect 73130 52420 73140 52480
rect 73200 52420 73210 52480
rect 72820 52412 73020 52418
rect 72710 52380 72790 52400
rect 72710 52320 72720 52380
rect 72780 52368 72790 52380
rect 72820 52378 72832 52412
rect 73008 52410 73020 52412
rect 73130 52410 73210 52420
rect 73680 52550 73690 52790
rect 73730 52550 73750 52790
rect 73680 52470 73750 52550
rect 73318 52412 73518 52418
rect 73318 52410 73330 52412
rect 73008 52380 73330 52410
rect 73008 52378 73020 52380
rect 72820 52372 73020 52378
rect 73318 52378 73330 52380
rect 73506 52378 73518 52412
rect 73318 52372 73518 52378
rect 73550 52380 73630 52400
rect 72782 52334 72790 52368
rect 72780 52320 72790 52334
rect 72710 52300 72790 52320
rect 72820 52324 73020 52330
rect 72820 52290 72832 52324
rect 73008 52320 73020 52324
rect 73318 52324 73518 52330
rect 73318 52320 73330 52324
rect 73008 52310 73330 52320
rect 73008 52290 73140 52310
rect 72820 52284 73020 52290
rect 73130 52250 73140 52290
rect 73200 52290 73330 52310
rect 73506 52290 73518 52324
rect 73550 52320 73560 52380
rect 73620 52320 73630 52380
rect 73550 52300 73630 52320
rect 73200 52250 73210 52290
rect 73318 52284 73518 52290
rect 73130 52240 73210 52250
rect 72600 51080 72670 52230
rect 72600 50820 72620 51080
rect 72660 50820 72670 51080
rect 73680 52230 73690 52470
rect 73730 52230 73750 52470
rect 73680 51080 73750 52230
rect 73130 51050 73210 51060
rect 72820 51012 73020 51018
rect 72710 50980 72790 51000
rect 72710 50920 72720 50980
rect 72780 50968 72790 50980
rect 72820 50978 72832 51012
rect 73008 51010 73020 51012
rect 73130 51010 73140 51050
rect 73008 50990 73140 51010
rect 73200 51010 73210 51050
rect 73318 51012 73518 51018
rect 73318 51010 73330 51012
rect 73200 50990 73330 51010
rect 73008 50980 73330 50990
rect 73008 50978 73020 50980
rect 72820 50972 73020 50978
rect 73318 50978 73330 50980
rect 73506 50978 73518 51012
rect 73318 50972 73518 50978
rect 73550 50980 73630 51000
rect 72782 50934 72790 50968
rect 72780 50920 72790 50934
rect 72710 50900 72790 50920
rect 72820 50924 73020 50930
rect 72820 50890 72832 50924
rect 73008 50920 73020 50924
rect 73318 50924 73518 50930
rect 73318 50920 73330 50924
rect 73008 50890 73330 50920
rect 73506 50890 73518 50924
rect 73550 50920 73560 50980
rect 73620 50920 73630 50980
rect 73550 50900 73630 50920
rect 72820 50884 73020 50890
rect 72600 50760 72670 50820
rect 72600 50520 72620 50760
rect 72660 50520 72670 50760
rect 73130 50880 73210 50890
rect 73318 50884 73518 50890
rect 73130 50820 73140 50880
rect 73200 50820 73210 50880
rect 73130 50770 73210 50820
rect 73130 50710 73140 50770
rect 73200 50710 73210 50770
rect 72820 50702 73020 50708
rect 72710 50670 72790 50690
rect 72710 50610 72720 50670
rect 72780 50658 72790 50670
rect 72820 50668 72832 50702
rect 73008 50700 73020 50702
rect 73130 50700 73210 50710
rect 73680 50840 73690 51080
rect 73730 50840 73750 51080
rect 73680 50760 73750 50840
rect 73318 50702 73518 50708
rect 73318 50700 73330 50702
rect 73008 50670 73330 50700
rect 73008 50668 73020 50670
rect 72820 50662 73020 50668
rect 73318 50668 73330 50670
rect 73506 50668 73518 50702
rect 73318 50662 73518 50668
rect 73550 50670 73630 50690
rect 72782 50624 72790 50658
rect 72780 50610 72790 50624
rect 72710 50590 72790 50610
rect 72820 50614 73020 50620
rect 72820 50580 72832 50614
rect 73008 50610 73020 50614
rect 73318 50614 73518 50620
rect 73318 50610 73330 50614
rect 73008 50600 73330 50610
rect 73008 50580 73140 50600
rect 72820 50574 73020 50580
rect 73130 50540 73140 50580
rect 73200 50580 73330 50600
rect 73506 50580 73518 50614
rect 73550 50610 73560 50670
rect 73620 50610 73630 50670
rect 73550 50590 73630 50610
rect 73200 50540 73210 50580
rect 73318 50574 73518 50580
rect 73130 50530 73210 50540
rect 72600 49370 72670 50520
rect 72600 49110 72620 49370
rect 72660 49110 72670 49370
rect 73680 50520 73690 50760
rect 73730 50520 73750 50760
rect 73680 49370 73750 50520
rect 73130 49340 73210 49350
rect 72820 49302 73020 49308
rect 72710 49270 72790 49290
rect 72710 49210 72720 49270
rect 72780 49258 72790 49270
rect 72820 49268 72832 49302
rect 73008 49300 73020 49302
rect 73130 49300 73140 49340
rect 73008 49280 73140 49300
rect 73200 49300 73210 49340
rect 73318 49302 73518 49308
rect 73318 49300 73330 49302
rect 73200 49280 73330 49300
rect 73008 49270 73330 49280
rect 73008 49268 73020 49270
rect 72820 49262 73020 49268
rect 73318 49268 73330 49270
rect 73506 49268 73518 49302
rect 73318 49262 73518 49268
rect 73550 49270 73630 49290
rect 72782 49224 72790 49258
rect 72780 49210 72790 49224
rect 72710 49190 72790 49210
rect 72820 49214 73020 49220
rect 72820 49180 72832 49214
rect 73008 49210 73020 49214
rect 73318 49214 73518 49220
rect 73318 49210 73330 49214
rect 73008 49180 73330 49210
rect 73506 49180 73518 49214
rect 73550 49210 73560 49270
rect 73620 49210 73630 49270
rect 73550 49190 73630 49210
rect 72820 49174 73020 49180
rect 72600 49050 72670 49110
rect 72600 48810 72620 49050
rect 72660 48810 72670 49050
rect 73130 49170 73210 49180
rect 73318 49174 73518 49180
rect 73130 49110 73140 49170
rect 73200 49110 73210 49170
rect 73130 49060 73210 49110
rect 73130 49000 73140 49060
rect 73200 49000 73210 49060
rect 72820 48992 73020 48998
rect 72710 48960 72790 48980
rect 72710 48900 72720 48960
rect 72780 48948 72790 48960
rect 72820 48958 72832 48992
rect 73008 48990 73020 48992
rect 73130 48990 73210 49000
rect 73680 49130 73690 49370
rect 73730 49130 73750 49370
rect 73680 49050 73750 49130
rect 73318 48992 73518 48998
rect 73318 48990 73330 48992
rect 73008 48960 73330 48990
rect 73008 48958 73020 48960
rect 72820 48952 73020 48958
rect 73318 48958 73330 48960
rect 73506 48958 73518 48992
rect 73318 48952 73518 48958
rect 73550 48960 73630 48980
rect 72782 48914 72790 48948
rect 72780 48900 72790 48914
rect 72710 48880 72790 48900
rect 72820 48904 73020 48910
rect 72820 48870 72832 48904
rect 73008 48900 73020 48904
rect 73318 48904 73518 48910
rect 73318 48900 73330 48904
rect 73008 48890 73330 48900
rect 73008 48870 73140 48890
rect 72820 48864 73020 48870
rect 73130 48830 73140 48870
rect 73200 48870 73330 48890
rect 73506 48870 73518 48904
rect 73550 48900 73560 48960
rect 73620 48900 73630 48960
rect 73550 48880 73630 48900
rect 73200 48830 73210 48870
rect 73318 48864 73518 48870
rect 73130 48820 73210 48830
rect 72600 47660 72670 48810
rect 72600 47400 72620 47660
rect 72660 47400 72670 47660
rect 73680 48810 73690 49050
rect 73730 48810 73750 49050
rect 73680 47660 73750 48810
rect 73130 47630 73210 47640
rect 72820 47592 73020 47598
rect 72710 47560 72790 47580
rect 72710 47500 72720 47560
rect 72780 47548 72790 47560
rect 72820 47558 72832 47592
rect 73008 47590 73020 47592
rect 73130 47590 73140 47630
rect 73008 47570 73140 47590
rect 73200 47590 73210 47630
rect 73318 47592 73518 47598
rect 73318 47590 73330 47592
rect 73200 47570 73330 47590
rect 73008 47560 73330 47570
rect 73008 47558 73020 47560
rect 72820 47552 73020 47558
rect 73318 47558 73330 47560
rect 73506 47558 73518 47592
rect 73318 47552 73518 47558
rect 73550 47560 73630 47580
rect 72782 47514 72790 47548
rect 72780 47500 72790 47514
rect 72710 47480 72790 47500
rect 72820 47504 73020 47510
rect 72820 47470 72832 47504
rect 73008 47500 73020 47504
rect 73318 47504 73518 47510
rect 73318 47500 73330 47504
rect 73008 47470 73330 47500
rect 73506 47470 73518 47504
rect 73550 47500 73560 47560
rect 73620 47500 73630 47560
rect 73550 47480 73630 47500
rect 72820 47464 73020 47470
rect 72600 47340 72670 47400
rect 72600 47100 72620 47340
rect 72660 47100 72670 47340
rect 73130 47460 73210 47470
rect 73318 47464 73518 47470
rect 73130 47400 73140 47460
rect 73200 47400 73210 47460
rect 73130 47350 73210 47400
rect 73130 47290 73140 47350
rect 73200 47290 73210 47350
rect 72820 47282 73020 47288
rect 72710 47250 72790 47270
rect 72710 47190 72720 47250
rect 72780 47238 72790 47250
rect 72820 47248 72832 47282
rect 73008 47280 73020 47282
rect 73130 47280 73210 47290
rect 73680 47420 73690 47660
rect 73730 47420 73750 47660
rect 73680 47340 73750 47420
rect 73318 47282 73518 47288
rect 73318 47280 73330 47282
rect 73008 47250 73330 47280
rect 73008 47248 73020 47250
rect 72820 47242 73020 47248
rect 73318 47248 73330 47250
rect 73506 47248 73518 47282
rect 73318 47242 73518 47248
rect 73550 47250 73630 47270
rect 72782 47204 72790 47238
rect 72780 47190 72790 47204
rect 72710 47170 72790 47190
rect 72820 47194 73020 47200
rect 72820 47160 72832 47194
rect 73008 47190 73020 47194
rect 73318 47194 73518 47200
rect 73318 47190 73330 47194
rect 73008 47180 73330 47190
rect 73008 47160 73140 47180
rect 72820 47154 73020 47160
rect 73130 47120 73140 47160
rect 73200 47160 73330 47180
rect 73506 47160 73518 47194
rect 73550 47190 73560 47250
rect 73620 47190 73630 47250
rect 73550 47170 73630 47190
rect 73200 47120 73210 47160
rect 73318 47154 73518 47160
rect 73130 47110 73210 47120
rect 72600 45950 72670 47100
rect 72600 45690 72620 45950
rect 72660 45690 72670 45950
rect 73680 47100 73690 47340
rect 73730 47100 73750 47340
rect 73680 45950 73750 47100
rect 73130 45920 73210 45930
rect 72820 45882 73020 45888
rect 72710 45850 72790 45870
rect 72710 45790 72720 45850
rect 72780 45838 72790 45850
rect 72820 45848 72832 45882
rect 73008 45880 73020 45882
rect 73130 45880 73140 45920
rect 73008 45860 73140 45880
rect 73200 45880 73210 45920
rect 73318 45882 73518 45888
rect 73318 45880 73330 45882
rect 73200 45860 73330 45880
rect 73008 45850 73330 45860
rect 73008 45848 73020 45850
rect 72820 45842 73020 45848
rect 73318 45848 73330 45850
rect 73506 45848 73518 45882
rect 73318 45842 73518 45848
rect 73550 45850 73630 45870
rect 72782 45804 72790 45838
rect 72780 45790 72790 45804
rect 72710 45770 72790 45790
rect 72820 45794 73020 45800
rect 72820 45760 72832 45794
rect 73008 45790 73020 45794
rect 73318 45794 73518 45800
rect 73318 45790 73330 45794
rect 73008 45760 73330 45790
rect 73506 45760 73518 45794
rect 73550 45790 73560 45850
rect 73620 45790 73630 45850
rect 73550 45770 73630 45790
rect 72820 45754 73020 45760
rect 72600 45630 72670 45690
rect 72600 45390 72620 45630
rect 72660 45390 72670 45630
rect 73130 45750 73210 45760
rect 73318 45754 73518 45760
rect 73130 45690 73140 45750
rect 73200 45690 73210 45750
rect 73130 45640 73210 45690
rect 73130 45580 73140 45640
rect 73200 45580 73210 45640
rect 72820 45572 73020 45578
rect 72710 45540 72790 45560
rect 72710 45480 72720 45540
rect 72780 45528 72790 45540
rect 72820 45538 72832 45572
rect 73008 45570 73020 45572
rect 73130 45570 73210 45580
rect 73680 45710 73690 45950
rect 73730 45710 73750 45950
rect 73680 45630 73750 45710
rect 73318 45572 73518 45578
rect 73318 45570 73330 45572
rect 73008 45540 73330 45570
rect 73008 45538 73020 45540
rect 72820 45532 73020 45538
rect 73318 45538 73330 45540
rect 73506 45538 73518 45572
rect 73318 45532 73518 45538
rect 73550 45540 73630 45560
rect 72782 45494 72790 45528
rect 72780 45480 72790 45494
rect 72710 45460 72790 45480
rect 72820 45484 73020 45490
rect 72820 45450 72832 45484
rect 73008 45480 73020 45484
rect 73318 45484 73518 45490
rect 73318 45480 73330 45484
rect 73008 45470 73330 45480
rect 73008 45450 73140 45470
rect 72820 45444 73020 45450
rect 73130 45410 73140 45450
rect 73200 45450 73330 45470
rect 73506 45450 73518 45484
rect 73550 45480 73560 45540
rect 73620 45480 73630 45540
rect 73550 45460 73630 45480
rect 73200 45410 73210 45450
rect 73318 45444 73518 45450
rect 73130 45400 73210 45410
rect 72600 44240 72670 45390
rect 72600 43980 72620 44240
rect 72660 43980 72670 44240
rect 73680 45390 73690 45630
rect 73730 45390 73750 45630
rect 73680 44240 73750 45390
rect 73130 44210 73210 44220
rect 72820 44172 73020 44178
rect 72710 44140 72790 44160
rect 72710 44080 72720 44140
rect 72780 44128 72790 44140
rect 72820 44138 72832 44172
rect 73008 44170 73020 44172
rect 73130 44170 73140 44210
rect 73008 44150 73140 44170
rect 73200 44170 73210 44210
rect 73318 44172 73518 44178
rect 73318 44170 73330 44172
rect 73200 44150 73330 44170
rect 73008 44140 73330 44150
rect 73008 44138 73020 44140
rect 72820 44132 73020 44138
rect 73318 44138 73330 44140
rect 73506 44138 73518 44172
rect 73318 44132 73518 44138
rect 73550 44140 73630 44160
rect 72782 44094 72790 44128
rect 72780 44080 72790 44094
rect 72710 44060 72790 44080
rect 72820 44084 73020 44090
rect 72820 44050 72832 44084
rect 73008 44080 73020 44084
rect 73318 44084 73518 44090
rect 73318 44080 73330 44084
rect 73008 44050 73330 44080
rect 73506 44050 73518 44084
rect 73550 44080 73560 44140
rect 73620 44080 73630 44140
rect 73550 44060 73630 44080
rect 72820 44044 73020 44050
rect 72600 43920 72670 43980
rect 72600 43680 72620 43920
rect 72660 43680 72670 43920
rect 73130 44040 73210 44050
rect 73318 44044 73518 44050
rect 73130 43980 73140 44040
rect 73200 43980 73210 44040
rect 73130 43930 73210 43980
rect 73130 43870 73140 43930
rect 73200 43870 73210 43930
rect 72820 43862 73020 43868
rect 72710 43830 72790 43850
rect 72710 43770 72720 43830
rect 72780 43818 72790 43830
rect 72820 43828 72832 43862
rect 73008 43860 73020 43862
rect 73130 43860 73210 43870
rect 73680 44000 73690 44240
rect 73730 44000 73750 44240
rect 73680 43920 73750 44000
rect 73318 43862 73518 43868
rect 73318 43860 73330 43862
rect 73008 43830 73330 43860
rect 73008 43828 73020 43830
rect 72820 43822 73020 43828
rect 73318 43828 73330 43830
rect 73506 43828 73518 43862
rect 73318 43822 73518 43828
rect 73550 43830 73630 43850
rect 72782 43784 72790 43818
rect 72780 43770 72790 43784
rect 72710 43750 72790 43770
rect 72820 43774 73020 43780
rect 72820 43740 72832 43774
rect 73008 43770 73020 43774
rect 73318 43774 73518 43780
rect 73318 43770 73330 43774
rect 73008 43760 73330 43770
rect 73008 43740 73140 43760
rect 72820 43734 73020 43740
rect 73130 43700 73140 43740
rect 73200 43740 73330 43760
rect 73506 43740 73518 43774
rect 73550 43770 73560 43830
rect 73620 43770 73630 43830
rect 73550 43750 73630 43770
rect 73200 43700 73210 43740
rect 73318 43734 73518 43740
rect 73130 43690 73210 43700
rect 72600 42530 72670 43680
rect 72600 42270 72620 42530
rect 72660 42270 72670 42530
rect 73680 43680 73690 43920
rect 73730 43680 73750 43920
rect 73680 42530 73750 43680
rect 73130 42500 73210 42510
rect 72820 42462 73020 42468
rect 72710 42430 72790 42450
rect 72710 42370 72720 42430
rect 72780 42418 72790 42430
rect 72820 42428 72832 42462
rect 73008 42460 73020 42462
rect 73130 42460 73140 42500
rect 73008 42440 73140 42460
rect 73200 42460 73210 42500
rect 73318 42462 73518 42468
rect 73318 42460 73330 42462
rect 73200 42440 73330 42460
rect 73008 42430 73330 42440
rect 73008 42428 73020 42430
rect 72820 42422 73020 42428
rect 73318 42428 73330 42430
rect 73506 42428 73518 42462
rect 73318 42422 73518 42428
rect 73550 42430 73630 42450
rect 72782 42384 72790 42418
rect 72780 42370 72790 42384
rect 72710 42350 72790 42370
rect 72820 42374 73020 42380
rect 72820 42340 72832 42374
rect 73008 42370 73020 42374
rect 73318 42374 73518 42380
rect 73318 42370 73330 42374
rect 73008 42340 73330 42370
rect 73506 42340 73518 42374
rect 73550 42370 73560 42430
rect 73620 42370 73630 42430
rect 73550 42350 73630 42370
rect 72820 42334 73020 42340
rect 72600 42210 72670 42270
rect 72600 41970 72620 42210
rect 72660 41970 72670 42210
rect 73130 42330 73210 42340
rect 73318 42334 73518 42340
rect 73130 42270 73140 42330
rect 73200 42270 73210 42330
rect 73130 42220 73210 42270
rect 73130 42160 73140 42220
rect 73200 42160 73210 42220
rect 72820 42152 73020 42158
rect 72710 42120 72790 42140
rect 72710 42060 72720 42120
rect 72780 42108 72790 42120
rect 72820 42118 72832 42152
rect 73008 42150 73020 42152
rect 73130 42150 73210 42160
rect 73680 42290 73690 42530
rect 73730 42290 73750 42530
rect 73680 42210 73750 42290
rect 73318 42152 73518 42158
rect 73318 42150 73330 42152
rect 73008 42120 73330 42150
rect 73008 42118 73020 42120
rect 72820 42112 73020 42118
rect 73318 42118 73330 42120
rect 73506 42118 73518 42152
rect 73318 42112 73518 42118
rect 73550 42120 73630 42140
rect 72782 42074 72790 42108
rect 72780 42060 72790 42074
rect 72710 42040 72790 42060
rect 72820 42064 73020 42070
rect 72820 42030 72832 42064
rect 73008 42060 73020 42064
rect 73318 42064 73518 42070
rect 73318 42060 73330 42064
rect 73008 42050 73330 42060
rect 73008 42030 73140 42050
rect 72820 42024 73020 42030
rect 73130 41990 73140 42030
rect 73200 42030 73330 42050
rect 73506 42030 73518 42064
rect 73550 42060 73560 42120
rect 73620 42060 73630 42120
rect 73550 42040 73630 42060
rect 73200 41990 73210 42030
rect 73318 42024 73518 42030
rect 73130 41980 73210 41990
rect 72600 40820 72670 41970
rect 72600 40560 72620 40820
rect 72660 40560 72670 40820
rect 73680 41970 73690 42210
rect 73730 41970 73750 42210
rect 73680 40820 73750 41970
rect 73130 40790 73210 40800
rect 72820 40752 73020 40758
rect 72710 40720 72790 40740
rect 72710 40660 72720 40720
rect 72780 40708 72790 40720
rect 72820 40718 72832 40752
rect 73008 40750 73020 40752
rect 73130 40750 73140 40790
rect 73008 40730 73140 40750
rect 73200 40750 73210 40790
rect 73318 40752 73518 40758
rect 73318 40750 73330 40752
rect 73200 40730 73330 40750
rect 73008 40720 73330 40730
rect 73008 40718 73020 40720
rect 72820 40712 73020 40718
rect 73318 40718 73330 40720
rect 73506 40718 73518 40752
rect 73318 40712 73518 40718
rect 73550 40720 73630 40740
rect 72782 40674 72790 40708
rect 72780 40660 72790 40674
rect 72710 40640 72790 40660
rect 72820 40664 73020 40670
rect 72820 40630 72832 40664
rect 73008 40660 73020 40664
rect 73318 40664 73518 40670
rect 73318 40660 73330 40664
rect 73008 40630 73330 40660
rect 73506 40630 73518 40664
rect 73550 40660 73560 40720
rect 73620 40660 73630 40720
rect 73550 40640 73630 40660
rect 72820 40624 73020 40630
rect 72600 40500 72670 40560
rect 72600 40260 72620 40500
rect 72660 40260 72670 40500
rect 73130 40620 73210 40630
rect 73318 40624 73518 40630
rect 73130 40560 73140 40620
rect 73200 40560 73210 40620
rect 73130 40510 73210 40560
rect 73130 40450 73140 40510
rect 73200 40450 73210 40510
rect 72820 40442 73020 40448
rect 72710 40410 72790 40430
rect 72710 40350 72720 40410
rect 72780 40398 72790 40410
rect 72820 40408 72832 40442
rect 73008 40440 73020 40442
rect 73130 40440 73210 40450
rect 73680 40580 73690 40820
rect 73730 40580 73750 40820
rect 73680 40500 73750 40580
rect 73318 40442 73518 40448
rect 73318 40440 73330 40442
rect 73008 40410 73330 40440
rect 73008 40408 73020 40410
rect 72820 40402 73020 40408
rect 73318 40408 73330 40410
rect 73506 40408 73518 40442
rect 73318 40402 73518 40408
rect 73550 40410 73630 40430
rect 72782 40364 72790 40398
rect 72780 40350 72790 40364
rect 72710 40330 72790 40350
rect 72820 40354 73020 40360
rect 72820 40320 72832 40354
rect 73008 40350 73020 40354
rect 73318 40354 73518 40360
rect 73318 40350 73330 40354
rect 73008 40340 73330 40350
rect 73008 40320 73140 40340
rect 72820 40314 73020 40320
rect 73130 40280 73140 40320
rect 73200 40320 73330 40340
rect 73506 40320 73518 40354
rect 73550 40350 73560 40410
rect 73620 40350 73630 40410
rect 73550 40330 73630 40350
rect 73200 40280 73210 40320
rect 73318 40314 73518 40320
rect 73130 40270 73210 40280
rect 72600 39690 72670 40260
rect 73680 40260 73690 40500
rect 73730 40260 73750 40500
rect 73680 39690 73750 40260
rect 72600 39680 72680 39690
rect 72600 39620 72610 39680
rect 72670 39620 72680 39680
rect 73670 39680 73750 39690
rect 73670 39620 73680 39680
rect 73740 39620 73750 39680
rect 73670 39610 73750 39620
rect 73780 66480 73810 67050
rect 73780 66470 73840 66480
rect 73780 66400 73840 66410
rect 73780 64770 73810 66400
rect 73870 65950 73900 67050
rect 73840 65940 73900 65950
rect 73840 65870 73900 65880
rect 73780 64760 73840 64770
rect 73780 64690 73840 64700
rect 73780 63060 73810 64690
rect 73870 64240 73900 65870
rect 73840 64230 73900 64240
rect 73840 64160 73900 64170
rect 73780 63050 73840 63060
rect 73780 62980 73840 62990
rect 73780 61350 73810 62980
rect 73870 62530 73900 64160
rect 73840 62520 73900 62530
rect 73840 62450 73900 62460
rect 73780 61340 73840 61350
rect 73780 61270 73840 61280
rect 73780 59640 73810 61270
rect 73870 60820 73900 62450
rect 73840 60810 73900 60820
rect 73840 60740 73900 60750
rect 73780 59630 73840 59640
rect 73780 59560 73840 59570
rect 73780 57930 73810 59560
rect 73870 59110 73900 60740
rect 73840 59100 73900 59110
rect 73840 59030 73900 59040
rect 73780 57920 73840 57930
rect 73780 57850 73840 57860
rect 73780 56220 73810 57850
rect 73870 57400 73900 59030
rect 73840 57390 73900 57400
rect 73840 57320 73900 57330
rect 73780 56210 73840 56220
rect 73780 56140 73840 56150
rect 73780 54510 73810 56140
rect 73870 55690 73900 57320
rect 73840 55680 73900 55690
rect 73840 55610 73900 55620
rect 73780 54500 73840 54510
rect 73780 54430 73840 54440
rect 73780 52800 73810 54430
rect 73870 53980 73900 55610
rect 73840 53970 73900 53980
rect 73840 53900 73900 53910
rect 73780 52790 73840 52800
rect 73780 52720 73840 52730
rect 73780 51090 73810 52720
rect 73870 52270 73900 53900
rect 73840 52260 73900 52270
rect 73840 52190 73900 52200
rect 73780 51080 73840 51090
rect 73780 51010 73840 51020
rect 73780 49380 73810 51010
rect 73870 50560 73900 52190
rect 73840 50550 73900 50560
rect 73840 50480 73900 50490
rect 73780 49370 73840 49380
rect 73780 49300 73840 49310
rect 73780 47670 73810 49300
rect 73870 48850 73900 50480
rect 73840 48840 73900 48850
rect 73840 48770 73900 48780
rect 73780 47660 73840 47670
rect 73780 47590 73840 47600
rect 73780 45960 73810 47590
rect 73870 47140 73900 48770
rect 73840 47130 73900 47140
rect 73840 47060 73900 47070
rect 73780 45950 73840 45960
rect 73780 45880 73840 45890
rect 73780 44250 73810 45880
rect 73870 45430 73900 47060
rect 73840 45420 73900 45430
rect 73840 45350 73900 45360
rect 73780 44240 73840 44250
rect 73780 44170 73840 44180
rect 73780 42540 73810 44170
rect 73870 43720 73900 45350
rect 73840 43710 73900 43720
rect 73840 43640 73900 43650
rect 73780 42530 73840 42540
rect 73780 42460 73840 42470
rect 73780 40830 73810 42460
rect 73870 42010 73900 43640
rect 73840 42000 73900 42010
rect 73840 41930 73900 41940
rect 73780 40820 73840 40830
rect 73780 40750 73840 40760
rect 69320 39220 69380 39230
rect 72310 39230 72570 39240
rect 69140 39160 69200 39170
rect 72370 39210 72570 39230
rect 72310 39160 72370 39170
rect 73780 38840 73810 40750
rect 73870 40300 73900 41930
rect 73840 40290 73900 40300
rect 73840 40220 73900 40230
rect 73870 39690 73900 40220
rect 73840 39680 73900 39690
rect 73840 39610 73900 39620
rect 73930 66390 73960 67050
rect 73930 66380 73990 66390
rect 73930 66310 73990 66320
rect 73930 64680 73960 66310
rect 73930 64670 73990 64680
rect 73930 64600 73990 64610
rect 73930 62970 73960 64600
rect 73930 62960 73990 62970
rect 73930 62890 73990 62900
rect 73930 61260 73960 62890
rect 73930 61250 73990 61260
rect 73930 61180 73990 61190
rect 73930 59550 73960 61180
rect 73930 59540 73990 59550
rect 73930 59470 73990 59480
rect 73930 57840 73960 59470
rect 73930 57830 73990 57840
rect 73930 57760 73990 57770
rect 73930 56130 73960 57760
rect 73930 56120 73990 56130
rect 73930 56050 73990 56060
rect 73930 54420 73960 56050
rect 73930 54410 73990 54420
rect 73930 54340 73990 54350
rect 73930 52710 73960 54340
rect 73930 52700 73990 52710
rect 73930 52630 73990 52640
rect 73930 51000 73960 52630
rect 73930 50990 73990 51000
rect 73930 50920 73990 50930
rect 73930 49290 73960 50920
rect 73930 49280 73990 49290
rect 73930 49210 73990 49220
rect 73930 47580 73960 49210
rect 73930 47570 73990 47580
rect 73930 47500 73990 47510
rect 73930 45870 73960 47500
rect 73930 45860 73990 45870
rect 73930 45790 73990 45800
rect 73930 44160 73960 45790
rect 73930 44150 73990 44160
rect 73930 44080 73990 44090
rect 73930 42450 73960 44080
rect 73930 42440 73990 42450
rect 73930 42370 73990 42380
rect 73930 40740 73960 42370
rect 73930 40730 73990 40740
rect 73930 40660 73990 40670
rect 73930 39240 73960 40660
rect 74050 39690 74080 67050
rect 74170 39690 74200 67050
rect 74290 39690 74320 67050
rect 74410 39690 74440 67050
rect 74530 39690 74560 67050
rect 74650 39690 74680 67050
rect 76810 39690 76840 67050
rect 76930 39690 76960 67050
rect 77050 39690 77080 67050
rect 77170 39690 77200 67050
rect 77290 39690 77320 67050
rect 77410 39690 77440 67050
rect 77530 66390 77560 67050
rect 77500 66380 77560 66390
rect 77500 66310 77560 66320
rect 77530 64680 77560 66310
rect 77500 64670 77560 64680
rect 77500 64600 77560 64610
rect 77530 62970 77560 64600
rect 77500 62960 77560 62970
rect 77500 62890 77560 62900
rect 77530 61260 77560 62890
rect 77500 61250 77560 61260
rect 77500 61180 77560 61190
rect 77530 59550 77560 61180
rect 77500 59540 77560 59550
rect 77500 59470 77560 59480
rect 77530 57840 77560 59470
rect 77500 57830 77560 57840
rect 77500 57760 77560 57770
rect 77530 56130 77560 57760
rect 77500 56120 77560 56130
rect 77500 56050 77560 56060
rect 77530 54420 77560 56050
rect 77500 54410 77560 54420
rect 77500 54340 77560 54350
rect 77530 52710 77560 54340
rect 77500 52700 77560 52710
rect 77500 52630 77560 52640
rect 77530 51000 77560 52630
rect 77500 50990 77560 51000
rect 77500 50920 77560 50930
rect 77530 49290 77560 50920
rect 77500 49280 77560 49290
rect 77500 49210 77560 49220
rect 77530 47580 77560 49210
rect 77500 47570 77560 47580
rect 77500 47500 77560 47510
rect 77530 45870 77560 47500
rect 77500 45860 77560 45870
rect 77500 45790 77560 45800
rect 77530 44160 77560 45790
rect 77500 44150 77560 44160
rect 77500 44080 77560 44090
rect 77530 42450 77560 44080
rect 77500 42440 77560 42450
rect 77500 42370 77560 42380
rect 77530 40740 77560 42370
rect 77500 40730 77560 40740
rect 77500 40660 77560 40670
rect 77530 39240 77560 40660
rect 77590 66470 77660 67050
rect 77590 66210 77610 66470
rect 77650 66210 77660 66470
rect 78670 66470 78740 67050
rect 78120 66440 78200 66450
rect 77810 66402 78010 66408
rect 77700 66370 77780 66390
rect 77700 66310 77710 66370
rect 77770 66358 77780 66370
rect 77810 66368 77822 66402
rect 77998 66400 78010 66402
rect 78120 66400 78130 66440
rect 77998 66380 78130 66400
rect 78190 66400 78200 66440
rect 78308 66402 78508 66408
rect 78308 66400 78320 66402
rect 78190 66380 78320 66400
rect 77998 66370 78320 66380
rect 77998 66368 78010 66370
rect 77810 66362 78010 66368
rect 78308 66368 78320 66370
rect 78496 66368 78508 66402
rect 78308 66362 78508 66368
rect 78540 66370 78620 66390
rect 77772 66324 77780 66358
rect 77770 66310 77780 66324
rect 77700 66290 77780 66310
rect 77810 66314 78010 66320
rect 77810 66280 77822 66314
rect 77998 66310 78010 66314
rect 78308 66314 78508 66320
rect 78308 66310 78320 66314
rect 77998 66280 78320 66310
rect 78496 66280 78508 66314
rect 78540 66310 78550 66370
rect 78610 66310 78620 66370
rect 78540 66290 78620 66310
rect 77810 66274 78010 66280
rect 77590 66150 77660 66210
rect 77590 65910 77610 66150
rect 77650 65910 77660 66150
rect 78120 66270 78200 66280
rect 78308 66274 78508 66280
rect 78120 66210 78130 66270
rect 78190 66210 78200 66270
rect 78120 66160 78200 66210
rect 78120 66100 78130 66160
rect 78190 66100 78200 66160
rect 77810 66092 78010 66098
rect 77700 66060 77780 66080
rect 77700 66000 77710 66060
rect 77770 66048 77780 66060
rect 77810 66058 77822 66092
rect 77998 66090 78010 66092
rect 78120 66090 78200 66100
rect 78670 66230 78680 66470
rect 78720 66230 78740 66470
rect 78670 66150 78740 66230
rect 78308 66092 78508 66098
rect 78308 66090 78320 66092
rect 77998 66060 78320 66090
rect 77998 66058 78010 66060
rect 77810 66052 78010 66058
rect 78308 66058 78320 66060
rect 78496 66058 78508 66092
rect 78308 66052 78508 66058
rect 78540 66060 78620 66080
rect 77772 66014 77780 66048
rect 77770 66000 77780 66014
rect 77700 65980 77780 66000
rect 77810 66004 78010 66010
rect 77810 65970 77822 66004
rect 77998 66000 78010 66004
rect 78308 66004 78508 66010
rect 78308 66000 78320 66004
rect 77998 65990 78320 66000
rect 77998 65970 78130 65990
rect 77810 65964 78010 65970
rect 78120 65930 78130 65970
rect 78190 65970 78320 65990
rect 78496 65970 78508 66004
rect 78540 66000 78550 66060
rect 78610 66000 78620 66060
rect 78540 65980 78620 66000
rect 78190 65930 78200 65970
rect 78308 65964 78508 65970
rect 78120 65920 78200 65930
rect 77590 64760 77660 65910
rect 77590 64500 77610 64760
rect 77650 64500 77660 64760
rect 78670 65910 78680 66150
rect 78720 65910 78740 66150
rect 78670 64760 78740 65910
rect 78120 64730 78200 64740
rect 77810 64692 78010 64698
rect 77700 64660 77780 64680
rect 77700 64600 77710 64660
rect 77770 64648 77780 64660
rect 77810 64658 77822 64692
rect 77998 64690 78010 64692
rect 78120 64690 78130 64730
rect 77998 64670 78130 64690
rect 78190 64690 78200 64730
rect 78308 64692 78508 64698
rect 78308 64690 78320 64692
rect 78190 64670 78320 64690
rect 77998 64660 78320 64670
rect 77998 64658 78010 64660
rect 77810 64652 78010 64658
rect 78308 64658 78320 64660
rect 78496 64658 78508 64692
rect 78308 64652 78508 64658
rect 78540 64660 78620 64680
rect 77772 64614 77780 64648
rect 77770 64600 77780 64614
rect 77700 64580 77780 64600
rect 77810 64604 78010 64610
rect 77810 64570 77822 64604
rect 77998 64600 78010 64604
rect 78308 64604 78508 64610
rect 78308 64600 78320 64604
rect 77998 64570 78320 64600
rect 78496 64570 78508 64604
rect 78540 64600 78550 64660
rect 78610 64600 78620 64660
rect 78540 64580 78620 64600
rect 77810 64564 78010 64570
rect 77590 64440 77660 64500
rect 77590 64200 77610 64440
rect 77650 64200 77660 64440
rect 78120 64560 78200 64570
rect 78308 64564 78508 64570
rect 78120 64500 78130 64560
rect 78190 64500 78200 64560
rect 78120 64450 78200 64500
rect 78120 64390 78130 64450
rect 78190 64390 78200 64450
rect 77810 64382 78010 64388
rect 77700 64350 77780 64370
rect 77700 64290 77710 64350
rect 77770 64338 77780 64350
rect 77810 64348 77822 64382
rect 77998 64380 78010 64382
rect 78120 64380 78200 64390
rect 78670 64520 78680 64760
rect 78720 64520 78740 64760
rect 78670 64440 78740 64520
rect 78308 64382 78508 64388
rect 78308 64380 78320 64382
rect 77998 64350 78320 64380
rect 77998 64348 78010 64350
rect 77810 64342 78010 64348
rect 78308 64348 78320 64350
rect 78496 64348 78508 64382
rect 78308 64342 78508 64348
rect 78540 64350 78620 64370
rect 77772 64304 77780 64338
rect 77770 64290 77780 64304
rect 77700 64270 77780 64290
rect 77810 64294 78010 64300
rect 77810 64260 77822 64294
rect 77998 64290 78010 64294
rect 78308 64294 78508 64300
rect 78308 64290 78320 64294
rect 77998 64280 78320 64290
rect 77998 64260 78130 64280
rect 77810 64254 78010 64260
rect 78120 64220 78130 64260
rect 78190 64260 78320 64280
rect 78496 64260 78508 64294
rect 78540 64290 78550 64350
rect 78610 64290 78620 64350
rect 78540 64270 78620 64290
rect 78190 64220 78200 64260
rect 78308 64254 78508 64260
rect 78120 64210 78200 64220
rect 77590 63050 77660 64200
rect 77590 62790 77610 63050
rect 77650 62790 77660 63050
rect 78670 64200 78680 64440
rect 78720 64200 78740 64440
rect 78670 63050 78740 64200
rect 78120 63020 78200 63030
rect 77810 62982 78010 62988
rect 77700 62950 77780 62970
rect 77700 62890 77710 62950
rect 77770 62938 77780 62950
rect 77810 62948 77822 62982
rect 77998 62980 78010 62982
rect 78120 62980 78130 63020
rect 77998 62960 78130 62980
rect 78190 62980 78200 63020
rect 78308 62982 78508 62988
rect 78308 62980 78320 62982
rect 78190 62960 78320 62980
rect 77998 62950 78320 62960
rect 77998 62948 78010 62950
rect 77810 62942 78010 62948
rect 78308 62948 78320 62950
rect 78496 62948 78508 62982
rect 78308 62942 78508 62948
rect 78540 62950 78620 62970
rect 77772 62904 77780 62938
rect 77770 62890 77780 62904
rect 77700 62870 77780 62890
rect 77810 62894 78010 62900
rect 77810 62860 77822 62894
rect 77998 62890 78010 62894
rect 78308 62894 78508 62900
rect 78308 62890 78320 62894
rect 77998 62860 78320 62890
rect 78496 62860 78508 62894
rect 78540 62890 78550 62950
rect 78610 62890 78620 62950
rect 78540 62870 78620 62890
rect 77810 62854 78010 62860
rect 77590 62730 77660 62790
rect 77590 62490 77610 62730
rect 77650 62490 77660 62730
rect 78120 62850 78200 62860
rect 78308 62854 78508 62860
rect 78120 62790 78130 62850
rect 78190 62790 78200 62850
rect 78120 62740 78200 62790
rect 78120 62680 78130 62740
rect 78190 62680 78200 62740
rect 77810 62672 78010 62678
rect 77700 62640 77780 62660
rect 77700 62580 77710 62640
rect 77770 62628 77780 62640
rect 77810 62638 77822 62672
rect 77998 62670 78010 62672
rect 78120 62670 78200 62680
rect 78670 62810 78680 63050
rect 78720 62810 78740 63050
rect 78670 62730 78740 62810
rect 78308 62672 78508 62678
rect 78308 62670 78320 62672
rect 77998 62640 78320 62670
rect 77998 62638 78010 62640
rect 77810 62632 78010 62638
rect 78308 62638 78320 62640
rect 78496 62638 78508 62672
rect 78308 62632 78508 62638
rect 78540 62640 78620 62660
rect 77772 62594 77780 62628
rect 77770 62580 77780 62594
rect 77700 62560 77780 62580
rect 77810 62584 78010 62590
rect 77810 62550 77822 62584
rect 77998 62580 78010 62584
rect 78308 62584 78508 62590
rect 78308 62580 78320 62584
rect 77998 62570 78320 62580
rect 77998 62550 78130 62570
rect 77810 62544 78010 62550
rect 78120 62510 78130 62550
rect 78190 62550 78320 62570
rect 78496 62550 78508 62584
rect 78540 62580 78550 62640
rect 78610 62580 78620 62640
rect 78540 62560 78620 62580
rect 78190 62510 78200 62550
rect 78308 62544 78508 62550
rect 78120 62500 78200 62510
rect 77590 61340 77660 62490
rect 77590 61080 77610 61340
rect 77650 61080 77660 61340
rect 78670 62490 78680 62730
rect 78720 62490 78740 62730
rect 78670 61340 78740 62490
rect 78120 61310 78200 61320
rect 77810 61272 78010 61278
rect 77700 61240 77780 61260
rect 77700 61180 77710 61240
rect 77770 61228 77780 61240
rect 77810 61238 77822 61272
rect 77998 61270 78010 61272
rect 78120 61270 78130 61310
rect 77998 61250 78130 61270
rect 78190 61270 78200 61310
rect 78308 61272 78508 61278
rect 78308 61270 78320 61272
rect 78190 61250 78320 61270
rect 77998 61240 78320 61250
rect 77998 61238 78010 61240
rect 77810 61232 78010 61238
rect 78308 61238 78320 61240
rect 78496 61238 78508 61272
rect 78308 61232 78508 61238
rect 78540 61240 78620 61260
rect 77772 61194 77780 61228
rect 77770 61180 77780 61194
rect 77700 61160 77780 61180
rect 77810 61184 78010 61190
rect 77810 61150 77822 61184
rect 77998 61180 78010 61184
rect 78308 61184 78508 61190
rect 78308 61180 78320 61184
rect 77998 61150 78320 61180
rect 78496 61150 78508 61184
rect 78540 61180 78550 61240
rect 78610 61180 78620 61240
rect 78540 61160 78620 61180
rect 77810 61144 78010 61150
rect 77590 61020 77660 61080
rect 77590 60780 77610 61020
rect 77650 60780 77660 61020
rect 78120 61140 78200 61150
rect 78308 61144 78508 61150
rect 78120 61080 78130 61140
rect 78190 61080 78200 61140
rect 78120 61030 78200 61080
rect 78120 60970 78130 61030
rect 78190 60970 78200 61030
rect 77810 60962 78010 60968
rect 77700 60930 77780 60950
rect 77700 60870 77710 60930
rect 77770 60918 77780 60930
rect 77810 60928 77822 60962
rect 77998 60960 78010 60962
rect 78120 60960 78200 60970
rect 78670 61100 78680 61340
rect 78720 61100 78740 61340
rect 78670 61020 78740 61100
rect 78308 60962 78508 60968
rect 78308 60960 78320 60962
rect 77998 60930 78320 60960
rect 77998 60928 78010 60930
rect 77810 60922 78010 60928
rect 78308 60928 78320 60930
rect 78496 60928 78508 60962
rect 78308 60922 78508 60928
rect 78540 60930 78620 60950
rect 77772 60884 77780 60918
rect 77770 60870 77780 60884
rect 77700 60850 77780 60870
rect 77810 60874 78010 60880
rect 77810 60840 77822 60874
rect 77998 60870 78010 60874
rect 78308 60874 78508 60880
rect 78308 60870 78320 60874
rect 77998 60860 78320 60870
rect 77998 60840 78130 60860
rect 77810 60834 78010 60840
rect 78120 60800 78130 60840
rect 78190 60840 78320 60860
rect 78496 60840 78508 60874
rect 78540 60870 78550 60930
rect 78610 60870 78620 60930
rect 78540 60850 78620 60870
rect 78190 60800 78200 60840
rect 78308 60834 78508 60840
rect 78120 60790 78200 60800
rect 77590 59630 77660 60780
rect 77590 59370 77610 59630
rect 77650 59370 77660 59630
rect 78670 60780 78680 61020
rect 78720 60780 78740 61020
rect 78670 59630 78740 60780
rect 78120 59600 78200 59610
rect 77810 59562 78010 59568
rect 77700 59530 77780 59550
rect 77700 59470 77710 59530
rect 77770 59518 77780 59530
rect 77810 59528 77822 59562
rect 77998 59560 78010 59562
rect 78120 59560 78130 59600
rect 77998 59540 78130 59560
rect 78190 59560 78200 59600
rect 78308 59562 78508 59568
rect 78308 59560 78320 59562
rect 78190 59540 78320 59560
rect 77998 59530 78320 59540
rect 77998 59528 78010 59530
rect 77810 59522 78010 59528
rect 78308 59528 78320 59530
rect 78496 59528 78508 59562
rect 78308 59522 78508 59528
rect 78540 59530 78620 59550
rect 77772 59484 77780 59518
rect 77770 59470 77780 59484
rect 77700 59450 77780 59470
rect 77810 59474 78010 59480
rect 77810 59440 77822 59474
rect 77998 59470 78010 59474
rect 78308 59474 78508 59480
rect 78308 59470 78320 59474
rect 77998 59440 78320 59470
rect 78496 59440 78508 59474
rect 78540 59470 78550 59530
rect 78610 59470 78620 59530
rect 78540 59450 78620 59470
rect 77810 59434 78010 59440
rect 77590 59310 77660 59370
rect 77590 59070 77610 59310
rect 77650 59070 77660 59310
rect 78120 59430 78200 59440
rect 78308 59434 78508 59440
rect 78120 59370 78130 59430
rect 78190 59370 78200 59430
rect 78120 59320 78200 59370
rect 78120 59260 78130 59320
rect 78190 59260 78200 59320
rect 77810 59252 78010 59258
rect 77700 59220 77780 59240
rect 77700 59160 77710 59220
rect 77770 59208 77780 59220
rect 77810 59218 77822 59252
rect 77998 59250 78010 59252
rect 78120 59250 78200 59260
rect 78670 59390 78680 59630
rect 78720 59390 78740 59630
rect 78670 59310 78740 59390
rect 78308 59252 78508 59258
rect 78308 59250 78320 59252
rect 77998 59220 78320 59250
rect 77998 59218 78010 59220
rect 77810 59212 78010 59218
rect 78308 59218 78320 59220
rect 78496 59218 78508 59252
rect 78308 59212 78508 59218
rect 78540 59220 78620 59240
rect 77772 59174 77780 59208
rect 77770 59160 77780 59174
rect 77700 59140 77780 59160
rect 77810 59164 78010 59170
rect 77810 59130 77822 59164
rect 77998 59160 78010 59164
rect 78308 59164 78508 59170
rect 78308 59160 78320 59164
rect 77998 59150 78320 59160
rect 77998 59130 78130 59150
rect 77810 59124 78010 59130
rect 78120 59090 78130 59130
rect 78190 59130 78320 59150
rect 78496 59130 78508 59164
rect 78540 59160 78550 59220
rect 78610 59160 78620 59220
rect 78540 59140 78620 59160
rect 78190 59090 78200 59130
rect 78308 59124 78508 59130
rect 78120 59080 78200 59090
rect 77590 57920 77660 59070
rect 77590 57660 77610 57920
rect 77650 57660 77660 57920
rect 78670 59070 78680 59310
rect 78720 59070 78740 59310
rect 78670 57920 78740 59070
rect 78120 57890 78200 57900
rect 77810 57852 78010 57858
rect 77700 57820 77780 57840
rect 77700 57760 77710 57820
rect 77770 57808 77780 57820
rect 77810 57818 77822 57852
rect 77998 57850 78010 57852
rect 78120 57850 78130 57890
rect 77998 57830 78130 57850
rect 78190 57850 78200 57890
rect 78308 57852 78508 57858
rect 78308 57850 78320 57852
rect 78190 57830 78320 57850
rect 77998 57820 78320 57830
rect 77998 57818 78010 57820
rect 77810 57812 78010 57818
rect 78308 57818 78320 57820
rect 78496 57818 78508 57852
rect 78308 57812 78508 57818
rect 78540 57820 78620 57840
rect 77772 57774 77780 57808
rect 77770 57760 77780 57774
rect 77700 57740 77780 57760
rect 77810 57764 78010 57770
rect 77810 57730 77822 57764
rect 77998 57760 78010 57764
rect 78308 57764 78508 57770
rect 78308 57760 78320 57764
rect 77998 57730 78320 57760
rect 78496 57730 78508 57764
rect 78540 57760 78550 57820
rect 78610 57760 78620 57820
rect 78540 57740 78620 57760
rect 77810 57724 78010 57730
rect 77590 57600 77660 57660
rect 77590 57360 77610 57600
rect 77650 57360 77660 57600
rect 78120 57720 78200 57730
rect 78308 57724 78508 57730
rect 78120 57660 78130 57720
rect 78190 57660 78200 57720
rect 78120 57610 78200 57660
rect 78120 57550 78130 57610
rect 78190 57550 78200 57610
rect 77810 57542 78010 57548
rect 77700 57510 77780 57530
rect 77700 57450 77710 57510
rect 77770 57498 77780 57510
rect 77810 57508 77822 57542
rect 77998 57540 78010 57542
rect 78120 57540 78200 57550
rect 78670 57680 78680 57920
rect 78720 57680 78740 57920
rect 78670 57600 78740 57680
rect 78308 57542 78508 57548
rect 78308 57540 78320 57542
rect 77998 57510 78320 57540
rect 77998 57508 78010 57510
rect 77810 57502 78010 57508
rect 78308 57508 78320 57510
rect 78496 57508 78508 57542
rect 78308 57502 78508 57508
rect 78540 57510 78620 57530
rect 77772 57464 77780 57498
rect 77770 57450 77780 57464
rect 77700 57430 77780 57450
rect 77810 57454 78010 57460
rect 77810 57420 77822 57454
rect 77998 57450 78010 57454
rect 78308 57454 78508 57460
rect 78308 57450 78320 57454
rect 77998 57440 78320 57450
rect 77998 57420 78130 57440
rect 77810 57414 78010 57420
rect 78120 57380 78130 57420
rect 78190 57420 78320 57440
rect 78496 57420 78508 57454
rect 78540 57450 78550 57510
rect 78610 57450 78620 57510
rect 78540 57430 78620 57450
rect 78190 57380 78200 57420
rect 78308 57414 78508 57420
rect 78120 57370 78200 57380
rect 77590 56210 77660 57360
rect 77590 55950 77610 56210
rect 77650 55950 77660 56210
rect 78670 57360 78680 57600
rect 78720 57360 78740 57600
rect 78670 56210 78740 57360
rect 78120 56180 78200 56190
rect 77810 56142 78010 56148
rect 77700 56110 77780 56130
rect 77700 56050 77710 56110
rect 77770 56098 77780 56110
rect 77810 56108 77822 56142
rect 77998 56140 78010 56142
rect 78120 56140 78130 56180
rect 77998 56120 78130 56140
rect 78190 56140 78200 56180
rect 78308 56142 78508 56148
rect 78308 56140 78320 56142
rect 78190 56120 78320 56140
rect 77998 56110 78320 56120
rect 77998 56108 78010 56110
rect 77810 56102 78010 56108
rect 78308 56108 78320 56110
rect 78496 56108 78508 56142
rect 78308 56102 78508 56108
rect 78540 56110 78620 56130
rect 77772 56064 77780 56098
rect 77770 56050 77780 56064
rect 77700 56030 77780 56050
rect 77810 56054 78010 56060
rect 77810 56020 77822 56054
rect 77998 56050 78010 56054
rect 78308 56054 78508 56060
rect 78308 56050 78320 56054
rect 77998 56020 78320 56050
rect 78496 56020 78508 56054
rect 78540 56050 78550 56110
rect 78610 56050 78620 56110
rect 78540 56030 78620 56050
rect 77810 56014 78010 56020
rect 77590 55890 77660 55950
rect 77590 55650 77610 55890
rect 77650 55650 77660 55890
rect 78120 56010 78200 56020
rect 78308 56014 78508 56020
rect 78120 55950 78130 56010
rect 78190 55950 78200 56010
rect 78120 55900 78200 55950
rect 78120 55840 78130 55900
rect 78190 55840 78200 55900
rect 77810 55832 78010 55838
rect 77700 55800 77780 55820
rect 77700 55740 77710 55800
rect 77770 55788 77780 55800
rect 77810 55798 77822 55832
rect 77998 55830 78010 55832
rect 78120 55830 78200 55840
rect 78670 55970 78680 56210
rect 78720 55970 78740 56210
rect 78670 55890 78740 55970
rect 78308 55832 78508 55838
rect 78308 55830 78320 55832
rect 77998 55800 78320 55830
rect 77998 55798 78010 55800
rect 77810 55792 78010 55798
rect 78308 55798 78320 55800
rect 78496 55798 78508 55832
rect 78308 55792 78508 55798
rect 78540 55800 78620 55820
rect 77772 55754 77780 55788
rect 77770 55740 77780 55754
rect 77700 55720 77780 55740
rect 77810 55744 78010 55750
rect 77810 55710 77822 55744
rect 77998 55740 78010 55744
rect 78308 55744 78508 55750
rect 78308 55740 78320 55744
rect 77998 55730 78320 55740
rect 77998 55710 78130 55730
rect 77810 55704 78010 55710
rect 78120 55670 78130 55710
rect 78190 55710 78320 55730
rect 78496 55710 78508 55744
rect 78540 55740 78550 55800
rect 78610 55740 78620 55800
rect 78540 55720 78620 55740
rect 78190 55670 78200 55710
rect 78308 55704 78508 55710
rect 78120 55660 78200 55670
rect 77590 54500 77660 55650
rect 77590 54240 77610 54500
rect 77650 54240 77660 54500
rect 78670 55650 78680 55890
rect 78720 55650 78740 55890
rect 78670 54500 78740 55650
rect 78120 54470 78200 54480
rect 77810 54432 78010 54438
rect 77700 54400 77780 54420
rect 77700 54340 77710 54400
rect 77770 54388 77780 54400
rect 77810 54398 77822 54432
rect 77998 54430 78010 54432
rect 78120 54430 78130 54470
rect 77998 54410 78130 54430
rect 78190 54430 78200 54470
rect 78308 54432 78508 54438
rect 78308 54430 78320 54432
rect 78190 54410 78320 54430
rect 77998 54400 78320 54410
rect 77998 54398 78010 54400
rect 77810 54392 78010 54398
rect 78308 54398 78320 54400
rect 78496 54398 78508 54432
rect 78308 54392 78508 54398
rect 78540 54400 78620 54420
rect 77772 54354 77780 54388
rect 77770 54340 77780 54354
rect 77700 54320 77780 54340
rect 77810 54344 78010 54350
rect 77810 54310 77822 54344
rect 77998 54340 78010 54344
rect 78308 54344 78508 54350
rect 78308 54340 78320 54344
rect 77998 54310 78320 54340
rect 78496 54310 78508 54344
rect 78540 54340 78550 54400
rect 78610 54340 78620 54400
rect 78540 54320 78620 54340
rect 77810 54304 78010 54310
rect 77590 54180 77660 54240
rect 77590 53940 77610 54180
rect 77650 53940 77660 54180
rect 78120 54300 78200 54310
rect 78308 54304 78508 54310
rect 78120 54240 78130 54300
rect 78190 54240 78200 54300
rect 78120 54190 78200 54240
rect 78120 54130 78130 54190
rect 78190 54130 78200 54190
rect 77810 54122 78010 54128
rect 77700 54090 77780 54110
rect 77700 54030 77710 54090
rect 77770 54078 77780 54090
rect 77810 54088 77822 54122
rect 77998 54120 78010 54122
rect 78120 54120 78200 54130
rect 78670 54260 78680 54500
rect 78720 54260 78740 54500
rect 78670 54180 78740 54260
rect 78308 54122 78508 54128
rect 78308 54120 78320 54122
rect 77998 54090 78320 54120
rect 77998 54088 78010 54090
rect 77810 54082 78010 54088
rect 78308 54088 78320 54090
rect 78496 54088 78508 54122
rect 78308 54082 78508 54088
rect 78540 54090 78620 54110
rect 77772 54044 77780 54078
rect 77770 54030 77780 54044
rect 77700 54010 77780 54030
rect 77810 54034 78010 54040
rect 77810 54000 77822 54034
rect 77998 54030 78010 54034
rect 78308 54034 78508 54040
rect 78308 54030 78320 54034
rect 77998 54020 78320 54030
rect 77998 54000 78130 54020
rect 77810 53994 78010 54000
rect 78120 53960 78130 54000
rect 78190 54000 78320 54020
rect 78496 54000 78508 54034
rect 78540 54030 78550 54090
rect 78610 54030 78620 54090
rect 78540 54010 78620 54030
rect 78190 53960 78200 54000
rect 78308 53994 78508 54000
rect 78120 53950 78200 53960
rect 77590 52790 77660 53940
rect 77590 52530 77610 52790
rect 77650 52530 77660 52790
rect 78670 53940 78680 54180
rect 78720 53940 78740 54180
rect 78670 52790 78740 53940
rect 78120 52760 78200 52770
rect 77810 52722 78010 52728
rect 77700 52690 77780 52710
rect 77700 52630 77710 52690
rect 77770 52678 77780 52690
rect 77810 52688 77822 52722
rect 77998 52720 78010 52722
rect 78120 52720 78130 52760
rect 77998 52700 78130 52720
rect 78190 52720 78200 52760
rect 78308 52722 78508 52728
rect 78308 52720 78320 52722
rect 78190 52700 78320 52720
rect 77998 52690 78320 52700
rect 77998 52688 78010 52690
rect 77810 52682 78010 52688
rect 78308 52688 78320 52690
rect 78496 52688 78508 52722
rect 78308 52682 78508 52688
rect 78540 52690 78620 52710
rect 77772 52644 77780 52678
rect 77770 52630 77780 52644
rect 77700 52610 77780 52630
rect 77810 52634 78010 52640
rect 77810 52600 77822 52634
rect 77998 52630 78010 52634
rect 78308 52634 78508 52640
rect 78308 52630 78320 52634
rect 77998 52600 78320 52630
rect 78496 52600 78508 52634
rect 78540 52630 78550 52690
rect 78610 52630 78620 52690
rect 78540 52610 78620 52630
rect 77810 52594 78010 52600
rect 77590 52470 77660 52530
rect 77590 52230 77610 52470
rect 77650 52230 77660 52470
rect 78120 52590 78200 52600
rect 78308 52594 78508 52600
rect 78120 52530 78130 52590
rect 78190 52530 78200 52590
rect 78120 52480 78200 52530
rect 78120 52420 78130 52480
rect 78190 52420 78200 52480
rect 77810 52412 78010 52418
rect 77700 52380 77780 52400
rect 77700 52320 77710 52380
rect 77770 52368 77780 52380
rect 77810 52378 77822 52412
rect 77998 52410 78010 52412
rect 78120 52410 78200 52420
rect 78670 52550 78680 52790
rect 78720 52550 78740 52790
rect 78670 52470 78740 52550
rect 78308 52412 78508 52418
rect 78308 52410 78320 52412
rect 77998 52380 78320 52410
rect 77998 52378 78010 52380
rect 77810 52372 78010 52378
rect 78308 52378 78320 52380
rect 78496 52378 78508 52412
rect 78308 52372 78508 52378
rect 78540 52380 78620 52400
rect 77772 52334 77780 52368
rect 77770 52320 77780 52334
rect 77700 52300 77780 52320
rect 77810 52324 78010 52330
rect 77810 52290 77822 52324
rect 77998 52320 78010 52324
rect 78308 52324 78508 52330
rect 78308 52320 78320 52324
rect 77998 52310 78320 52320
rect 77998 52290 78130 52310
rect 77810 52284 78010 52290
rect 78120 52250 78130 52290
rect 78190 52290 78320 52310
rect 78496 52290 78508 52324
rect 78540 52320 78550 52380
rect 78610 52320 78620 52380
rect 78540 52300 78620 52320
rect 78190 52250 78200 52290
rect 78308 52284 78508 52290
rect 78120 52240 78200 52250
rect 77590 51080 77660 52230
rect 77590 50820 77610 51080
rect 77650 50820 77660 51080
rect 78670 52230 78680 52470
rect 78720 52230 78740 52470
rect 78670 51080 78740 52230
rect 78120 51050 78200 51060
rect 77810 51012 78010 51018
rect 77700 50980 77780 51000
rect 77700 50920 77710 50980
rect 77770 50968 77780 50980
rect 77810 50978 77822 51012
rect 77998 51010 78010 51012
rect 78120 51010 78130 51050
rect 77998 50990 78130 51010
rect 78190 51010 78200 51050
rect 78308 51012 78508 51018
rect 78308 51010 78320 51012
rect 78190 50990 78320 51010
rect 77998 50980 78320 50990
rect 77998 50978 78010 50980
rect 77810 50972 78010 50978
rect 78308 50978 78320 50980
rect 78496 50978 78508 51012
rect 78308 50972 78508 50978
rect 78540 50980 78620 51000
rect 77772 50934 77780 50968
rect 77770 50920 77780 50934
rect 77700 50900 77780 50920
rect 77810 50924 78010 50930
rect 77810 50890 77822 50924
rect 77998 50920 78010 50924
rect 78308 50924 78508 50930
rect 78308 50920 78320 50924
rect 77998 50890 78320 50920
rect 78496 50890 78508 50924
rect 78540 50920 78550 50980
rect 78610 50920 78620 50980
rect 78540 50900 78620 50920
rect 77810 50884 78010 50890
rect 77590 50760 77660 50820
rect 77590 50520 77610 50760
rect 77650 50520 77660 50760
rect 78120 50880 78200 50890
rect 78308 50884 78508 50890
rect 78120 50820 78130 50880
rect 78190 50820 78200 50880
rect 78120 50770 78200 50820
rect 78120 50710 78130 50770
rect 78190 50710 78200 50770
rect 77810 50702 78010 50708
rect 77700 50670 77780 50690
rect 77700 50610 77710 50670
rect 77770 50658 77780 50670
rect 77810 50668 77822 50702
rect 77998 50700 78010 50702
rect 78120 50700 78200 50710
rect 78670 50840 78680 51080
rect 78720 50840 78740 51080
rect 78670 50760 78740 50840
rect 78308 50702 78508 50708
rect 78308 50700 78320 50702
rect 77998 50670 78320 50700
rect 77998 50668 78010 50670
rect 77810 50662 78010 50668
rect 78308 50668 78320 50670
rect 78496 50668 78508 50702
rect 78308 50662 78508 50668
rect 78540 50670 78620 50690
rect 77772 50624 77780 50658
rect 77770 50610 77780 50624
rect 77700 50590 77780 50610
rect 77810 50614 78010 50620
rect 77810 50580 77822 50614
rect 77998 50610 78010 50614
rect 78308 50614 78508 50620
rect 78308 50610 78320 50614
rect 77998 50600 78320 50610
rect 77998 50580 78130 50600
rect 77810 50574 78010 50580
rect 78120 50540 78130 50580
rect 78190 50580 78320 50600
rect 78496 50580 78508 50614
rect 78540 50610 78550 50670
rect 78610 50610 78620 50670
rect 78540 50590 78620 50610
rect 78190 50540 78200 50580
rect 78308 50574 78508 50580
rect 78120 50530 78200 50540
rect 77590 49370 77660 50520
rect 77590 49110 77610 49370
rect 77650 49110 77660 49370
rect 78670 50520 78680 50760
rect 78720 50520 78740 50760
rect 78670 49370 78740 50520
rect 78120 49340 78200 49350
rect 77810 49302 78010 49308
rect 77700 49270 77780 49290
rect 77700 49210 77710 49270
rect 77770 49258 77780 49270
rect 77810 49268 77822 49302
rect 77998 49300 78010 49302
rect 78120 49300 78130 49340
rect 77998 49280 78130 49300
rect 78190 49300 78200 49340
rect 78308 49302 78508 49308
rect 78308 49300 78320 49302
rect 78190 49280 78320 49300
rect 77998 49270 78320 49280
rect 77998 49268 78010 49270
rect 77810 49262 78010 49268
rect 78308 49268 78320 49270
rect 78496 49268 78508 49302
rect 78308 49262 78508 49268
rect 78540 49270 78620 49290
rect 77772 49224 77780 49258
rect 77770 49210 77780 49224
rect 77700 49190 77780 49210
rect 77810 49214 78010 49220
rect 77810 49180 77822 49214
rect 77998 49210 78010 49214
rect 78308 49214 78508 49220
rect 78308 49210 78320 49214
rect 77998 49180 78320 49210
rect 78496 49180 78508 49214
rect 78540 49210 78550 49270
rect 78610 49210 78620 49270
rect 78540 49190 78620 49210
rect 77810 49174 78010 49180
rect 77590 49050 77660 49110
rect 77590 48810 77610 49050
rect 77650 48810 77660 49050
rect 78120 49170 78200 49180
rect 78308 49174 78508 49180
rect 78120 49110 78130 49170
rect 78190 49110 78200 49170
rect 78120 49060 78200 49110
rect 78120 49000 78130 49060
rect 78190 49000 78200 49060
rect 77810 48992 78010 48998
rect 77700 48960 77780 48980
rect 77700 48900 77710 48960
rect 77770 48948 77780 48960
rect 77810 48958 77822 48992
rect 77998 48990 78010 48992
rect 78120 48990 78200 49000
rect 78670 49130 78680 49370
rect 78720 49130 78740 49370
rect 78670 49050 78740 49130
rect 78308 48992 78508 48998
rect 78308 48990 78320 48992
rect 77998 48960 78320 48990
rect 77998 48958 78010 48960
rect 77810 48952 78010 48958
rect 78308 48958 78320 48960
rect 78496 48958 78508 48992
rect 78308 48952 78508 48958
rect 78540 48960 78620 48980
rect 77772 48914 77780 48948
rect 77770 48900 77780 48914
rect 77700 48880 77780 48900
rect 77810 48904 78010 48910
rect 77810 48870 77822 48904
rect 77998 48900 78010 48904
rect 78308 48904 78508 48910
rect 78308 48900 78320 48904
rect 77998 48890 78320 48900
rect 77998 48870 78130 48890
rect 77810 48864 78010 48870
rect 78120 48830 78130 48870
rect 78190 48870 78320 48890
rect 78496 48870 78508 48904
rect 78540 48900 78550 48960
rect 78610 48900 78620 48960
rect 78540 48880 78620 48900
rect 78190 48830 78200 48870
rect 78308 48864 78508 48870
rect 78120 48820 78200 48830
rect 77590 47660 77660 48810
rect 77590 47400 77610 47660
rect 77650 47400 77660 47660
rect 78670 48810 78680 49050
rect 78720 48810 78740 49050
rect 78670 47660 78740 48810
rect 78120 47630 78200 47640
rect 77810 47592 78010 47598
rect 77700 47560 77780 47580
rect 77700 47500 77710 47560
rect 77770 47548 77780 47560
rect 77810 47558 77822 47592
rect 77998 47590 78010 47592
rect 78120 47590 78130 47630
rect 77998 47570 78130 47590
rect 78190 47590 78200 47630
rect 78308 47592 78508 47598
rect 78308 47590 78320 47592
rect 78190 47570 78320 47590
rect 77998 47560 78320 47570
rect 77998 47558 78010 47560
rect 77810 47552 78010 47558
rect 78308 47558 78320 47560
rect 78496 47558 78508 47592
rect 78308 47552 78508 47558
rect 78540 47560 78620 47580
rect 77772 47514 77780 47548
rect 77770 47500 77780 47514
rect 77700 47480 77780 47500
rect 77810 47504 78010 47510
rect 77810 47470 77822 47504
rect 77998 47500 78010 47504
rect 78308 47504 78508 47510
rect 78308 47500 78320 47504
rect 77998 47470 78320 47500
rect 78496 47470 78508 47504
rect 78540 47500 78550 47560
rect 78610 47500 78620 47560
rect 78540 47480 78620 47500
rect 77810 47464 78010 47470
rect 77590 47340 77660 47400
rect 77590 47100 77610 47340
rect 77650 47100 77660 47340
rect 78120 47460 78200 47470
rect 78308 47464 78508 47470
rect 78120 47400 78130 47460
rect 78190 47400 78200 47460
rect 78120 47350 78200 47400
rect 78120 47290 78130 47350
rect 78190 47290 78200 47350
rect 77810 47282 78010 47288
rect 77700 47250 77780 47270
rect 77700 47190 77710 47250
rect 77770 47238 77780 47250
rect 77810 47248 77822 47282
rect 77998 47280 78010 47282
rect 78120 47280 78200 47290
rect 78670 47420 78680 47660
rect 78720 47420 78740 47660
rect 78670 47340 78740 47420
rect 78308 47282 78508 47288
rect 78308 47280 78320 47282
rect 77998 47250 78320 47280
rect 77998 47248 78010 47250
rect 77810 47242 78010 47248
rect 78308 47248 78320 47250
rect 78496 47248 78508 47282
rect 78308 47242 78508 47248
rect 78540 47250 78620 47270
rect 77772 47204 77780 47238
rect 77770 47190 77780 47204
rect 77700 47170 77780 47190
rect 77810 47194 78010 47200
rect 77810 47160 77822 47194
rect 77998 47190 78010 47194
rect 78308 47194 78508 47200
rect 78308 47190 78320 47194
rect 77998 47180 78320 47190
rect 77998 47160 78130 47180
rect 77810 47154 78010 47160
rect 78120 47120 78130 47160
rect 78190 47160 78320 47180
rect 78496 47160 78508 47194
rect 78540 47190 78550 47250
rect 78610 47190 78620 47250
rect 78540 47170 78620 47190
rect 78190 47120 78200 47160
rect 78308 47154 78508 47160
rect 78120 47110 78200 47120
rect 77590 45950 77660 47100
rect 77590 45690 77610 45950
rect 77650 45690 77660 45950
rect 78670 47100 78680 47340
rect 78720 47100 78740 47340
rect 78670 45950 78740 47100
rect 78120 45920 78200 45930
rect 77810 45882 78010 45888
rect 77700 45850 77780 45870
rect 77700 45790 77710 45850
rect 77770 45838 77780 45850
rect 77810 45848 77822 45882
rect 77998 45880 78010 45882
rect 78120 45880 78130 45920
rect 77998 45860 78130 45880
rect 78190 45880 78200 45920
rect 78308 45882 78508 45888
rect 78308 45880 78320 45882
rect 78190 45860 78320 45880
rect 77998 45850 78320 45860
rect 77998 45848 78010 45850
rect 77810 45842 78010 45848
rect 78308 45848 78320 45850
rect 78496 45848 78508 45882
rect 78308 45842 78508 45848
rect 78540 45850 78620 45870
rect 77772 45804 77780 45838
rect 77770 45790 77780 45804
rect 77700 45770 77780 45790
rect 77810 45794 78010 45800
rect 77810 45760 77822 45794
rect 77998 45790 78010 45794
rect 78308 45794 78508 45800
rect 78308 45790 78320 45794
rect 77998 45760 78320 45790
rect 78496 45760 78508 45794
rect 78540 45790 78550 45850
rect 78610 45790 78620 45850
rect 78540 45770 78620 45790
rect 77810 45754 78010 45760
rect 77590 45630 77660 45690
rect 77590 45390 77610 45630
rect 77650 45390 77660 45630
rect 78120 45750 78200 45760
rect 78308 45754 78508 45760
rect 78120 45690 78130 45750
rect 78190 45690 78200 45750
rect 78120 45640 78200 45690
rect 78120 45580 78130 45640
rect 78190 45580 78200 45640
rect 77810 45572 78010 45578
rect 77700 45540 77780 45560
rect 77700 45480 77710 45540
rect 77770 45528 77780 45540
rect 77810 45538 77822 45572
rect 77998 45570 78010 45572
rect 78120 45570 78200 45580
rect 78670 45710 78680 45950
rect 78720 45710 78740 45950
rect 78670 45630 78740 45710
rect 78308 45572 78508 45578
rect 78308 45570 78320 45572
rect 77998 45540 78320 45570
rect 77998 45538 78010 45540
rect 77810 45532 78010 45538
rect 78308 45538 78320 45540
rect 78496 45538 78508 45572
rect 78308 45532 78508 45538
rect 78540 45540 78620 45560
rect 77772 45494 77780 45528
rect 77770 45480 77780 45494
rect 77700 45460 77780 45480
rect 77810 45484 78010 45490
rect 77810 45450 77822 45484
rect 77998 45480 78010 45484
rect 78308 45484 78508 45490
rect 78308 45480 78320 45484
rect 77998 45470 78320 45480
rect 77998 45450 78130 45470
rect 77810 45444 78010 45450
rect 78120 45410 78130 45450
rect 78190 45450 78320 45470
rect 78496 45450 78508 45484
rect 78540 45480 78550 45540
rect 78610 45480 78620 45540
rect 78540 45460 78620 45480
rect 78190 45410 78200 45450
rect 78308 45444 78508 45450
rect 78120 45400 78200 45410
rect 77590 44240 77660 45390
rect 77590 43980 77610 44240
rect 77650 43980 77660 44240
rect 78670 45390 78680 45630
rect 78720 45390 78740 45630
rect 78670 44240 78740 45390
rect 78120 44210 78200 44220
rect 77810 44172 78010 44178
rect 77700 44140 77780 44160
rect 77700 44080 77710 44140
rect 77770 44128 77780 44140
rect 77810 44138 77822 44172
rect 77998 44170 78010 44172
rect 78120 44170 78130 44210
rect 77998 44150 78130 44170
rect 78190 44170 78200 44210
rect 78308 44172 78508 44178
rect 78308 44170 78320 44172
rect 78190 44150 78320 44170
rect 77998 44140 78320 44150
rect 77998 44138 78010 44140
rect 77810 44132 78010 44138
rect 78308 44138 78320 44140
rect 78496 44138 78508 44172
rect 78308 44132 78508 44138
rect 78540 44140 78620 44160
rect 77772 44094 77780 44128
rect 77770 44080 77780 44094
rect 77700 44060 77780 44080
rect 77810 44084 78010 44090
rect 77810 44050 77822 44084
rect 77998 44080 78010 44084
rect 78308 44084 78508 44090
rect 78308 44080 78320 44084
rect 77998 44050 78320 44080
rect 78496 44050 78508 44084
rect 78540 44080 78550 44140
rect 78610 44080 78620 44140
rect 78540 44060 78620 44080
rect 77810 44044 78010 44050
rect 77590 43920 77660 43980
rect 77590 43680 77610 43920
rect 77650 43680 77660 43920
rect 78120 44040 78200 44050
rect 78308 44044 78508 44050
rect 78120 43980 78130 44040
rect 78190 43980 78200 44040
rect 78120 43930 78200 43980
rect 78120 43870 78130 43930
rect 78190 43870 78200 43930
rect 77810 43862 78010 43868
rect 77700 43830 77780 43850
rect 77700 43770 77710 43830
rect 77770 43818 77780 43830
rect 77810 43828 77822 43862
rect 77998 43860 78010 43862
rect 78120 43860 78200 43870
rect 78670 44000 78680 44240
rect 78720 44000 78740 44240
rect 78670 43920 78740 44000
rect 78308 43862 78508 43868
rect 78308 43860 78320 43862
rect 77998 43830 78320 43860
rect 77998 43828 78010 43830
rect 77810 43822 78010 43828
rect 78308 43828 78320 43830
rect 78496 43828 78508 43862
rect 78308 43822 78508 43828
rect 78540 43830 78620 43850
rect 77772 43784 77780 43818
rect 77770 43770 77780 43784
rect 77700 43750 77780 43770
rect 77810 43774 78010 43780
rect 77810 43740 77822 43774
rect 77998 43770 78010 43774
rect 78308 43774 78508 43780
rect 78308 43770 78320 43774
rect 77998 43760 78320 43770
rect 77998 43740 78130 43760
rect 77810 43734 78010 43740
rect 78120 43700 78130 43740
rect 78190 43740 78320 43760
rect 78496 43740 78508 43774
rect 78540 43770 78550 43830
rect 78610 43770 78620 43830
rect 78540 43750 78620 43770
rect 78190 43700 78200 43740
rect 78308 43734 78508 43740
rect 78120 43690 78200 43700
rect 77590 42530 77660 43680
rect 77590 42270 77610 42530
rect 77650 42270 77660 42530
rect 78670 43680 78680 43920
rect 78720 43680 78740 43920
rect 78670 42530 78740 43680
rect 78120 42500 78200 42510
rect 77810 42462 78010 42468
rect 77700 42430 77780 42450
rect 77700 42370 77710 42430
rect 77770 42418 77780 42430
rect 77810 42428 77822 42462
rect 77998 42460 78010 42462
rect 78120 42460 78130 42500
rect 77998 42440 78130 42460
rect 78190 42460 78200 42500
rect 78308 42462 78508 42468
rect 78308 42460 78320 42462
rect 78190 42440 78320 42460
rect 77998 42430 78320 42440
rect 77998 42428 78010 42430
rect 77810 42422 78010 42428
rect 78308 42428 78320 42430
rect 78496 42428 78508 42462
rect 78308 42422 78508 42428
rect 78540 42430 78620 42450
rect 77772 42384 77780 42418
rect 77770 42370 77780 42384
rect 77700 42350 77780 42370
rect 77810 42374 78010 42380
rect 77810 42340 77822 42374
rect 77998 42370 78010 42374
rect 78308 42374 78508 42380
rect 78308 42370 78320 42374
rect 77998 42340 78320 42370
rect 78496 42340 78508 42374
rect 78540 42370 78550 42430
rect 78610 42370 78620 42430
rect 78540 42350 78620 42370
rect 77810 42334 78010 42340
rect 77590 42210 77660 42270
rect 77590 41970 77610 42210
rect 77650 41970 77660 42210
rect 78120 42330 78200 42340
rect 78308 42334 78508 42340
rect 78120 42270 78130 42330
rect 78190 42270 78200 42330
rect 78120 42220 78200 42270
rect 78120 42160 78130 42220
rect 78190 42160 78200 42220
rect 77810 42152 78010 42158
rect 77700 42120 77780 42140
rect 77700 42060 77710 42120
rect 77770 42108 77780 42120
rect 77810 42118 77822 42152
rect 77998 42150 78010 42152
rect 78120 42150 78200 42160
rect 78670 42290 78680 42530
rect 78720 42290 78740 42530
rect 78670 42210 78740 42290
rect 78308 42152 78508 42158
rect 78308 42150 78320 42152
rect 77998 42120 78320 42150
rect 77998 42118 78010 42120
rect 77810 42112 78010 42118
rect 78308 42118 78320 42120
rect 78496 42118 78508 42152
rect 78308 42112 78508 42118
rect 78540 42120 78620 42140
rect 77772 42074 77780 42108
rect 77770 42060 77780 42074
rect 77700 42040 77780 42060
rect 77810 42064 78010 42070
rect 77810 42030 77822 42064
rect 77998 42060 78010 42064
rect 78308 42064 78508 42070
rect 78308 42060 78320 42064
rect 77998 42050 78320 42060
rect 77998 42030 78130 42050
rect 77810 42024 78010 42030
rect 78120 41990 78130 42030
rect 78190 42030 78320 42050
rect 78496 42030 78508 42064
rect 78540 42060 78550 42120
rect 78610 42060 78620 42120
rect 78540 42040 78620 42060
rect 78190 41990 78200 42030
rect 78308 42024 78508 42030
rect 78120 41980 78200 41990
rect 77590 40820 77660 41970
rect 77590 40560 77610 40820
rect 77650 40560 77660 40820
rect 78670 41970 78680 42210
rect 78720 41970 78740 42210
rect 78670 40820 78740 41970
rect 78120 40790 78200 40800
rect 77810 40752 78010 40758
rect 77700 40720 77780 40740
rect 77700 40660 77710 40720
rect 77770 40708 77780 40720
rect 77810 40718 77822 40752
rect 77998 40750 78010 40752
rect 78120 40750 78130 40790
rect 77998 40730 78130 40750
rect 78190 40750 78200 40790
rect 78308 40752 78508 40758
rect 78308 40750 78320 40752
rect 78190 40730 78320 40750
rect 77998 40720 78320 40730
rect 77998 40718 78010 40720
rect 77810 40712 78010 40718
rect 78308 40718 78320 40720
rect 78496 40718 78508 40752
rect 78308 40712 78508 40718
rect 78540 40720 78620 40740
rect 77772 40674 77780 40708
rect 77770 40660 77780 40674
rect 77700 40640 77780 40660
rect 77810 40664 78010 40670
rect 77810 40630 77822 40664
rect 77998 40660 78010 40664
rect 78308 40664 78508 40670
rect 78308 40660 78320 40664
rect 77998 40630 78320 40660
rect 78496 40630 78508 40664
rect 78540 40660 78550 40720
rect 78610 40660 78620 40720
rect 78540 40640 78620 40660
rect 77810 40624 78010 40630
rect 77590 40500 77660 40560
rect 77590 40260 77610 40500
rect 77650 40260 77660 40500
rect 78120 40620 78200 40630
rect 78308 40624 78508 40630
rect 78120 40560 78130 40620
rect 78190 40560 78200 40620
rect 78120 40510 78200 40560
rect 78120 40450 78130 40510
rect 78190 40450 78200 40510
rect 77810 40442 78010 40448
rect 77700 40410 77780 40430
rect 77700 40350 77710 40410
rect 77770 40398 77780 40410
rect 77810 40408 77822 40442
rect 77998 40440 78010 40442
rect 78120 40440 78200 40450
rect 78670 40580 78680 40820
rect 78720 40580 78740 40820
rect 78670 40500 78740 40580
rect 78308 40442 78508 40448
rect 78308 40440 78320 40442
rect 77998 40410 78320 40440
rect 77998 40408 78010 40410
rect 77810 40402 78010 40408
rect 78308 40408 78320 40410
rect 78496 40408 78508 40442
rect 78308 40402 78508 40408
rect 78540 40410 78620 40430
rect 77772 40364 77780 40398
rect 77770 40350 77780 40364
rect 77700 40330 77780 40350
rect 77810 40354 78010 40360
rect 77810 40320 77822 40354
rect 77998 40350 78010 40354
rect 78308 40354 78508 40360
rect 78308 40350 78320 40354
rect 77998 40340 78320 40350
rect 77998 40320 78130 40340
rect 77810 40314 78010 40320
rect 78120 40280 78130 40320
rect 78190 40320 78320 40340
rect 78496 40320 78508 40354
rect 78540 40350 78550 40410
rect 78610 40350 78620 40410
rect 78540 40330 78620 40350
rect 78190 40280 78200 40320
rect 78308 40314 78508 40320
rect 78120 40270 78200 40280
rect 77590 39690 77660 40260
rect 78670 40260 78680 40500
rect 78720 40260 78740 40500
rect 78670 39690 78740 40260
rect 77590 39680 77670 39690
rect 77590 39620 77600 39680
rect 77660 39620 77670 39680
rect 78660 39680 78740 39690
rect 78660 39620 78670 39680
rect 78730 39620 78740 39680
rect 78660 39610 78740 39620
rect 78770 66480 78800 67050
rect 78770 66470 78830 66480
rect 78770 66400 78830 66410
rect 78770 64770 78800 66400
rect 78860 65950 78890 67050
rect 78830 65940 78890 65950
rect 78830 65870 78890 65880
rect 78770 64760 78830 64770
rect 78770 64690 78830 64700
rect 78770 63060 78800 64690
rect 78860 64240 78890 65870
rect 78830 64230 78890 64240
rect 78830 64160 78890 64170
rect 78770 63050 78830 63060
rect 78770 62980 78830 62990
rect 78770 61350 78800 62980
rect 78860 62530 78890 64160
rect 78830 62520 78890 62530
rect 78830 62450 78890 62460
rect 78770 61340 78830 61350
rect 78770 61270 78830 61280
rect 78770 59640 78800 61270
rect 78860 60820 78890 62450
rect 78830 60810 78890 60820
rect 78830 60740 78890 60750
rect 78770 59630 78830 59640
rect 78770 59560 78830 59570
rect 78770 57930 78800 59560
rect 78860 59110 78890 60740
rect 78830 59100 78890 59110
rect 78830 59030 78890 59040
rect 78770 57920 78830 57930
rect 78770 57850 78830 57860
rect 78770 56220 78800 57850
rect 78860 57400 78890 59030
rect 78830 57390 78890 57400
rect 78830 57320 78890 57330
rect 78770 56210 78830 56220
rect 78770 56140 78830 56150
rect 78770 54510 78800 56140
rect 78860 55690 78890 57320
rect 78830 55680 78890 55690
rect 78830 55610 78890 55620
rect 78770 54500 78830 54510
rect 78770 54430 78830 54440
rect 78770 52800 78800 54430
rect 78860 53980 78890 55610
rect 78830 53970 78890 53980
rect 78830 53900 78890 53910
rect 78770 52790 78830 52800
rect 78770 52720 78830 52730
rect 78770 51090 78800 52720
rect 78860 52270 78890 53900
rect 78830 52260 78890 52270
rect 78830 52190 78890 52200
rect 78770 51080 78830 51090
rect 78770 51010 78830 51020
rect 78770 49380 78800 51010
rect 78860 50560 78890 52190
rect 78830 50550 78890 50560
rect 78830 50480 78890 50490
rect 78770 49370 78830 49380
rect 78770 49300 78830 49310
rect 78770 47670 78800 49300
rect 78860 48850 78890 50480
rect 78830 48840 78890 48850
rect 78830 48770 78890 48780
rect 78770 47660 78830 47670
rect 78770 47590 78830 47600
rect 78770 45960 78800 47590
rect 78860 47140 78890 48770
rect 78830 47130 78890 47140
rect 78830 47060 78890 47070
rect 78770 45950 78830 45960
rect 78770 45880 78830 45890
rect 78770 44250 78800 45880
rect 78860 45430 78890 47060
rect 78830 45420 78890 45430
rect 78830 45350 78890 45360
rect 78770 44240 78830 44250
rect 78770 44170 78830 44180
rect 78770 42540 78800 44170
rect 78860 43720 78890 45350
rect 78830 43710 78890 43720
rect 78830 43640 78890 43650
rect 78770 42530 78830 42540
rect 78770 42460 78830 42470
rect 78770 40830 78800 42460
rect 78860 42010 78890 43640
rect 78830 42000 78890 42010
rect 78830 41930 78890 41940
rect 78770 40820 78830 40830
rect 78770 40750 78830 40760
rect 73930 39230 74190 39240
rect 73930 39210 74130 39230
rect 74130 39160 74190 39170
rect 77300 39230 77560 39240
rect 77360 39210 77560 39230
rect 77300 39160 77360 39170
rect 78770 38840 78800 40750
rect 78860 40300 78890 41930
rect 78830 40290 78890 40300
rect 78830 40220 78890 40230
rect 78860 39690 78890 40220
rect 78830 39680 78890 39690
rect 78830 39610 78890 39620
rect 78920 66390 78950 67050
rect 78920 66380 78980 66390
rect 78920 66310 78980 66320
rect 78920 64680 78950 66310
rect 78920 64670 78980 64680
rect 78920 64600 78980 64610
rect 78920 62970 78950 64600
rect 78920 62960 78980 62970
rect 78920 62890 78980 62900
rect 78920 61260 78950 62890
rect 78920 61250 78980 61260
rect 78920 61180 78980 61190
rect 78920 59550 78950 61180
rect 78920 59540 78980 59550
rect 78920 59470 78980 59480
rect 78920 57840 78950 59470
rect 78920 57830 78980 57840
rect 78920 57760 78980 57770
rect 78920 56130 78950 57760
rect 78920 56120 78980 56130
rect 78920 56050 78980 56060
rect 78920 54420 78950 56050
rect 78920 54410 78980 54420
rect 78920 54340 78980 54350
rect 78920 52710 78950 54340
rect 78920 52700 78980 52710
rect 78920 52630 78980 52640
rect 78920 51000 78950 52630
rect 78920 50990 78980 51000
rect 78920 50920 78980 50930
rect 78920 49290 78950 50920
rect 78920 49280 78980 49290
rect 78920 49210 78980 49220
rect 78920 47580 78950 49210
rect 78920 47570 78980 47580
rect 78920 47500 78980 47510
rect 78920 45870 78950 47500
rect 78920 45860 78980 45870
rect 78920 45790 78980 45800
rect 78920 44160 78950 45790
rect 78920 44150 78980 44160
rect 78920 44080 78980 44090
rect 78920 42450 78950 44080
rect 78920 42440 78980 42450
rect 78920 42370 78980 42380
rect 78920 40740 78950 42370
rect 78920 40730 78980 40740
rect 78920 40660 78980 40670
rect 78920 39240 78950 40660
rect 79040 39690 79070 67050
rect 79160 39690 79190 67050
rect 79280 39690 79310 67050
rect 79400 39690 79430 67050
rect 79520 39690 79550 67050
rect 79640 39690 79670 67050
rect 78920 39230 79180 39240
rect 78920 39210 79120 39230
rect 79120 39160 79180 39170
rect 40 38810 79800 38840
rect 40 38670 3970 38700
rect 3960 38640 3970 38670
rect 4030 38670 8960 38700
rect 4030 38640 4040 38670
rect 8950 38640 8960 38670
rect 9020 38670 13950 38700
rect 9020 38640 9030 38670
rect 13940 38640 13950 38670
rect 14010 38670 18940 38700
rect 14010 38640 14020 38670
rect 18930 38640 18940 38670
rect 19000 38670 23930 38700
rect 19000 38640 19010 38670
rect 23920 38640 23930 38670
rect 23990 38670 28920 38700
rect 23990 38640 24000 38670
rect 28910 38640 28920 38670
rect 28980 38670 33910 38700
rect 28980 38640 28990 38670
rect 33900 38640 33910 38670
rect 33970 38670 38900 38700
rect 33970 38640 33980 38670
rect 38890 38640 38900 38670
rect 38960 38670 43890 38700
rect 38960 38640 38970 38670
rect 43880 38640 43890 38670
rect 43950 38670 48880 38700
rect 43950 38640 43960 38670
rect 48870 38640 48880 38670
rect 48940 38670 53870 38700
rect 48940 38640 48950 38670
rect 53860 38640 53870 38670
rect 53930 38670 58860 38700
rect 53930 38640 53940 38670
rect 58850 38640 58860 38670
rect 58920 38670 63850 38700
rect 58920 38640 58930 38670
rect 63840 38640 63850 38670
rect 63910 38670 68840 38700
rect 63910 38640 63920 38670
rect 68830 38640 68840 38670
rect 68900 38670 73830 38700
rect 68900 38640 68910 38670
rect 73820 38640 73830 38670
rect 73890 38670 78820 38700
rect 73890 38640 73900 38670
rect 78810 38640 78820 38670
rect 78880 38670 79800 38700
rect 78880 38640 78890 38670
rect 40 38530 40200 38560
rect 36370 38490 36430 38530
rect 40190 38500 40200 38530
rect 40260 38530 79800 38560
rect 40260 38500 40270 38530
rect 40 38390 40270 38420
rect 36310 38350 36370 38390
rect 40260 38360 40270 38390
rect 40330 38390 79800 38420
rect 40330 38360 40340 38390
rect 40 38250 45020 38280
rect 45010 38220 45020 38250
rect 45080 38250 79800 38280
rect 45080 38220 45090 38250
rect 40 38110 45110 38140
rect 45100 38080 45110 38110
rect 45170 38110 79800 38140
rect 45170 38080 45180 38110
rect 40 37970 40030 38000
rect 36550 37930 36610 37970
rect 40020 37940 40030 37970
rect 40090 37970 45200 38000
rect 40090 37940 40100 37970
rect 45190 37940 45200 37970
rect 45260 37970 79800 38000
rect 45260 37940 45270 37970
rect 40 37830 40090 37860
rect 40080 37800 40090 37830
rect 40150 37830 45260 37860
rect 40150 37800 40160 37830
rect 45250 37800 45260 37830
rect 45320 37830 79800 37860
rect 45320 37800 45330 37830
rect 40 37690 34860 37720
rect 31740 37650 31800 37690
rect 34850 37660 34860 37690
rect 34920 37690 49830 37720
rect 34920 37660 34930 37690
rect 46710 37650 46770 37690
rect 49820 37660 49830 37690
rect 49890 37690 79800 37720
rect 49890 37660 49900 37690
rect 40 37550 34920 37580
rect 34910 37520 34920 37550
rect 34980 37550 49890 37580
rect 34980 37520 34990 37550
rect 49880 37520 49890 37550
rect 49950 37550 79800 37580
rect 49950 37520 49960 37550
rect 40 37410 35040 37440
rect 31560 37370 31620 37410
rect 35030 37380 35040 37410
rect 35100 37410 39850 37440
rect 35100 37380 35110 37410
rect 36730 37370 36790 37410
rect 39840 37380 39850 37410
rect 39910 37410 44840 37440
rect 39910 37380 39920 37410
rect 41720 37370 41780 37410
rect 44830 37380 44840 37410
rect 44900 37410 50010 37440
rect 44900 37380 44910 37410
rect 46530 37370 46590 37410
rect 50000 37380 50010 37410
rect 50070 37410 79800 37440
rect 50070 37380 50080 37410
rect 40 37270 35100 37300
rect 35090 37240 35100 37270
rect 35160 37270 39910 37300
rect 35160 37240 35170 37270
rect 39900 37240 39910 37270
rect 39970 37270 44900 37300
rect 39970 37240 39980 37270
rect 44890 37240 44900 37270
rect 44960 37270 50070 37300
rect 44960 37240 44970 37270
rect 50060 37240 50070 37270
rect 50130 37270 79800 37300
rect 50130 37240 50140 37270
rect 40 37130 24520 37160
rect 22120 37090 22180 37130
rect 24510 37100 24520 37130
rect 24580 37130 29510 37160
rect 24580 37100 24590 37130
rect 27110 37090 27170 37130
rect 29500 37100 29510 37130
rect 29570 37130 34680 37160
rect 29570 37100 29580 37130
rect 31920 37090 31980 37130
rect 34670 37100 34680 37130
rect 34740 37130 39670 37160
rect 34740 37100 34750 37130
rect 36910 37090 36970 37130
rect 39660 37100 39670 37130
rect 39730 37130 44660 37160
rect 39730 37100 39740 37130
rect 41900 37090 41960 37130
rect 44650 37100 44660 37130
rect 44720 37130 49650 37160
rect 44720 37100 44730 37130
rect 46890 37090 46950 37130
rect 49640 37100 49650 37130
rect 49710 37130 54460 37160
rect 49710 37100 49720 37130
rect 52060 37090 52120 37130
rect 54450 37100 54460 37130
rect 54520 37130 59450 37160
rect 54520 37100 54530 37130
rect 57050 37090 57110 37130
rect 59440 37100 59450 37130
rect 59510 37130 79800 37160
rect 59510 37100 59520 37130
rect 40 36990 24580 37020
rect 24570 36960 24580 36990
rect 24640 36990 29570 37020
rect 24640 36960 24650 36990
rect 29560 36960 29570 36990
rect 29630 36990 34740 37020
rect 29630 36960 29640 36990
rect 34730 36960 34740 36990
rect 34800 36990 39730 37020
rect 34800 36960 34810 36990
rect 39720 36960 39730 36990
rect 39790 36990 44720 37020
rect 39790 36960 39800 36990
rect 44710 36960 44720 36990
rect 44780 36990 49710 37020
rect 44780 36960 44790 36990
rect 49700 36960 49710 36990
rect 49770 36990 54520 37020
rect 49770 36960 49780 36990
rect 54510 36960 54520 36990
rect 54580 36990 59510 37020
rect 54580 36960 54590 36990
rect 59500 36960 59510 36990
rect 59570 36990 79800 37020
rect 59570 36960 59580 36990
rect 40 36850 24700 36880
rect 21940 36810 22000 36850
rect 24690 36820 24700 36850
rect 24760 36850 29690 36880
rect 24760 36820 24770 36850
rect 26930 36810 26990 36850
rect 29680 36820 29690 36850
rect 29750 36850 34500 36880
rect 29750 36820 29760 36850
rect 32100 36810 32160 36850
rect 34490 36820 34500 36850
rect 34560 36850 39490 36880
rect 34560 36820 34570 36850
rect 37090 36810 37150 36850
rect 39480 36820 39490 36850
rect 39550 36850 44480 36880
rect 39550 36820 39560 36850
rect 42080 36810 42140 36850
rect 44470 36820 44480 36850
rect 44540 36850 49470 36880
rect 44540 36820 44550 36850
rect 47070 36810 47130 36850
rect 49460 36820 49470 36850
rect 49530 36850 54640 36880
rect 49530 36820 49540 36850
rect 51880 36810 51940 36850
rect 54630 36820 54640 36850
rect 54700 36850 59630 36880
rect 54700 36820 54710 36850
rect 56870 36810 56930 36850
rect 59620 36820 59630 36850
rect 59690 36850 79800 36880
rect 59690 36820 59700 36850
rect 40 36710 24760 36740
rect 24750 36680 24760 36710
rect 24820 36710 29750 36740
rect 24820 36680 24830 36710
rect 29740 36680 29750 36710
rect 29810 36710 34560 36740
rect 29810 36680 29820 36710
rect 34550 36680 34560 36710
rect 34620 36710 39550 36740
rect 34620 36680 34630 36710
rect 39540 36680 39550 36710
rect 39610 36710 44540 36740
rect 39610 36680 39620 36710
rect 44530 36680 44540 36710
rect 44600 36710 49530 36740
rect 44600 36680 44610 36710
rect 49520 36680 49530 36710
rect 49590 36710 54700 36740
rect 49590 36680 49600 36710
rect 54690 36680 54700 36710
rect 54760 36710 59690 36740
rect 54760 36680 54770 36710
rect 59680 36680 59690 36710
rect 59750 36710 79800 36740
rect 59750 36680 59760 36710
rect 40 36570 14360 36600
rect 12320 36530 12380 36570
rect 14350 36540 14360 36570
rect 14420 36570 19350 36600
rect 14420 36540 14430 36570
rect 17310 36530 17370 36570
rect 19340 36540 19350 36570
rect 19410 36570 24340 36600
rect 19410 36540 19420 36570
rect 22300 36530 22360 36570
rect 24330 36540 24340 36570
rect 24400 36570 29330 36600
rect 24400 36540 24410 36570
rect 27290 36530 27350 36570
rect 29320 36540 29330 36570
rect 29390 36570 34320 36600
rect 29390 36540 29400 36570
rect 32280 36530 32340 36570
rect 34310 36540 34320 36570
rect 34380 36570 39310 36600
rect 34380 36540 34390 36570
rect 37270 36530 37330 36570
rect 39300 36540 39310 36570
rect 39370 36570 44300 36600
rect 39370 36540 39380 36570
rect 42260 36530 42320 36570
rect 44290 36540 44300 36570
rect 44360 36570 49290 36600
rect 44360 36540 44370 36570
rect 47250 36530 47310 36570
rect 49280 36540 49290 36570
rect 49350 36570 54280 36600
rect 49350 36540 49360 36570
rect 52240 36530 52300 36570
rect 54270 36540 54280 36570
rect 54340 36570 59270 36600
rect 54340 36540 54350 36570
rect 57230 36530 57290 36570
rect 59260 36540 59270 36570
rect 59330 36570 64260 36600
rect 59330 36540 59340 36570
rect 62220 36530 62280 36570
rect 64250 36540 64260 36570
rect 64320 36570 69250 36600
rect 64320 36540 64330 36570
rect 67210 36530 67270 36570
rect 69240 36540 69250 36570
rect 69310 36570 79800 36600
rect 69310 36540 69320 36570
rect 40 36430 14420 36460
rect 14410 36400 14420 36430
rect 14480 36430 19410 36460
rect 14480 36400 14490 36430
rect 19400 36400 19410 36430
rect 19470 36430 24400 36460
rect 19470 36400 19480 36430
rect 24390 36400 24400 36430
rect 24460 36430 29390 36460
rect 24460 36400 24470 36430
rect 29380 36400 29390 36430
rect 29450 36430 34380 36460
rect 29450 36400 29460 36430
rect 34370 36400 34380 36430
rect 34440 36430 39370 36460
rect 34440 36400 34450 36430
rect 39360 36400 39370 36430
rect 39430 36430 44360 36460
rect 39430 36400 39440 36430
rect 44350 36400 44360 36430
rect 44420 36430 49350 36460
rect 44420 36400 44430 36430
rect 49340 36400 49350 36430
rect 49410 36430 54340 36460
rect 49410 36400 49420 36430
rect 54330 36400 54340 36430
rect 54400 36430 59330 36460
rect 54400 36400 54410 36430
rect 59320 36400 59330 36430
rect 59390 36430 64320 36460
rect 59390 36400 59400 36430
rect 64310 36400 64320 36430
rect 64380 36430 69310 36460
rect 64380 36400 64390 36430
rect 69300 36400 69310 36430
rect 69370 36430 79800 36460
rect 69370 36400 69380 36430
rect 40 36290 4200 36320
rect 2520 36250 2580 36290
rect 4190 36260 4200 36290
rect 4260 36290 9190 36320
rect 4260 36260 4270 36290
rect 7510 36250 7570 36290
rect 9180 36260 9190 36290
rect 9250 36290 14180 36320
rect 9250 36260 9260 36290
rect 12500 36250 12560 36290
rect 14170 36260 14180 36290
rect 14240 36290 19170 36320
rect 14240 36260 14250 36290
rect 17490 36250 17550 36290
rect 19160 36260 19170 36290
rect 19230 36290 24160 36320
rect 19230 36260 19240 36290
rect 22480 36250 22540 36290
rect 24150 36260 24160 36290
rect 24220 36290 29150 36320
rect 24220 36260 24230 36290
rect 27470 36250 27530 36290
rect 29140 36260 29150 36290
rect 29210 36290 34140 36320
rect 29210 36260 29220 36290
rect 32460 36250 32520 36290
rect 34130 36260 34140 36290
rect 34200 36290 39130 36320
rect 34200 36260 34210 36290
rect 37450 36250 37510 36290
rect 39120 36260 39130 36290
rect 39190 36290 44120 36320
rect 39190 36260 39200 36290
rect 42440 36250 42500 36290
rect 44110 36260 44120 36290
rect 44180 36290 49110 36320
rect 44180 36260 44190 36290
rect 47430 36250 47490 36290
rect 49100 36260 49110 36290
rect 49170 36290 54100 36320
rect 49170 36260 49180 36290
rect 52420 36250 52480 36290
rect 54090 36260 54100 36290
rect 54160 36290 59090 36320
rect 54160 36260 54170 36290
rect 57410 36250 57470 36290
rect 59080 36260 59090 36290
rect 59150 36290 64080 36320
rect 59150 36260 59160 36290
rect 62400 36250 62460 36290
rect 64070 36260 64080 36290
rect 64140 36290 69070 36320
rect 64140 36260 64150 36290
rect 67390 36250 67450 36290
rect 69060 36260 69070 36290
rect 69130 36290 74060 36320
rect 69130 36260 69140 36290
rect 72380 36250 72440 36290
rect 74050 36260 74060 36290
rect 74120 36290 79050 36320
rect 74120 36260 74130 36290
rect 77370 36250 77430 36290
rect 79040 36260 79050 36290
rect 79110 36290 79800 36320
rect 79110 36260 79120 36290
rect 40 36150 4260 36180
rect 4250 36120 4260 36150
rect 4320 36150 9250 36180
rect 4320 36120 4330 36150
rect 9240 36120 9250 36150
rect 9310 36150 14240 36180
rect 9310 36120 9320 36150
rect 14230 36120 14240 36150
rect 14300 36150 19230 36180
rect 14300 36120 14310 36150
rect 19220 36120 19230 36150
rect 19290 36150 24220 36180
rect 19290 36120 19300 36150
rect 24210 36120 24220 36150
rect 24280 36150 29210 36180
rect 24280 36120 24290 36150
rect 29200 36120 29210 36150
rect 29270 36150 34200 36180
rect 29270 36120 29280 36150
rect 34190 36120 34200 36150
rect 34260 36150 39190 36180
rect 34260 36120 34270 36150
rect 39180 36120 39190 36150
rect 39250 36150 44180 36180
rect 39250 36120 39260 36150
rect 44170 36120 44180 36150
rect 44240 36150 49170 36180
rect 44240 36120 44250 36150
rect 49160 36120 49170 36150
rect 49230 36150 54160 36180
rect 49230 36120 49240 36150
rect 54150 36120 54160 36150
rect 54220 36150 59150 36180
rect 54220 36120 54230 36150
rect 59140 36120 59150 36150
rect 59210 36150 64140 36180
rect 59210 36120 59220 36150
rect 64130 36120 64140 36150
rect 64200 36150 69130 36180
rect 64200 36120 64210 36150
rect 69120 36120 69130 36150
rect 69190 36150 74120 36180
rect 69190 36120 69200 36150
rect 74110 36120 74120 36150
rect 74180 36150 79110 36180
rect 74180 36120 74190 36150
rect 79100 36120 79110 36150
rect 79170 36150 79800 36180
rect 79170 36120 79180 36150
rect 4150 30900 4160 30930
rect -60 30870 4160 30900
rect 4220 30900 4230 30930
rect 9140 30900 9150 30930
rect 4220 30870 9150 30900
rect 9210 30900 9220 30930
rect 14130 30900 14140 30930
rect 9210 30870 14140 30900
rect 14200 30900 14210 30930
rect 19120 30900 19130 30930
rect 14200 30870 19130 30900
rect 19190 30900 19200 30930
rect 24110 30900 24120 30930
rect 19190 30870 24120 30900
rect 24180 30900 24190 30930
rect 29100 30900 29110 30930
rect 24180 30870 29110 30900
rect 29170 30900 29180 30930
rect 34090 30900 34100 30930
rect 29170 30870 34100 30900
rect 34160 30900 34170 30930
rect 39080 30900 39090 30930
rect 34160 30870 39090 30900
rect 39150 30900 39160 30930
rect 44070 30900 44080 30930
rect 39150 30870 44080 30900
rect 44140 30900 44150 30930
rect 49060 30900 49070 30930
rect 44140 30870 49070 30900
rect 49130 30900 49140 30930
rect 54050 30900 54060 30930
rect 49130 30870 54060 30900
rect 54120 30900 54130 30930
rect 59040 30900 59050 30930
rect 54120 30870 59050 30900
rect 59110 30900 59120 30930
rect 64030 30900 64040 30930
rect 59110 30870 64040 30900
rect 64100 30900 64110 30930
rect 69020 30900 69030 30930
rect 64100 30870 69030 30900
rect 69090 30900 69100 30930
rect 74010 30900 74020 30930
rect 69090 30870 74020 30900
rect 74080 30900 74090 30930
rect 79000 30900 79010 30930
rect 74080 30870 79010 30900
rect 79070 30900 79080 30930
rect 79070 30870 79700 30900
rect 2420 30760 2480 30800
rect 4090 30760 4100 30790
rect -60 30730 4100 30760
rect 4160 30760 4170 30790
rect 7410 30760 7470 30800
rect 9080 30760 9090 30790
rect 4160 30730 9090 30760
rect 9150 30760 9160 30790
rect 12400 30760 12460 30800
rect 14070 30760 14080 30790
rect 9150 30730 14080 30760
rect 14140 30760 14150 30790
rect 17390 30760 17450 30800
rect 19060 30760 19070 30790
rect 14140 30730 19070 30760
rect 19130 30760 19140 30790
rect 22380 30760 22440 30800
rect 24050 30760 24060 30790
rect 19130 30730 24060 30760
rect 24120 30760 24130 30790
rect 27370 30760 27430 30800
rect 29040 30760 29050 30790
rect 24120 30730 29050 30760
rect 29110 30760 29120 30790
rect 32360 30760 32420 30800
rect 34030 30760 34040 30790
rect 29110 30730 34040 30760
rect 34100 30760 34110 30790
rect 37350 30760 37410 30800
rect 39020 30760 39030 30790
rect 34100 30730 39030 30760
rect 39090 30760 39100 30790
rect 42340 30760 42400 30800
rect 44010 30760 44020 30790
rect 39090 30730 44020 30760
rect 44080 30760 44090 30790
rect 47330 30760 47390 30800
rect 49000 30760 49010 30790
rect 44080 30730 49010 30760
rect 49070 30760 49080 30790
rect 52320 30760 52380 30800
rect 53990 30760 54000 30790
rect 49070 30730 54000 30760
rect 54060 30760 54070 30790
rect 57310 30760 57370 30800
rect 58980 30760 58990 30790
rect 54060 30730 58990 30760
rect 59050 30760 59060 30790
rect 62300 30760 62360 30800
rect 63970 30760 63980 30790
rect 59050 30730 63980 30760
rect 64040 30760 64050 30790
rect 67290 30760 67350 30800
rect 68960 30760 68970 30790
rect 64040 30730 68970 30760
rect 69030 30760 69040 30790
rect 72280 30760 72340 30800
rect 73950 30760 73960 30790
rect 69030 30730 73960 30760
rect 74020 30760 74030 30790
rect 77270 30760 77330 30800
rect 78940 30760 78950 30790
rect 74020 30730 78950 30760
rect 79010 30760 79020 30790
rect 79010 30730 79700 30760
rect -9652 12618 -1736 30652
rect 14310 30620 14320 30650
rect -60 30590 14320 30620
rect 14380 30620 14390 30650
rect 19300 30620 19310 30650
rect 14380 30590 19310 30620
rect 19370 30620 19380 30650
rect 24290 30620 24300 30650
rect 19370 30590 24300 30620
rect 24360 30620 24370 30650
rect 29280 30620 29290 30650
rect 24360 30590 29290 30620
rect 29350 30620 29360 30650
rect 34270 30620 34280 30650
rect 29350 30590 34280 30620
rect 34340 30620 34350 30650
rect 39260 30620 39270 30650
rect 34340 30590 39270 30620
rect 39330 30620 39340 30650
rect 44250 30620 44260 30650
rect 39330 30590 44260 30620
rect 44320 30620 44330 30650
rect 49240 30620 49250 30650
rect 44320 30590 49250 30620
rect 49310 30620 49320 30650
rect 54230 30620 54240 30650
rect 49310 30590 54240 30620
rect 54300 30620 54310 30650
rect 59220 30620 59230 30650
rect 54300 30590 59230 30620
rect 59290 30620 59300 30650
rect 64210 30620 64220 30650
rect 59290 30590 64220 30620
rect 64280 30620 64290 30650
rect 69200 30620 69210 30650
rect 64280 30590 69210 30620
rect 69270 30620 69280 30650
rect 69270 30590 79700 30620
rect 12220 30480 12280 30520
rect 14250 30480 14260 30510
rect -60 30450 14260 30480
rect 14320 30480 14330 30510
rect 17210 30480 17270 30520
rect 19240 30480 19250 30510
rect 14320 30450 19250 30480
rect 19310 30480 19320 30510
rect 22200 30480 22260 30520
rect 24230 30480 24240 30510
rect 19310 30450 24240 30480
rect 24300 30480 24310 30510
rect 27190 30480 27250 30520
rect 29220 30480 29230 30510
rect 24300 30450 29230 30480
rect 29290 30480 29300 30510
rect 32180 30480 32240 30520
rect 34210 30480 34220 30510
rect 29290 30450 34220 30480
rect 34280 30480 34290 30510
rect 37170 30480 37230 30520
rect 39200 30480 39210 30510
rect 34280 30450 39210 30480
rect 39270 30480 39280 30510
rect 42160 30480 42220 30520
rect 44190 30480 44200 30510
rect 39270 30450 44200 30480
rect 44260 30480 44270 30510
rect 47150 30480 47210 30520
rect 49180 30480 49190 30510
rect 44260 30450 49190 30480
rect 49250 30480 49260 30510
rect 52140 30480 52200 30520
rect 54170 30480 54180 30510
rect 49250 30450 54180 30480
rect 54240 30480 54250 30510
rect 57130 30480 57190 30520
rect 59160 30480 59170 30510
rect 54240 30450 59170 30480
rect 59230 30480 59240 30510
rect 62120 30480 62180 30520
rect 64150 30480 64160 30510
rect 59230 30450 64160 30480
rect 64220 30480 64230 30510
rect 67110 30480 67170 30520
rect 69140 30480 69150 30510
rect 64220 30450 69150 30480
rect 69210 30480 69220 30510
rect 69210 30450 79700 30480
rect 24650 30340 24660 30370
rect -60 30310 24660 30340
rect 24720 30340 24730 30370
rect 29640 30340 29650 30370
rect 24720 30310 29650 30340
rect 29710 30340 29720 30370
rect 34450 30340 34460 30370
rect 29710 30310 34460 30340
rect 34520 30340 34530 30370
rect 39440 30340 39450 30370
rect 34520 30310 39450 30340
rect 39510 30340 39520 30370
rect 44430 30340 44440 30370
rect 39510 30310 44440 30340
rect 44500 30340 44510 30370
rect 49420 30340 49430 30370
rect 44500 30310 49430 30340
rect 49490 30340 49500 30370
rect 54590 30340 54600 30370
rect 49490 30310 54600 30340
rect 54660 30340 54670 30370
rect 59580 30340 59590 30370
rect 54660 30310 59590 30340
rect 59650 30340 59660 30370
rect 59650 30310 79700 30340
rect 21840 30200 21900 30240
rect 24590 30200 24600 30230
rect -60 30170 24600 30200
rect 24660 30200 24670 30230
rect 26830 30200 26890 30240
rect 29580 30200 29590 30230
rect 24660 30170 29590 30200
rect 29650 30200 29660 30230
rect 32000 30200 32060 30240
rect 34390 30200 34400 30230
rect 29650 30170 34400 30200
rect 34460 30200 34470 30230
rect 36990 30200 37050 30240
rect 39380 30200 39390 30230
rect 34460 30170 39390 30200
rect 39450 30200 39460 30230
rect 41980 30200 42040 30240
rect 44370 30200 44380 30230
rect 39450 30170 44380 30200
rect 44440 30200 44450 30230
rect 46970 30200 47030 30240
rect 49360 30200 49370 30230
rect 44440 30170 49370 30200
rect 49430 30200 49440 30230
rect 51780 30200 51840 30240
rect 54530 30200 54540 30230
rect 49430 30170 54540 30200
rect 54600 30200 54610 30230
rect 56770 30200 56830 30240
rect 59520 30200 59530 30230
rect 54600 30170 59530 30200
rect 59590 30200 59600 30230
rect 59590 30170 79700 30200
rect 24470 30060 24480 30090
rect -60 30030 24480 30060
rect 24540 30060 24550 30090
rect 29460 30060 29470 30090
rect 24540 30030 29470 30060
rect 29530 30060 29540 30090
rect 34630 30060 34640 30090
rect 29530 30030 34640 30060
rect 34700 30060 34710 30090
rect 39620 30060 39630 30090
rect 34700 30030 39630 30060
rect 39690 30060 39700 30090
rect 44610 30060 44620 30090
rect 39690 30030 44620 30060
rect 44680 30060 44690 30090
rect 49600 30060 49610 30090
rect 44680 30030 49610 30060
rect 49670 30060 49680 30090
rect 54410 30060 54420 30090
rect 49670 30030 54420 30060
rect 54480 30060 54490 30090
rect 59400 30060 59410 30090
rect 54480 30030 59410 30060
rect 59470 30060 59480 30090
rect 59470 30030 79700 30060
rect 22020 29920 22080 29960
rect 24410 29920 24420 29950
rect -60 29890 24420 29920
rect 24480 29920 24490 29950
rect 27010 29920 27070 29960
rect 29400 29920 29410 29950
rect 24480 29890 29410 29920
rect 29470 29920 29480 29950
rect 31820 29920 31880 29960
rect 34570 29920 34580 29950
rect 29470 29890 34580 29920
rect 34640 29920 34650 29950
rect 36810 29920 36870 29960
rect 39560 29920 39570 29950
rect 34640 29890 39570 29920
rect 39630 29920 39640 29950
rect 41800 29920 41860 29960
rect 44550 29920 44560 29950
rect 39630 29890 44560 29920
rect 44620 29920 44630 29950
rect 46790 29920 46850 29960
rect 49540 29920 49550 29950
rect 44620 29890 49550 29920
rect 49610 29920 49620 29950
rect 51960 29920 52020 29960
rect 54350 29920 54360 29950
rect 49610 29890 54360 29920
rect 54420 29920 54430 29950
rect 56950 29920 57010 29960
rect 59340 29920 59350 29950
rect 54420 29890 59350 29920
rect 59410 29920 59420 29950
rect 59410 29890 79700 29920
rect 34990 29780 35000 29810
rect -60 29750 35000 29780
rect 35060 29780 35070 29810
rect 39800 29780 39810 29810
rect 35060 29750 39810 29780
rect 39870 29780 39880 29810
rect 44790 29780 44800 29810
rect 39870 29750 44800 29780
rect 44860 29780 44870 29810
rect 49960 29780 49970 29810
rect 44860 29750 49970 29780
rect 50030 29780 50040 29810
rect 50030 29750 79700 29780
rect 31460 29640 31520 29680
rect 34930 29640 34940 29670
rect -60 29610 34940 29640
rect 35000 29640 35010 29670
rect 36630 29640 36690 29680
rect 39740 29640 39750 29670
rect 35000 29610 39750 29640
rect 39810 29640 39820 29670
rect 41620 29640 41680 29680
rect 44730 29640 44740 29670
rect 39810 29610 44740 29640
rect 44800 29640 44810 29670
rect 46430 29640 46490 29680
rect 49900 29640 49910 29670
rect 44800 29610 49910 29640
rect 49970 29640 49980 29670
rect 49970 29610 79700 29640
rect 34810 29500 34820 29530
rect -60 29470 34820 29500
rect 34880 29500 34890 29530
rect 49780 29500 49790 29530
rect 34880 29470 49790 29500
rect 49850 29500 49860 29530
rect 49850 29470 79700 29500
rect 31640 29360 31700 29400
rect 34750 29360 34760 29390
rect -60 29330 34760 29360
rect 34820 29360 34830 29390
rect 46610 29360 46670 29400
rect 49720 29360 49730 29390
rect 34820 29330 49730 29360
rect 49790 29360 49800 29390
rect 49790 29330 79700 29360
rect 39980 29220 39990 29250
rect -60 29190 39990 29220
rect 40050 29220 40060 29250
rect 45150 29220 45160 29250
rect 40050 29190 45160 29220
rect 45220 29220 45230 29250
rect 45220 29190 79700 29220
rect 36450 29080 36510 29120
rect 39920 29080 39930 29110
rect -60 29050 39930 29080
rect 39990 29080 40000 29110
rect 45090 29080 45100 29110
rect 39990 29050 45100 29080
rect 45160 29080 45170 29110
rect 45160 29050 79700 29080
rect 45000 28940 45010 28970
rect -60 28910 45010 28940
rect 45070 28940 45080 28970
rect 45070 28910 79700 28940
rect 44910 28800 44920 28830
rect -60 28770 44920 28800
rect 44980 28800 44990 28830
rect 44980 28770 79700 28800
rect 36210 28660 36270 28700
rect 40160 28660 40170 28690
rect -60 28630 40170 28660
rect 40230 28660 40240 28690
rect 40230 28630 79700 28660
rect 36270 28520 36330 28560
rect 40090 28520 40100 28550
rect -60 28490 40100 28520
rect 40160 28520 40170 28550
rect 40160 28490 79700 28520
rect -58 28420 3872 28450
rect 3860 28380 3870 28410
rect -60 28350 3870 28380
rect 3930 28380 3940 28410
rect 8850 28380 8860 28410
rect 3930 28350 8860 28380
rect 8920 28380 8930 28410
rect 13840 28380 13850 28410
rect 8920 28350 13850 28380
rect 13910 28380 13920 28410
rect 18830 28380 18840 28410
rect 13910 28350 18840 28380
rect 18900 28380 18910 28410
rect 23820 28380 23830 28410
rect 18900 28350 23830 28380
rect 23890 28380 23900 28410
rect 28810 28380 28820 28410
rect 23890 28350 28820 28380
rect 28880 28380 28890 28410
rect 33800 28380 33810 28410
rect 28880 28350 33810 28380
rect 33870 28380 33880 28410
rect 38790 28380 38800 28410
rect 33870 28350 38800 28380
rect 38860 28380 38870 28410
rect 43780 28380 43790 28410
rect 38860 28350 43790 28380
rect 43850 28380 43860 28410
rect 48770 28380 48780 28410
rect 43850 28350 48780 28380
rect 48840 28380 48850 28410
rect 53760 28380 53770 28410
rect 48840 28350 53770 28380
rect 53830 28380 53840 28410
rect 58750 28380 58760 28410
rect 53830 28350 58760 28380
rect 58820 28380 58830 28410
rect 63740 28380 63750 28410
rect 58820 28350 63750 28380
rect 63810 28380 63820 28410
rect 68730 28380 68740 28410
rect 63810 28350 68740 28380
rect 68800 28380 68810 28410
rect 73720 28380 73730 28410
rect 68800 28350 73730 28380
rect 73790 28380 73800 28410
rect 78710 28380 78720 28410
rect 73790 28350 78720 28380
rect 78780 28380 78790 28410
rect 78780 28350 79700 28380
rect -60 28210 79700 28240
rect 2350 27880 2410 27890
rect 2410 27820 2610 27840
rect 2350 27810 2610 27820
rect 2580 27360 2610 27810
rect 3710 27430 3790 27440
rect 2640 27370 2650 27430
rect 2710 27370 2720 27430
rect 2640 27360 2720 27370
rect 3710 27370 3720 27430
rect 3780 27370 3790 27430
rect 3710 27360 3790 27370
rect 3820 27360 3850 28210
rect 4170 27880 4230 27890
rect 3970 27820 4170 27840
rect 3970 27810 4230 27820
rect 7340 27880 7400 27890
rect 7400 27820 7600 27840
rect 7340 27810 7600 27820
rect 3880 27430 3940 27440
rect 3880 27360 3940 27370
rect 3970 27360 4000 27810
rect 7570 27360 7600 27810
rect 8700 27430 8780 27440
rect 7630 27370 7640 27430
rect 7700 27370 7710 27430
rect 7630 27360 7710 27370
rect 8700 27370 8710 27430
rect 8770 27370 8780 27430
rect 8700 27360 8780 27370
rect 8810 27360 8840 28210
rect 9160 27880 9220 27890
rect 8960 27820 9160 27840
rect 12330 27880 12390 27890
rect 8960 27810 9220 27820
rect 12150 27820 12210 27830
rect 8870 27430 8930 27440
rect 8870 27360 8930 27370
rect 8960 27360 8990 27810
rect 12390 27820 12590 27840
rect 12330 27810 12590 27820
rect 12210 27760 12470 27780
rect 12150 27750 12470 27760
rect 12440 27360 12470 27750
rect 12560 27360 12590 27810
rect 13690 27430 13770 27440
rect 12620 27370 12630 27430
rect 12690 27370 12700 27430
rect 12620 27360 12700 27370
rect 13690 27370 13700 27430
rect 13760 27370 13770 27430
rect 13690 27360 13770 27370
rect 13800 27360 13830 28210
rect 14150 27880 14210 27890
rect 13950 27820 14150 27840
rect 17320 27880 17380 27890
rect 13950 27810 14210 27820
rect 14330 27820 14390 27830
rect 13860 27430 13920 27440
rect 13860 27360 13920 27370
rect 13950 27360 13980 27810
rect 14070 27760 14330 27780
rect 14070 27750 14390 27760
rect 17140 27820 17200 27830
rect 17380 27820 17580 27840
rect 17320 27810 17580 27820
rect 17200 27760 17460 27780
rect 17140 27750 17460 27760
rect 14070 27360 14100 27750
rect 17430 27360 17460 27750
rect 17550 27360 17580 27810
rect 18680 27430 18760 27440
rect 17610 27370 17620 27430
rect 17680 27370 17690 27430
rect 17610 27360 17690 27370
rect 18680 27370 18690 27430
rect 18750 27370 18760 27430
rect 18680 27360 18760 27370
rect 18790 27360 18820 28210
rect 19140 27880 19200 27890
rect 18940 27820 19140 27840
rect 22310 27880 22370 27890
rect 18940 27810 19200 27820
rect 19320 27820 19380 27830
rect 18850 27430 18910 27440
rect 18850 27360 18910 27370
rect 18940 27360 18970 27810
rect 19060 27760 19320 27780
rect 22130 27820 22190 27830
rect 19060 27750 19380 27760
rect 21950 27760 22010 27770
rect 19060 27360 19090 27750
rect 21770 27700 21830 27710
rect 22370 27820 22570 27840
rect 22310 27810 22570 27820
rect 22190 27760 22450 27780
rect 22130 27750 22450 27760
rect 22010 27700 22330 27720
rect 21950 27690 22330 27700
rect 21830 27640 22210 27660
rect 21770 27630 22210 27640
rect 22180 27360 22210 27630
rect 22300 27360 22330 27690
rect 22420 27360 22450 27750
rect 22540 27360 22570 27810
rect 23670 27430 23750 27440
rect 22600 27370 22610 27430
rect 22670 27370 22680 27430
rect 22600 27360 22680 27370
rect 23670 27370 23680 27430
rect 23740 27370 23750 27430
rect 23670 27360 23750 27370
rect 23780 27360 23810 28210
rect 24130 27880 24190 27890
rect 23930 27820 24130 27840
rect 27300 27880 27360 27890
rect 23930 27810 24190 27820
rect 24310 27820 24370 27830
rect 23840 27430 23900 27440
rect 23840 27360 23900 27370
rect 23930 27360 23960 27810
rect 24050 27760 24310 27780
rect 27120 27820 27180 27830
rect 24050 27750 24370 27760
rect 24490 27760 24550 27770
rect 24050 27360 24080 27750
rect 24170 27700 24490 27720
rect 26940 27760 27000 27770
rect 24170 27690 24550 27700
rect 24670 27700 24730 27710
rect 24170 27360 24200 27690
rect 24290 27640 24670 27660
rect 24290 27630 24730 27640
rect 26760 27700 26820 27710
rect 27360 27820 27560 27840
rect 27300 27810 27560 27820
rect 27180 27760 27440 27780
rect 27120 27750 27440 27760
rect 27000 27700 27320 27720
rect 26940 27690 27320 27700
rect 26820 27640 27200 27660
rect 26760 27630 27200 27640
rect 24290 27360 24320 27630
rect 27170 27360 27200 27630
rect 27290 27360 27320 27690
rect 27410 27360 27440 27750
rect 27530 27360 27560 27810
rect 28660 27430 28740 27440
rect 27590 27370 27600 27430
rect 27660 27370 27670 27430
rect 27590 27360 27670 27370
rect 28660 27370 28670 27430
rect 28730 27370 28740 27430
rect 28660 27360 28740 27370
rect 28770 27360 28800 28210
rect 29120 27880 29180 27890
rect 28920 27820 29120 27840
rect 32290 27880 32350 27890
rect 28920 27810 29180 27820
rect 29300 27820 29360 27830
rect 28830 27430 28890 27440
rect 28830 27360 28890 27370
rect 28920 27360 28950 27810
rect 29040 27760 29300 27780
rect 32110 27820 32170 27830
rect 29040 27750 29360 27760
rect 29480 27760 29540 27770
rect 29040 27360 29070 27750
rect 29160 27700 29480 27720
rect 31930 27760 31990 27770
rect 29160 27690 29540 27700
rect 29660 27700 29720 27710
rect 29160 27360 29190 27690
rect 29280 27640 29660 27660
rect 31750 27700 31810 27710
rect 29280 27630 29720 27640
rect 31570 27640 31630 27650
rect 29280 27360 29310 27630
rect 31390 27580 31450 27590
rect 32350 27820 32550 27840
rect 32290 27810 32550 27820
rect 32170 27760 32430 27780
rect 32110 27750 32430 27760
rect 31990 27700 32310 27720
rect 31930 27690 32310 27700
rect 31810 27640 32190 27660
rect 31750 27630 32190 27640
rect 31630 27580 32070 27600
rect 31570 27570 32070 27580
rect 31450 27520 31950 27540
rect 31390 27510 31950 27520
rect 31920 27360 31950 27510
rect 32040 27360 32070 27570
rect 32160 27360 32190 27630
rect 32280 27360 32310 27690
rect 32400 27360 32430 27750
rect 32520 27360 32550 27810
rect 33650 27430 33730 27440
rect 32580 27370 32590 27430
rect 32650 27370 32660 27430
rect 32580 27360 32660 27370
rect 33650 27370 33660 27430
rect 33720 27370 33730 27430
rect 33650 27360 33730 27370
rect 33760 27360 33790 28210
rect 34110 27880 34170 27890
rect 33910 27820 34110 27840
rect 37280 27880 37340 27890
rect 33910 27810 34170 27820
rect 34290 27820 34350 27830
rect 33820 27430 33880 27440
rect 33820 27360 33880 27370
rect 33910 27360 33940 27810
rect 34030 27760 34290 27780
rect 37100 27820 37160 27830
rect 34030 27750 34350 27760
rect 34470 27760 34530 27770
rect 34030 27360 34060 27750
rect 34150 27700 34470 27720
rect 36920 27760 36980 27770
rect 34150 27690 34530 27700
rect 34650 27700 34710 27710
rect 34150 27360 34180 27690
rect 34270 27640 34650 27660
rect 36740 27700 36800 27710
rect 34270 27630 34710 27640
rect 34830 27640 34890 27650
rect 34270 27360 34300 27630
rect 34390 27580 34830 27600
rect 36560 27640 36620 27650
rect 34390 27570 34890 27580
rect 35010 27580 35070 27590
rect 34390 27360 34420 27570
rect 34510 27520 35010 27540
rect 36380 27580 36440 27590
rect 34510 27510 35070 27520
rect 36200 27520 36260 27530
rect 34510 27360 34540 27510
rect 37340 27820 37540 27840
rect 37280 27810 37540 27820
rect 37160 27760 37420 27780
rect 37100 27750 37420 27760
rect 36980 27700 37300 27720
rect 36920 27690 37300 27700
rect 36800 27640 37180 27660
rect 36740 27630 37180 27640
rect 36620 27580 37060 27600
rect 36560 27570 37060 27580
rect 36440 27520 36940 27540
rect 36380 27510 36940 27520
rect 36260 27460 36820 27480
rect 36200 27450 36820 27460
rect 36790 27360 36820 27450
rect 36910 27360 36940 27510
rect 37030 27360 37060 27570
rect 37150 27360 37180 27630
rect 37270 27360 37300 27690
rect 37390 27360 37420 27750
rect 37510 27360 37540 27810
rect 38640 27430 38720 27440
rect 37570 27370 37580 27430
rect 37640 27370 37650 27430
rect 37570 27360 37650 27370
rect 38640 27370 38650 27430
rect 38710 27370 38720 27430
rect 38640 27360 38720 27370
rect 38750 27360 38780 28210
rect 39100 27880 39160 27890
rect 38900 27820 39100 27840
rect 42270 27880 42330 27890
rect 38900 27810 39160 27820
rect 39280 27820 39340 27830
rect 38810 27430 38870 27440
rect 38810 27360 38870 27370
rect 38900 27360 38930 27810
rect 39020 27760 39280 27780
rect 42090 27820 42150 27830
rect 39020 27750 39340 27760
rect 39460 27760 39520 27770
rect 39020 27360 39050 27750
rect 39140 27700 39460 27720
rect 41910 27760 41970 27770
rect 39140 27690 39520 27700
rect 39640 27700 39700 27710
rect 39140 27360 39170 27690
rect 39260 27640 39640 27660
rect 41730 27700 41790 27710
rect 39260 27630 39700 27640
rect 39820 27640 39880 27650
rect 39260 27360 39290 27630
rect 39380 27580 39820 27600
rect 41550 27640 41610 27650
rect 39380 27570 39880 27580
rect 40000 27580 40060 27590
rect 39380 27360 39410 27570
rect 39500 27520 40000 27540
rect 41370 27580 41430 27590
rect 39500 27510 40060 27520
rect 40180 27520 40240 27530
rect 39500 27360 39530 27510
rect 39620 27460 40180 27480
rect 39620 27450 40240 27460
rect 41190 27520 41250 27530
rect 42330 27820 42530 27840
rect 42270 27810 42530 27820
rect 42150 27760 42410 27780
rect 42090 27750 42410 27760
rect 41970 27700 42290 27720
rect 41910 27690 42290 27700
rect 41790 27640 42170 27660
rect 41730 27630 42170 27640
rect 41610 27580 42050 27600
rect 41550 27570 42050 27580
rect 41430 27520 41930 27540
rect 41370 27510 41930 27520
rect 41250 27460 41810 27480
rect 41190 27450 41810 27460
rect 39620 27360 39650 27450
rect 41780 27360 41810 27450
rect 41900 27360 41930 27510
rect 42020 27360 42050 27570
rect 42140 27360 42170 27630
rect 42260 27360 42290 27690
rect 42380 27360 42410 27750
rect 42500 27360 42530 27810
rect 43630 27430 43710 27440
rect 42560 27370 42570 27430
rect 42630 27370 42640 27430
rect 42560 27360 42640 27370
rect 43630 27370 43640 27430
rect 43700 27370 43710 27430
rect 43630 27360 43710 27370
rect 43740 27360 43770 28210
rect 44090 27880 44150 27890
rect 43890 27820 44090 27840
rect 47260 27880 47320 27890
rect 43890 27810 44150 27820
rect 44270 27820 44330 27830
rect 43800 27430 43860 27440
rect 43800 27360 43860 27370
rect 43890 27360 43920 27810
rect 44010 27760 44270 27780
rect 47080 27820 47140 27830
rect 44010 27750 44330 27760
rect 44450 27760 44510 27770
rect 44010 27360 44040 27750
rect 44130 27700 44450 27720
rect 46900 27760 46960 27770
rect 44130 27690 44510 27700
rect 44630 27700 44690 27710
rect 44130 27360 44160 27690
rect 44250 27640 44630 27660
rect 46720 27700 46780 27710
rect 44250 27630 44690 27640
rect 44810 27640 44870 27650
rect 44250 27360 44280 27630
rect 44370 27580 44810 27600
rect 46540 27640 46600 27650
rect 44370 27570 44870 27580
rect 44990 27580 45050 27590
rect 44370 27330 44400 27570
rect 44490 27520 44990 27540
rect 46360 27580 46420 27590
rect 44490 27510 45050 27520
rect 45170 27520 45230 27530
rect 44490 27360 44520 27510
rect 44610 27460 45170 27480
rect 47320 27820 47520 27840
rect 47260 27810 47520 27820
rect 47140 27760 47400 27780
rect 47080 27750 47400 27760
rect 46960 27700 47280 27720
rect 46900 27690 47280 27700
rect 46780 27640 47160 27660
rect 46720 27630 47160 27640
rect 46600 27580 47040 27600
rect 46540 27570 47040 27580
rect 46420 27520 46920 27540
rect 46360 27510 46920 27520
rect 44610 27450 45230 27460
rect 44610 27360 44640 27450
rect 46890 27360 46920 27510
rect 47010 27360 47040 27570
rect 47130 27360 47160 27630
rect 47250 27360 47280 27690
rect 47370 27360 47400 27750
rect 47490 27360 47520 27810
rect 48620 27430 48700 27440
rect 47550 27370 47560 27430
rect 47620 27370 47630 27430
rect 47550 27360 47630 27370
rect 48620 27370 48630 27430
rect 48690 27370 48700 27430
rect 48620 27360 48700 27370
rect 48730 27360 48760 28210
rect 49080 27880 49140 27890
rect 48880 27820 49080 27840
rect 52250 27880 52310 27890
rect 48880 27810 49140 27820
rect 49260 27820 49320 27830
rect 48790 27430 48850 27440
rect 48790 27360 48850 27370
rect 48880 27360 48910 27810
rect 49000 27760 49260 27780
rect 52070 27820 52130 27830
rect 49000 27750 49320 27760
rect 49440 27760 49500 27770
rect 49000 27360 49030 27750
rect 49120 27700 49440 27720
rect 51890 27760 51950 27770
rect 49120 27690 49500 27700
rect 49620 27700 49680 27710
rect 49120 27360 49150 27690
rect 49240 27640 49620 27660
rect 51710 27700 51770 27710
rect 49240 27630 49680 27640
rect 49800 27640 49860 27650
rect 49240 27360 49270 27630
rect 49360 27580 49800 27600
rect 52310 27820 52510 27840
rect 52250 27810 52510 27820
rect 52130 27760 52390 27780
rect 52070 27750 52390 27760
rect 51950 27700 52270 27720
rect 51890 27690 52270 27700
rect 51770 27640 52150 27660
rect 51710 27630 52150 27640
rect 49360 27570 49860 27580
rect 49980 27580 50040 27590
rect 49360 27360 49390 27570
rect 49480 27520 49980 27540
rect 49480 27510 50040 27520
rect 49480 27360 49510 27510
rect 52120 27360 52150 27630
rect 52240 27360 52270 27690
rect 52360 27360 52390 27750
rect 52480 27360 52510 27810
rect 53610 27430 53690 27440
rect 52540 27370 52550 27430
rect 52610 27370 52620 27430
rect 52540 27360 52620 27370
rect 53610 27370 53620 27430
rect 53680 27370 53690 27430
rect 53610 27360 53690 27370
rect 53720 27360 53750 28210
rect 54070 27880 54130 27890
rect 53870 27820 54070 27840
rect 57240 27880 57300 27890
rect 53870 27810 54130 27820
rect 54250 27820 54310 27830
rect 53780 27430 53840 27440
rect 53780 27360 53840 27370
rect 53870 27360 53900 27810
rect 53990 27760 54250 27780
rect 57060 27820 57120 27830
rect 53990 27750 54310 27760
rect 54430 27760 54490 27770
rect 53990 27360 54020 27750
rect 54110 27700 54430 27720
rect 56880 27760 56940 27770
rect 54110 27690 54490 27700
rect 54610 27700 54670 27710
rect 54110 27360 54140 27690
rect 54230 27640 54610 27660
rect 54230 27630 54670 27640
rect 56700 27700 56760 27710
rect 57300 27820 57500 27840
rect 57240 27810 57500 27820
rect 57120 27760 57380 27780
rect 57060 27750 57380 27760
rect 56940 27700 57260 27720
rect 56880 27690 57260 27700
rect 56760 27640 57140 27660
rect 56700 27630 57140 27640
rect 54230 27360 54260 27630
rect 57110 27360 57140 27630
rect 57230 27360 57260 27690
rect 57350 27360 57380 27750
rect 57470 27360 57500 27810
rect 58600 27430 58680 27440
rect 57530 27370 57540 27430
rect 57600 27370 57610 27430
rect 57530 27360 57610 27370
rect 58600 27370 58610 27430
rect 58670 27370 58680 27430
rect 58600 27360 58680 27370
rect 58710 27360 58740 28210
rect 59060 27880 59120 27890
rect 58860 27820 59060 27840
rect 62230 27880 62290 27890
rect 58860 27810 59120 27820
rect 59240 27820 59300 27830
rect 58770 27430 58830 27440
rect 58770 27360 58830 27370
rect 58860 27360 58890 27810
rect 58980 27760 59240 27780
rect 62050 27820 62110 27830
rect 58980 27750 59300 27760
rect 59420 27760 59480 27770
rect 58980 27360 59010 27750
rect 59100 27700 59420 27720
rect 62290 27820 62490 27840
rect 62230 27810 62490 27820
rect 62110 27760 62370 27780
rect 62050 27750 62370 27760
rect 59100 27690 59480 27700
rect 59600 27700 59660 27710
rect 59100 27360 59130 27690
rect 59220 27640 59600 27660
rect 59220 27630 59660 27640
rect 59220 27360 59250 27630
rect 62340 27360 62370 27750
rect 62460 27360 62490 27810
rect 63590 27430 63670 27440
rect 62520 27370 62530 27430
rect 62590 27370 62600 27430
rect 62520 27360 62600 27370
rect 63590 27370 63600 27430
rect 63660 27370 63670 27430
rect 63590 27360 63670 27370
rect 63700 27360 63730 28210
rect 64050 27880 64110 27890
rect 63850 27820 64050 27840
rect 67220 27880 67280 27890
rect 63850 27810 64110 27820
rect 64230 27820 64290 27830
rect 63760 27430 63820 27440
rect 63760 27360 63820 27370
rect 63850 27360 63880 27810
rect 63970 27760 64230 27780
rect 63970 27750 64290 27760
rect 67040 27820 67100 27830
rect 67280 27820 67480 27840
rect 67220 27810 67480 27820
rect 67100 27760 67360 27780
rect 67040 27750 67360 27760
rect 63970 27360 64000 27750
rect 67330 27360 67360 27750
rect 67450 27360 67480 27810
rect 68580 27430 68660 27440
rect 67510 27370 67520 27430
rect 67580 27370 67590 27430
rect 67510 27360 67590 27370
rect 68580 27370 68590 27430
rect 68650 27370 68660 27430
rect 68580 27360 68660 27370
rect 68690 27360 68720 28210
rect 69040 27880 69100 27890
rect 68840 27820 69040 27840
rect 72210 27880 72270 27890
rect 68840 27810 69100 27820
rect 69220 27820 69280 27830
rect 68750 27430 68810 27440
rect 68750 27360 68810 27370
rect 68840 27360 68870 27810
rect 68960 27760 69220 27780
rect 72270 27820 72470 27840
rect 72210 27810 72470 27820
rect 68960 27750 69280 27760
rect 68960 27360 68990 27750
rect 72440 27360 72470 27810
rect 73570 27430 73650 27440
rect 72500 27370 72510 27430
rect 72570 27370 72580 27430
rect 72500 27360 72580 27370
rect 73570 27370 73580 27430
rect 73640 27370 73650 27430
rect 73570 27360 73650 27370
rect 73680 27360 73710 28210
rect 74030 27880 74090 27890
rect 73830 27820 74030 27840
rect 73830 27810 74090 27820
rect 77200 27880 77260 27890
rect 77260 27820 77460 27840
rect 77200 27810 77460 27820
rect 73740 27430 73800 27440
rect 73740 27360 73800 27370
rect 73830 27360 73860 27810
rect 77430 27360 77460 27810
rect 78560 27430 78640 27440
rect 77490 27370 77500 27430
rect 77560 27370 77570 27430
rect 77490 27360 77570 27370
rect 78560 27370 78570 27430
rect 78630 27370 78640 27430
rect 78560 27360 78640 27370
rect 78670 27360 78700 28210
rect 79020 27880 79080 27890
rect 78820 27820 79020 27840
rect 78820 27810 79080 27820
rect 78730 27430 78790 27440
rect 78730 27360 78790 27370
rect 78820 27360 78850 27810
rect 82714 16840 104970 52994
<< via1 >>
rect 2650 66320 2710 66380
rect 2650 64610 2710 64670
rect 2650 62900 2710 62960
rect 2650 61190 2710 61250
rect 2650 59480 2710 59540
rect 2650 57770 2710 57830
rect 2650 56060 2710 56120
rect 2650 54350 2710 54410
rect 2650 52640 2710 52700
rect 2650 50930 2710 50990
rect 2650 49220 2710 49280
rect 2650 47510 2710 47570
rect 2650 45800 2710 45860
rect 2650 44090 2710 44150
rect 2650 42380 2710 42440
rect 2650 40670 2710 40730
rect 2860 66358 2920 66370
rect 3280 66380 3340 66440
rect 2860 66324 2888 66358
rect 2888 66324 2920 66358
rect 2860 66310 2920 66324
rect 3700 66358 3760 66370
rect 3700 66324 3705 66358
rect 3705 66324 3739 66358
rect 3739 66324 3760 66358
rect 3700 66310 3760 66324
rect 3280 66210 3340 66270
rect 3280 66100 3340 66160
rect 2860 66048 2920 66060
rect 2860 66014 2888 66048
rect 2888 66014 2920 66048
rect 2860 66000 2920 66014
rect 3280 65930 3340 65990
rect 3700 66048 3760 66060
rect 3700 66014 3705 66048
rect 3705 66014 3739 66048
rect 3739 66014 3760 66048
rect 3700 66000 3760 66014
rect 2860 64648 2920 64660
rect 3280 64670 3340 64730
rect 2860 64614 2888 64648
rect 2888 64614 2920 64648
rect 2860 64600 2920 64614
rect 3700 64648 3760 64660
rect 3700 64614 3705 64648
rect 3705 64614 3739 64648
rect 3739 64614 3760 64648
rect 3700 64600 3760 64614
rect 3280 64500 3340 64560
rect 3280 64390 3340 64450
rect 2860 64338 2920 64350
rect 2860 64304 2888 64338
rect 2888 64304 2920 64338
rect 2860 64290 2920 64304
rect 3280 64220 3340 64280
rect 3700 64338 3760 64350
rect 3700 64304 3705 64338
rect 3705 64304 3739 64338
rect 3739 64304 3760 64338
rect 3700 64290 3760 64304
rect 2860 62938 2920 62950
rect 3280 62960 3340 63020
rect 2860 62904 2888 62938
rect 2888 62904 2920 62938
rect 2860 62890 2920 62904
rect 3700 62938 3760 62950
rect 3700 62904 3705 62938
rect 3705 62904 3739 62938
rect 3739 62904 3760 62938
rect 3700 62890 3760 62904
rect 3280 62790 3340 62850
rect 3280 62680 3340 62740
rect 2860 62628 2920 62640
rect 2860 62594 2888 62628
rect 2888 62594 2920 62628
rect 2860 62580 2920 62594
rect 3280 62510 3340 62570
rect 3700 62628 3760 62640
rect 3700 62594 3705 62628
rect 3705 62594 3739 62628
rect 3739 62594 3760 62628
rect 3700 62580 3760 62594
rect 2860 61228 2920 61240
rect 3280 61250 3340 61310
rect 2860 61194 2888 61228
rect 2888 61194 2920 61228
rect 2860 61180 2920 61194
rect 3700 61228 3760 61240
rect 3700 61194 3705 61228
rect 3705 61194 3739 61228
rect 3739 61194 3760 61228
rect 3700 61180 3760 61194
rect 3280 61080 3340 61140
rect 3280 60970 3340 61030
rect 2860 60918 2920 60930
rect 2860 60884 2888 60918
rect 2888 60884 2920 60918
rect 2860 60870 2920 60884
rect 3280 60800 3340 60860
rect 3700 60918 3760 60930
rect 3700 60884 3705 60918
rect 3705 60884 3739 60918
rect 3739 60884 3760 60918
rect 3700 60870 3760 60884
rect 2860 59518 2920 59530
rect 3280 59540 3340 59600
rect 2860 59484 2888 59518
rect 2888 59484 2920 59518
rect 2860 59470 2920 59484
rect 3700 59518 3760 59530
rect 3700 59484 3705 59518
rect 3705 59484 3739 59518
rect 3739 59484 3760 59518
rect 3700 59470 3760 59484
rect 3280 59370 3340 59430
rect 3280 59260 3340 59320
rect 2860 59208 2920 59220
rect 2860 59174 2888 59208
rect 2888 59174 2920 59208
rect 2860 59160 2920 59174
rect 3280 59090 3340 59150
rect 3700 59208 3760 59220
rect 3700 59174 3705 59208
rect 3705 59174 3739 59208
rect 3739 59174 3760 59208
rect 3700 59160 3760 59174
rect 2860 57808 2920 57820
rect 3280 57830 3340 57890
rect 2860 57774 2888 57808
rect 2888 57774 2920 57808
rect 2860 57760 2920 57774
rect 3700 57808 3760 57820
rect 3700 57774 3705 57808
rect 3705 57774 3739 57808
rect 3739 57774 3760 57808
rect 3700 57760 3760 57774
rect 3280 57660 3340 57720
rect 3280 57550 3340 57610
rect 2860 57498 2920 57510
rect 2860 57464 2888 57498
rect 2888 57464 2920 57498
rect 2860 57450 2920 57464
rect 3280 57380 3340 57440
rect 3700 57498 3760 57510
rect 3700 57464 3705 57498
rect 3705 57464 3739 57498
rect 3739 57464 3760 57498
rect 3700 57450 3760 57464
rect 2860 56098 2920 56110
rect 3280 56120 3340 56180
rect 2860 56064 2888 56098
rect 2888 56064 2920 56098
rect 2860 56050 2920 56064
rect 3700 56098 3760 56110
rect 3700 56064 3705 56098
rect 3705 56064 3739 56098
rect 3739 56064 3760 56098
rect 3700 56050 3760 56064
rect 3280 55950 3340 56010
rect 3280 55840 3340 55900
rect 2860 55788 2920 55800
rect 2860 55754 2888 55788
rect 2888 55754 2920 55788
rect 2860 55740 2920 55754
rect 3280 55670 3340 55730
rect 3700 55788 3760 55800
rect 3700 55754 3705 55788
rect 3705 55754 3739 55788
rect 3739 55754 3760 55788
rect 3700 55740 3760 55754
rect 2860 54388 2920 54400
rect 3280 54410 3340 54470
rect 2860 54354 2888 54388
rect 2888 54354 2920 54388
rect 2860 54340 2920 54354
rect 3700 54388 3760 54400
rect 3700 54354 3705 54388
rect 3705 54354 3739 54388
rect 3739 54354 3760 54388
rect 3700 54340 3760 54354
rect 3280 54240 3340 54300
rect 3280 54130 3340 54190
rect 2860 54078 2920 54090
rect 2860 54044 2888 54078
rect 2888 54044 2920 54078
rect 2860 54030 2920 54044
rect 3280 53960 3340 54020
rect 3700 54078 3760 54090
rect 3700 54044 3705 54078
rect 3705 54044 3739 54078
rect 3739 54044 3760 54078
rect 3700 54030 3760 54044
rect 2860 52678 2920 52690
rect 3280 52700 3340 52760
rect 2860 52644 2888 52678
rect 2888 52644 2920 52678
rect 2860 52630 2920 52644
rect 3700 52678 3760 52690
rect 3700 52644 3705 52678
rect 3705 52644 3739 52678
rect 3739 52644 3760 52678
rect 3700 52630 3760 52644
rect 3280 52530 3340 52590
rect 3280 52420 3340 52480
rect 2860 52368 2920 52380
rect 2860 52334 2888 52368
rect 2888 52334 2920 52368
rect 2860 52320 2920 52334
rect 3280 52250 3340 52310
rect 3700 52368 3760 52380
rect 3700 52334 3705 52368
rect 3705 52334 3739 52368
rect 3739 52334 3760 52368
rect 3700 52320 3760 52334
rect 2860 50968 2920 50980
rect 3280 50990 3340 51050
rect 2860 50934 2888 50968
rect 2888 50934 2920 50968
rect 2860 50920 2920 50934
rect 3700 50968 3760 50980
rect 3700 50934 3705 50968
rect 3705 50934 3739 50968
rect 3739 50934 3760 50968
rect 3700 50920 3760 50934
rect 3280 50820 3340 50880
rect 3280 50710 3340 50770
rect 2860 50658 2920 50670
rect 2860 50624 2888 50658
rect 2888 50624 2920 50658
rect 2860 50610 2920 50624
rect 3280 50540 3340 50600
rect 3700 50658 3760 50670
rect 3700 50624 3705 50658
rect 3705 50624 3739 50658
rect 3739 50624 3760 50658
rect 3700 50610 3760 50624
rect 2860 49258 2920 49270
rect 3280 49280 3340 49340
rect 2860 49224 2888 49258
rect 2888 49224 2920 49258
rect 2860 49210 2920 49224
rect 3700 49258 3760 49270
rect 3700 49224 3705 49258
rect 3705 49224 3739 49258
rect 3739 49224 3760 49258
rect 3700 49210 3760 49224
rect 3280 49110 3340 49170
rect 3280 49000 3340 49060
rect 2860 48948 2920 48960
rect 2860 48914 2888 48948
rect 2888 48914 2920 48948
rect 2860 48900 2920 48914
rect 3280 48830 3340 48890
rect 3700 48948 3760 48960
rect 3700 48914 3705 48948
rect 3705 48914 3739 48948
rect 3739 48914 3760 48948
rect 3700 48900 3760 48914
rect 2860 47548 2920 47560
rect 3280 47570 3340 47630
rect 2860 47514 2888 47548
rect 2888 47514 2920 47548
rect 2860 47500 2920 47514
rect 3700 47548 3760 47560
rect 3700 47514 3705 47548
rect 3705 47514 3739 47548
rect 3739 47514 3760 47548
rect 3700 47500 3760 47514
rect 3280 47400 3340 47460
rect 3280 47290 3340 47350
rect 2860 47238 2920 47250
rect 2860 47204 2888 47238
rect 2888 47204 2920 47238
rect 2860 47190 2920 47204
rect 3280 47120 3340 47180
rect 3700 47238 3760 47250
rect 3700 47204 3705 47238
rect 3705 47204 3739 47238
rect 3739 47204 3760 47238
rect 3700 47190 3760 47204
rect 2860 45838 2920 45850
rect 3280 45860 3340 45920
rect 2860 45804 2888 45838
rect 2888 45804 2920 45838
rect 2860 45790 2920 45804
rect 3700 45838 3760 45850
rect 3700 45804 3705 45838
rect 3705 45804 3739 45838
rect 3739 45804 3760 45838
rect 3700 45790 3760 45804
rect 3280 45690 3340 45750
rect 3280 45580 3340 45640
rect 2860 45528 2920 45540
rect 2860 45494 2888 45528
rect 2888 45494 2920 45528
rect 2860 45480 2920 45494
rect 3280 45410 3340 45470
rect 3700 45528 3760 45540
rect 3700 45494 3705 45528
rect 3705 45494 3739 45528
rect 3739 45494 3760 45528
rect 3700 45480 3760 45494
rect 2860 44128 2920 44140
rect 3280 44150 3340 44210
rect 2860 44094 2888 44128
rect 2888 44094 2920 44128
rect 2860 44080 2920 44094
rect 3700 44128 3760 44140
rect 3700 44094 3705 44128
rect 3705 44094 3739 44128
rect 3739 44094 3760 44128
rect 3700 44080 3760 44094
rect 3280 43980 3340 44040
rect 3280 43870 3340 43930
rect 2860 43818 2920 43830
rect 2860 43784 2888 43818
rect 2888 43784 2920 43818
rect 2860 43770 2920 43784
rect 3280 43700 3340 43760
rect 3700 43818 3760 43830
rect 3700 43784 3705 43818
rect 3705 43784 3739 43818
rect 3739 43784 3760 43818
rect 3700 43770 3760 43784
rect 2860 42418 2920 42430
rect 3280 42440 3340 42500
rect 2860 42384 2888 42418
rect 2888 42384 2920 42418
rect 2860 42370 2920 42384
rect 3700 42418 3760 42430
rect 3700 42384 3705 42418
rect 3705 42384 3739 42418
rect 3739 42384 3760 42418
rect 3700 42370 3760 42384
rect 3280 42270 3340 42330
rect 3280 42160 3340 42220
rect 2860 42108 2920 42120
rect 2860 42074 2888 42108
rect 2888 42074 2920 42108
rect 2860 42060 2920 42074
rect 3280 41990 3340 42050
rect 3700 42108 3760 42120
rect 3700 42074 3705 42108
rect 3705 42074 3739 42108
rect 3739 42074 3760 42108
rect 3700 42060 3760 42074
rect 2860 40708 2920 40720
rect 3280 40730 3340 40790
rect 2860 40674 2888 40708
rect 2888 40674 2920 40708
rect 2860 40660 2920 40674
rect 3700 40708 3760 40720
rect 3700 40674 3705 40708
rect 3705 40674 3739 40708
rect 3739 40674 3760 40708
rect 3700 40660 3760 40674
rect 3280 40560 3340 40620
rect 3280 40450 3340 40510
rect 2860 40398 2920 40410
rect 2860 40364 2888 40398
rect 2888 40364 2920 40398
rect 2860 40350 2920 40364
rect 3280 40280 3340 40340
rect 3700 40398 3760 40410
rect 3700 40364 3705 40398
rect 3705 40364 3739 40398
rect 3739 40364 3760 40398
rect 3700 40350 3760 40364
rect 2750 39620 2810 39680
rect 3820 39620 3880 39680
rect 3920 66410 3980 66470
rect 3980 65880 4040 65940
rect 3920 64700 3980 64760
rect 3980 64170 4040 64230
rect 3920 62990 3980 63050
rect 3980 62460 4040 62520
rect 3920 61280 3980 61340
rect 3980 60750 4040 60810
rect 3920 59570 3980 59630
rect 3980 59040 4040 59100
rect 3920 57860 3980 57920
rect 3980 57330 4040 57390
rect 3920 56150 3980 56210
rect 3980 55620 4040 55680
rect 3920 54440 3980 54500
rect 3980 53910 4040 53970
rect 3920 52730 3980 52790
rect 3980 52200 4040 52260
rect 3920 51020 3980 51080
rect 3980 50490 4040 50550
rect 3920 49310 3980 49370
rect 3980 48780 4040 48840
rect 3920 47600 3980 47660
rect 3980 47070 4040 47130
rect 3920 45890 3980 45950
rect 3980 45360 4040 45420
rect 3920 44180 3980 44240
rect 3980 43650 4040 43710
rect 3920 42470 3980 42530
rect 3980 41940 4040 42000
rect 3920 40760 3980 40820
rect 2450 39170 2510 39230
rect 3980 40230 4040 40290
rect 3980 39620 4040 39680
rect 4070 66320 4130 66380
rect 4070 64610 4130 64670
rect 4070 62900 4130 62960
rect 4070 61190 4130 61250
rect 4070 59480 4130 59540
rect 4070 57770 4130 57830
rect 4070 56060 4130 56120
rect 4070 54350 4130 54410
rect 4070 52640 4130 52700
rect 4070 50930 4130 50990
rect 4070 49220 4130 49280
rect 4070 47510 4130 47570
rect 4070 45800 4130 45860
rect 4070 44090 4130 44150
rect 4070 42380 4130 42440
rect 4070 40670 4130 40730
rect 7640 66320 7700 66380
rect 7640 64610 7700 64670
rect 7640 62900 7700 62960
rect 7640 61190 7700 61250
rect 7640 59480 7700 59540
rect 7640 57770 7700 57830
rect 7640 56060 7700 56120
rect 7640 54350 7700 54410
rect 7640 52640 7700 52700
rect 7640 50930 7700 50990
rect 7640 49220 7700 49280
rect 7640 47510 7700 47570
rect 7640 45800 7700 45860
rect 7640 44090 7700 44150
rect 7640 42380 7700 42440
rect 7640 40670 7700 40730
rect 7850 66358 7910 66370
rect 8270 66380 8330 66440
rect 7850 66324 7878 66358
rect 7878 66324 7910 66358
rect 7850 66310 7910 66324
rect 8690 66358 8750 66370
rect 8690 66324 8695 66358
rect 8695 66324 8729 66358
rect 8729 66324 8750 66358
rect 8690 66310 8750 66324
rect 8270 66210 8330 66270
rect 8270 66100 8330 66160
rect 7850 66048 7910 66060
rect 7850 66014 7878 66048
rect 7878 66014 7910 66048
rect 7850 66000 7910 66014
rect 8270 65930 8330 65990
rect 8690 66048 8750 66060
rect 8690 66014 8695 66048
rect 8695 66014 8729 66048
rect 8729 66014 8750 66048
rect 8690 66000 8750 66014
rect 7850 64648 7910 64660
rect 8270 64670 8330 64730
rect 7850 64614 7878 64648
rect 7878 64614 7910 64648
rect 7850 64600 7910 64614
rect 8690 64648 8750 64660
rect 8690 64614 8695 64648
rect 8695 64614 8729 64648
rect 8729 64614 8750 64648
rect 8690 64600 8750 64614
rect 8270 64500 8330 64560
rect 8270 64390 8330 64450
rect 7850 64338 7910 64350
rect 7850 64304 7878 64338
rect 7878 64304 7910 64338
rect 7850 64290 7910 64304
rect 8270 64220 8330 64280
rect 8690 64338 8750 64350
rect 8690 64304 8695 64338
rect 8695 64304 8729 64338
rect 8729 64304 8750 64338
rect 8690 64290 8750 64304
rect 7850 62938 7910 62950
rect 8270 62960 8330 63020
rect 7850 62904 7878 62938
rect 7878 62904 7910 62938
rect 7850 62890 7910 62904
rect 8690 62938 8750 62950
rect 8690 62904 8695 62938
rect 8695 62904 8729 62938
rect 8729 62904 8750 62938
rect 8690 62890 8750 62904
rect 8270 62790 8330 62850
rect 8270 62680 8330 62740
rect 7850 62628 7910 62640
rect 7850 62594 7878 62628
rect 7878 62594 7910 62628
rect 7850 62580 7910 62594
rect 8270 62510 8330 62570
rect 8690 62628 8750 62640
rect 8690 62594 8695 62628
rect 8695 62594 8729 62628
rect 8729 62594 8750 62628
rect 8690 62580 8750 62594
rect 7850 61228 7910 61240
rect 8270 61250 8330 61310
rect 7850 61194 7878 61228
rect 7878 61194 7910 61228
rect 7850 61180 7910 61194
rect 8690 61228 8750 61240
rect 8690 61194 8695 61228
rect 8695 61194 8729 61228
rect 8729 61194 8750 61228
rect 8690 61180 8750 61194
rect 8270 61080 8330 61140
rect 8270 60970 8330 61030
rect 7850 60918 7910 60930
rect 7850 60884 7878 60918
rect 7878 60884 7910 60918
rect 7850 60870 7910 60884
rect 8270 60800 8330 60860
rect 8690 60918 8750 60930
rect 8690 60884 8695 60918
rect 8695 60884 8729 60918
rect 8729 60884 8750 60918
rect 8690 60870 8750 60884
rect 7850 59518 7910 59530
rect 8270 59540 8330 59600
rect 7850 59484 7878 59518
rect 7878 59484 7910 59518
rect 7850 59470 7910 59484
rect 8690 59518 8750 59530
rect 8690 59484 8695 59518
rect 8695 59484 8729 59518
rect 8729 59484 8750 59518
rect 8690 59470 8750 59484
rect 8270 59370 8330 59430
rect 8270 59260 8330 59320
rect 7850 59208 7910 59220
rect 7850 59174 7878 59208
rect 7878 59174 7910 59208
rect 7850 59160 7910 59174
rect 8270 59090 8330 59150
rect 8690 59208 8750 59220
rect 8690 59174 8695 59208
rect 8695 59174 8729 59208
rect 8729 59174 8750 59208
rect 8690 59160 8750 59174
rect 7850 57808 7910 57820
rect 8270 57830 8330 57890
rect 7850 57774 7878 57808
rect 7878 57774 7910 57808
rect 7850 57760 7910 57774
rect 8690 57808 8750 57820
rect 8690 57774 8695 57808
rect 8695 57774 8729 57808
rect 8729 57774 8750 57808
rect 8690 57760 8750 57774
rect 8270 57660 8330 57720
rect 8270 57550 8330 57610
rect 7850 57498 7910 57510
rect 7850 57464 7878 57498
rect 7878 57464 7910 57498
rect 7850 57450 7910 57464
rect 8270 57380 8330 57440
rect 8690 57498 8750 57510
rect 8690 57464 8695 57498
rect 8695 57464 8729 57498
rect 8729 57464 8750 57498
rect 8690 57450 8750 57464
rect 7850 56098 7910 56110
rect 8270 56120 8330 56180
rect 7850 56064 7878 56098
rect 7878 56064 7910 56098
rect 7850 56050 7910 56064
rect 8690 56098 8750 56110
rect 8690 56064 8695 56098
rect 8695 56064 8729 56098
rect 8729 56064 8750 56098
rect 8690 56050 8750 56064
rect 8270 55950 8330 56010
rect 8270 55840 8330 55900
rect 7850 55788 7910 55800
rect 7850 55754 7878 55788
rect 7878 55754 7910 55788
rect 7850 55740 7910 55754
rect 8270 55670 8330 55730
rect 8690 55788 8750 55800
rect 8690 55754 8695 55788
rect 8695 55754 8729 55788
rect 8729 55754 8750 55788
rect 8690 55740 8750 55754
rect 7850 54388 7910 54400
rect 8270 54410 8330 54470
rect 7850 54354 7878 54388
rect 7878 54354 7910 54388
rect 7850 54340 7910 54354
rect 8690 54388 8750 54400
rect 8690 54354 8695 54388
rect 8695 54354 8729 54388
rect 8729 54354 8750 54388
rect 8690 54340 8750 54354
rect 8270 54240 8330 54300
rect 8270 54130 8330 54190
rect 7850 54078 7910 54090
rect 7850 54044 7878 54078
rect 7878 54044 7910 54078
rect 7850 54030 7910 54044
rect 8270 53960 8330 54020
rect 8690 54078 8750 54090
rect 8690 54044 8695 54078
rect 8695 54044 8729 54078
rect 8729 54044 8750 54078
rect 8690 54030 8750 54044
rect 7850 52678 7910 52690
rect 8270 52700 8330 52760
rect 7850 52644 7878 52678
rect 7878 52644 7910 52678
rect 7850 52630 7910 52644
rect 8690 52678 8750 52690
rect 8690 52644 8695 52678
rect 8695 52644 8729 52678
rect 8729 52644 8750 52678
rect 8690 52630 8750 52644
rect 8270 52530 8330 52590
rect 8270 52420 8330 52480
rect 7850 52368 7910 52380
rect 7850 52334 7878 52368
rect 7878 52334 7910 52368
rect 7850 52320 7910 52334
rect 8270 52250 8330 52310
rect 8690 52368 8750 52380
rect 8690 52334 8695 52368
rect 8695 52334 8729 52368
rect 8729 52334 8750 52368
rect 8690 52320 8750 52334
rect 7850 50968 7910 50980
rect 8270 50990 8330 51050
rect 7850 50934 7878 50968
rect 7878 50934 7910 50968
rect 7850 50920 7910 50934
rect 8690 50968 8750 50980
rect 8690 50934 8695 50968
rect 8695 50934 8729 50968
rect 8729 50934 8750 50968
rect 8690 50920 8750 50934
rect 8270 50820 8330 50880
rect 8270 50710 8330 50770
rect 7850 50658 7910 50670
rect 7850 50624 7878 50658
rect 7878 50624 7910 50658
rect 7850 50610 7910 50624
rect 8270 50540 8330 50600
rect 8690 50658 8750 50670
rect 8690 50624 8695 50658
rect 8695 50624 8729 50658
rect 8729 50624 8750 50658
rect 8690 50610 8750 50624
rect 7850 49258 7910 49270
rect 8270 49280 8330 49340
rect 7850 49224 7878 49258
rect 7878 49224 7910 49258
rect 7850 49210 7910 49224
rect 8690 49258 8750 49270
rect 8690 49224 8695 49258
rect 8695 49224 8729 49258
rect 8729 49224 8750 49258
rect 8690 49210 8750 49224
rect 8270 49110 8330 49170
rect 8270 49000 8330 49060
rect 7850 48948 7910 48960
rect 7850 48914 7878 48948
rect 7878 48914 7910 48948
rect 7850 48900 7910 48914
rect 8270 48830 8330 48890
rect 8690 48948 8750 48960
rect 8690 48914 8695 48948
rect 8695 48914 8729 48948
rect 8729 48914 8750 48948
rect 8690 48900 8750 48914
rect 7850 47548 7910 47560
rect 8270 47570 8330 47630
rect 7850 47514 7878 47548
rect 7878 47514 7910 47548
rect 7850 47500 7910 47514
rect 8690 47548 8750 47560
rect 8690 47514 8695 47548
rect 8695 47514 8729 47548
rect 8729 47514 8750 47548
rect 8690 47500 8750 47514
rect 8270 47400 8330 47460
rect 8270 47290 8330 47350
rect 7850 47238 7910 47250
rect 7850 47204 7878 47238
rect 7878 47204 7910 47238
rect 7850 47190 7910 47204
rect 8270 47120 8330 47180
rect 8690 47238 8750 47250
rect 8690 47204 8695 47238
rect 8695 47204 8729 47238
rect 8729 47204 8750 47238
rect 8690 47190 8750 47204
rect 7850 45838 7910 45850
rect 8270 45860 8330 45920
rect 7850 45804 7878 45838
rect 7878 45804 7910 45838
rect 7850 45790 7910 45804
rect 8690 45838 8750 45850
rect 8690 45804 8695 45838
rect 8695 45804 8729 45838
rect 8729 45804 8750 45838
rect 8690 45790 8750 45804
rect 8270 45690 8330 45750
rect 8270 45580 8330 45640
rect 7850 45528 7910 45540
rect 7850 45494 7878 45528
rect 7878 45494 7910 45528
rect 7850 45480 7910 45494
rect 8270 45410 8330 45470
rect 8690 45528 8750 45540
rect 8690 45494 8695 45528
rect 8695 45494 8729 45528
rect 8729 45494 8750 45528
rect 8690 45480 8750 45494
rect 7850 44128 7910 44140
rect 8270 44150 8330 44210
rect 7850 44094 7878 44128
rect 7878 44094 7910 44128
rect 7850 44080 7910 44094
rect 8690 44128 8750 44140
rect 8690 44094 8695 44128
rect 8695 44094 8729 44128
rect 8729 44094 8750 44128
rect 8690 44080 8750 44094
rect 8270 43980 8330 44040
rect 8270 43870 8330 43930
rect 7850 43818 7910 43830
rect 7850 43784 7878 43818
rect 7878 43784 7910 43818
rect 7850 43770 7910 43784
rect 8270 43700 8330 43760
rect 8690 43818 8750 43830
rect 8690 43784 8695 43818
rect 8695 43784 8729 43818
rect 8729 43784 8750 43818
rect 8690 43770 8750 43784
rect 7850 42418 7910 42430
rect 8270 42440 8330 42500
rect 7850 42384 7878 42418
rect 7878 42384 7910 42418
rect 7850 42370 7910 42384
rect 8690 42418 8750 42430
rect 8690 42384 8695 42418
rect 8695 42384 8729 42418
rect 8729 42384 8750 42418
rect 8690 42370 8750 42384
rect 8270 42270 8330 42330
rect 8270 42160 8330 42220
rect 7850 42108 7910 42120
rect 7850 42074 7878 42108
rect 7878 42074 7910 42108
rect 7850 42060 7910 42074
rect 8270 41990 8330 42050
rect 8690 42108 8750 42120
rect 8690 42074 8695 42108
rect 8695 42074 8729 42108
rect 8729 42074 8750 42108
rect 8690 42060 8750 42074
rect 7850 40708 7910 40720
rect 8270 40730 8330 40790
rect 7850 40674 7878 40708
rect 7878 40674 7910 40708
rect 7850 40660 7910 40674
rect 8690 40708 8750 40720
rect 8690 40674 8695 40708
rect 8695 40674 8729 40708
rect 8729 40674 8750 40708
rect 8690 40660 8750 40674
rect 8270 40560 8330 40620
rect 8270 40450 8330 40510
rect 7850 40398 7910 40410
rect 7850 40364 7878 40398
rect 7878 40364 7910 40398
rect 7850 40350 7910 40364
rect 8270 40280 8330 40340
rect 8690 40398 8750 40410
rect 8690 40364 8695 40398
rect 8695 40364 8729 40398
rect 8729 40364 8750 40398
rect 8690 40350 8750 40364
rect 7740 39620 7800 39680
rect 8810 39620 8870 39680
rect 8910 66410 8970 66470
rect 8970 65880 9030 65940
rect 8910 64700 8970 64760
rect 8970 64170 9030 64230
rect 8910 62990 8970 63050
rect 8970 62460 9030 62520
rect 8910 61280 8970 61340
rect 8970 60750 9030 60810
rect 8910 59570 8970 59630
rect 8970 59040 9030 59100
rect 8910 57860 8970 57920
rect 8970 57330 9030 57390
rect 8910 56150 8970 56210
rect 8970 55620 9030 55680
rect 8910 54440 8970 54500
rect 8970 53910 9030 53970
rect 8910 52730 8970 52790
rect 8970 52200 9030 52260
rect 8910 51020 8970 51080
rect 8970 50490 9030 50550
rect 8910 49310 8970 49370
rect 8970 48780 9030 48840
rect 8910 47600 8970 47660
rect 8970 47070 9030 47130
rect 8910 45890 8970 45950
rect 8970 45360 9030 45420
rect 8910 44180 8970 44240
rect 8970 43650 9030 43710
rect 8910 42470 8970 42530
rect 8970 41940 9030 42000
rect 8910 40760 8970 40820
rect 4270 39170 4330 39230
rect 7440 39170 7500 39230
rect 8970 40230 9030 40290
rect 8970 39620 9030 39680
rect 9060 66320 9120 66380
rect 9060 64610 9120 64670
rect 9060 62900 9120 62960
rect 9060 61190 9120 61250
rect 9060 59480 9120 59540
rect 9060 57770 9120 57830
rect 9060 56060 9120 56120
rect 9060 54350 9120 54410
rect 9060 52640 9120 52700
rect 9060 50930 9120 50990
rect 9060 49220 9120 49280
rect 9060 47510 9120 47570
rect 9060 45800 9120 45860
rect 9060 44090 9120 44150
rect 9060 42380 9120 42440
rect 9060 40670 9120 40730
rect 12630 66320 12690 66380
rect 12630 64610 12690 64670
rect 12630 62900 12690 62960
rect 12630 61190 12690 61250
rect 12510 59480 12570 59540
rect 12510 57770 12570 57830
rect 12510 56060 12570 56120
rect 12510 54350 12570 54410
rect 12510 52640 12570 52700
rect 12510 50930 12570 50990
rect 12510 49220 12570 49280
rect 12510 47510 12570 47570
rect 12630 45800 12690 45860
rect 12630 44090 12690 44150
rect 12630 42380 12690 42440
rect 12630 40670 12690 40730
rect 9260 39170 9320 39230
rect 12250 39230 12310 39290
rect 12840 66358 12900 66370
rect 13260 66380 13320 66440
rect 12840 66324 12868 66358
rect 12868 66324 12900 66358
rect 12840 66310 12900 66324
rect 13680 66358 13740 66370
rect 13680 66324 13685 66358
rect 13685 66324 13719 66358
rect 13719 66324 13740 66358
rect 13680 66310 13740 66324
rect 13260 66210 13320 66270
rect 13260 66100 13320 66160
rect 12840 66048 12900 66060
rect 12840 66014 12868 66048
rect 12868 66014 12900 66048
rect 12840 66000 12900 66014
rect 13260 65930 13320 65990
rect 13680 66048 13740 66060
rect 13680 66014 13685 66048
rect 13685 66014 13719 66048
rect 13719 66014 13740 66048
rect 13680 66000 13740 66014
rect 12840 64648 12900 64660
rect 13260 64670 13320 64730
rect 12840 64614 12868 64648
rect 12868 64614 12900 64648
rect 12840 64600 12900 64614
rect 13680 64648 13740 64660
rect 13680 64614 13685 64648
rect 13685 64614 13719 64648
rect 13719 64614 13740 64648
rect 13680 64600 13740 64614
rect 13260 64500 13320 64560
rect 13260 64390 13320 64450
rect 12840 64338 12900 64350
rect 12840 64304 12868 64338
rect 12868 64304 12900 64338
rect 12840 64290 12900 64304
rect 13260 64220 13320 64280
rect 13680 64338 13740 64350
rect 13680 64304 13685 64338
rect 13685 64304 13719 64338
rect 13719 64304 13740 64338
rect 13680 64290 13740 64304
rect 12840 62938 12900 62950
rect 13260 62960 13320 63020
rect 12840 62904 12868 62938
rect 12868 62904 12900 62938
rect 12840 62890 12900 62904
rect 13680 62938 13740 62950
rect 13680 62904 13685 62938
rect 13685 62904 13719 62938
rect 13719 62904 13740 62938
rect 13680 62890 13740 62904
rect 13260 62790 13320 62850
rect 13260 62680 13320 62740
rect 12840 62628 12900 62640
rect 12840 62594 12868 62628
rect 12868 62594 12900 62628
rect 12840 62580 12900 62594
rect 13260 62510 13320 62570
rect 13680 62628 13740 62640
rect 13680 62594 13685 62628
rect 13685 62594 13719 62628
rect 13719 62594 13740 62628
rect 13680 62580 13740 62594
rect 12840 61228 12900 61240
rect 13260 61250 13320 61310
rect 12840 61194 12868 61228
rect 12868 61194 12900 61228
rect 12840 61180 12900 61194
rect 13680 61228 13740 61240
rect 13680 61194 13685 61228
rect 13685 61194 13719 61228
rect 13719 61194 13740 61228
rect 13680 61180 13740 61194
rect 13260 61080 13320 61140
rect 13260 60970 13320 61030
rect 12840 60918 12900 60930
rect 12840 60884 12868 60918
rect 12868 60884 12900 60918
rect 12840 60870 12900 60884
rect 13260 60800 13320 60860
rect 13680 60918 13740 60930
rect 13680 60884 13685 60918
rect 13685 60884 13719 60918
rect 13719 60884 13740 60918
rect 13680 60870 13740 60884
rect 12840 59518 12900 59530
rect 13260 59540 13320 59600
rect 12840 59484 12868 59518
rect 12868 59484 12900 59518
rect 12840 59470 12900 59484
rect 13680 59518 13740 59530
rect 13680 59484 13685 59518
rect 13685 59484 13719 59518
rect 13719 59484 13740 59518
rect 13680 59470 13740 59484
rect 13260 59370 13320 59430
rect 13260 59260 13320 59320
rect 12840 59208 12900 59220
rect 12840 59174 12868 59208
rect 12868 59174 12900 59208
rect 12840 59160 12900 59174
rect 13260 59090 13320 59150
rect 13680 59208 13740 59220
rect 13680 59174 13685 59208
rect 13685 59174 13719 59208
rect 13719 59174 13740 59208
rect 13680 59160 13740 59174
rect 12840 57808 12900 57820
rect 13260 57830 13320 57890
rect 12840 57774 12868 57808
rect 12868 57774 12900 57808
rect 12840 57760 12900 57774
rect 13680 57808 13740 57820
rect 13680 57774 13685 57808
rect 13685 57774 13719 57808
rect 13719 57774 13740 57808
rect 13680 57760 13740 57774
rect 13260 57660 13320 57720
rect 13260 57550 13320 57610
rect 12840 57498 12900 57510
rect 12840 57464 12868 57498
rect 12868 57464 12900 57498
rect 12840 57450 12900 57464
rect 13260 57380 13320 57440
rect 13680 57498 13740 57510
rect 13680 57464 13685 57498
rect 13685 57464 13719 57498
rect 13719 57464 13740 57498
rect 13680 57450 13740 57464
rect 12840 56098 12900 56110
rect 13260 56120 13320 56180
rect 12840 56064 12868 56098
rect 12868 56064 12900 56098
rect 12840 56050 12900 56064
rect 13680 56098 13740 56110
rect 13680 56064 13685 56098
rect 13685 56064 13719 56098
rect 13719 56064 13740 56098
rect 13680 56050 13740 56064
rect 13260 55950 13320 56010
rect 13260 55840 13320 55900
rect 12840 55788 12900 55800
rect 12840 55754 12868 55788
rect 12868 55754 12900 55788
rect 12840 55740 12900 55754
rect 13260 55670 13320 55730
rect 13680 55788 13740 55800
rect 13680 55754 13685 55788
rect 13685 55754 13719 55788
rect 13719 55754 13740 55788
rect 13680 55740 13740 55754
rect 12840 54388 12900 54400
rect 13260 54410 13320 54470
rect 12840 54354 12868 54388
rect 12868 54354 12900 54388
rect 12840 54340 12900 54354
rect 13680 54388 13740 54400
rect 13680 54354 13685 54388
rect 13685 54354 13719 54388
rect 13719 54354 13740 54388
rect 13680 54340 13740 54354
rect 13260 54240 13320 54300
rect 13260 54130 13320 54190
rect 12840 54078 12900 54090
rect 12840 54044 12868 54078
rect 12868 54044 12900 54078
rect 12840 54030 12900 54044
rect 13260 53960 13320 54020
rect 13680 54078 13740 54090
rect 13680 54044 13685 54078
rect 13685 54044 13719 54078
rect 13719 54044 13740 54078
rect 13680 54030 13740 54044
rect 12840 52678 12900 52690
rect 13260 52700 13320 52760
rect 12840 52644 12868 52678
rect 12868 52644 12900 52678
rect 12840 52630 12900 52644
rect 13680 52678 13740 52690
rect 13680 52644 13685 52678
rect 13685 52644 13719 52678
rect 13719 52644 13740 52678
rect 13680 52630 13740 52644
rect 13260 52530 13320 52590
rect 13260 52420 13320 52480
rect 12840 52368 12900 52380
rect 12840 52334 12868 52368
rect 12868 52334 12900 52368
rect 12840 52320 12900 52334
rect 13260 52250 13320 52310
rect 13680 52368 13740 52380
rect 13680 52334 13685 52368
rect 13685 52334 13719 52368
rect 13719 52334 13740 52368
rect 13680 52320 13740 52334
rect 12840 50968 12900 50980
rect 13260 50990 13320 51050
rect 12840 50934 12868 50968
rect 12868 50934 12900 50968
rect 12840 50920 12900 50934
rect 13680 50968 13740 50980
rect 13680 50934 13685 50968
rect 13685 50934 13719 50968
rect 13719 50934 13740 50968
rect 13680 50920 13740 50934
rect 13260 50820 13320 50880
rect 13260 50710 13320 50770
rect 12840 50658 12900 50670
rect 12840 50624 12868 50658
rect 12868 50624 12900 50658
rect 12840 50610 12900 50624
rect 13260 50540 13320 50600
rect 13680 50658 13740 50670
rect 13680 50624 13685 50658
rect 13685 50624 13719 50658
rect 13719 50624 13740 50658
rect 13680 50610 13740 50624
rect 12840 49258 12900 49270
rect 13260 49280 13320 49340
rect 12840 49224 12868 49258
rect 12868 49224 12900 49258
rect 12840 49210 12900 49224
rect 13680 49258 13740 49270
rect 13680 49224 13685 49258
rect 13685 49224 13719 49258
rect 13719 49224 13740 49258
rect 13680 49210 13740 49224
rect 13260 49110 13320 49170
rect 13260 49000 13320 49060
rect 12840 48948 12900 48960
rect 12840 48914 12868 48948
rect 12868 48914 12900 48948
rect 12840 48900 12900 48914
rect 13260 48830 13320 48890
rect 13680 48948 13740 48960
rect 13680 48914 13685 48948
rect 13685 48914 13719 48948
rect 13719 48914 13740 48948
rect 13680 48900 13740 48914
rect 12840 47548 12900 47560
rect 13260 47570 13320 47630
rect 12840 47514 12868 47548
rect 12868 47514 12900 47548
rect 12840 47500 12900 47514
rect 13680 47548 13740 47560
rect 13680 47514 13685 47548
rect 13685 47514 13719 47548
rect 13719 47514 13740 47548
rect 13680 47500 13740 47514
rect 13260 47400 13320 47460
rect 13260 47290 13320 47350
rect 12840 47238 12900 47250
rect 12840 47204 12868 47238
rect 12868 47204 12900 47238
rect 12840 47190 12900 47204
rect 13260 47120 13320 47180
rect 13680 47238 13740 47250
rect 13680 47204 13685 47238
rect 13685 47204 13719 47238
rect 13719 47204 13740 47238
rect 13680 47190 13740 47204
rect 12840 45838 12900 45850
rect 13260 45860 13320 45920
rect 12840 45804 12868 45838
rect 12868 45804 12900 45838
rect 12840 45790 12900 45804
rect 13680 45838 13740 45850
rect 13680 45804 13685 45838
rect 13685 45804 13719 45838
rect 13719 45804 13740 45838
rect 13680 45790 13740 45804
rect 13260 45690 13320 45750
rect 13260 45580 13320 45640
rect 12840 45528 12900 45540
rect 12840 45494 12868 45528
rect 12868 45494 12900 45528
rect 12840 45480 12900 45494
rect 13260 45410 13320 45470
rect 13680 45528 13740 45540
rect 13680 45494 13685 45528
rect 13685 45494 13719 45528
rect 13719 45494 13740 45528
rect 13680 45480 13740 45494
rect 12840 44128 12900 44140
rect 13260 44150 13320 44210
rect 12840 44094 12868 44128
rect 12868 44094 12900 44128
rect 12840 44080 12900 44094
rect 13680 44128 13740 44140
rect 13680 44094 13685 44128
rect 13685 44094 13719 44128
rect 13719 44094 13740 44128
rect 13680 44080 13740 44094
rect 13260 43980 13320 44040
rect 13260 43870 13320 43930
rect 12840 43818 12900 43830
rect 12840 43784 12868 43818
rect 12868 43784 12900 43818
rect 12840 43770 12900 43784
rect 13260 43700 13320 43760
rect 13680 43818 13740 43830
rect 13680 43784 13685 43818
rect 13685 43784 13719 43818
rect 13719 43784 13740 43818
rect 13680 43770 13740 43784
rect 12840 42418 12900 42430
rect 13260 42440 13320 42500
rect 12840 42384 12868 42418
rect 12868 42384 12900 42418
rect 12840 42370 12900 42384
rect 13680 42418 13740 42430
rect 13680 42384 13685 42418
rect 13685 42384 13719 42418
rect 13719 42384 13740 42418
rect 13680 42370 13740 42384
rect 13260 42270 13320 42330
rect 13260 42160 13320 42220
rect 12840 42108 12900 42120
rect 12840 42074 12868 42108
rect 12868 42074 12900 42108
rect 12840 42060 12900 42074
rect 13260 41990 13320 42050
rect 13680 42108 13740 42120
rect 13680 42074 13685 42108
rect 13685 42074 13719 42108
rect 13719 42074 13740 42108
rect 13680 42060 13740 42074
rect 12840 40708 12900 40720
rect 13260 40730 13320 40790
rect 12840 40674 12868 40708
rect 12868 40674 12900 40708
rect 12840 40660 12900 40674
rect 13680 40708 13740 40720
rect 13680 40674 13685 40708
rect 13685 40674 13719 40708
rect 13719 40674 13740 40708
rect 13680 40660 13740 40674
rect 13260 40560 13320 40620
rect 13260 40450 13320 40510
rect 12840 40398 12900 40410
rect 12840 40364 12868 40398
rect 12868 40364 12900 40398
rect 12840 40350 12900 40364
rect 13260 40280 13320 40340
rect 13680 40398 13740 40410
rect 13680 40364 13685 40398
rect 13685 40364 13719 40398
rect 13719 40364 13740 40398
rect 13680 40350 13740 40364
rect 12730 39620 12790 39680
rect 13800 39620 13860 39680
rect 13900 66410 13960 66470
rect 13960 65880 14020 65940
rect 13900 64700 13960 64760
rect 13960 64170 14020 64230
rect 13900 62990 13960 63050
rect 13960 62460 14020 62520
rect 13900 61280 13960 61340
rect 13960 60750 14020 60810
rect 13900 59570 13960 59630
rect 13960 59040 14020 59100
rect 13900 57860 13960 57920
rect 13960 57330 14020 57390
rect 13900 56150 13960 56210
rect 13960 55620 14020 55680
rect 13900 54440 13960 54500
rect 13960 53910 14020 53970
rect 13900 52730 13960 52790
rect 13960 52200 14020 52260
rect 13900 51020 13960 51080
rect 13960 50490 14020 50550
rect 13900 49310 13960 49370
rect 13960 48780 14020 48840
rect 13900 47600 13960 47660
rect 13960 47070 14020 47130
rect 13900 45890 13960 45950
rect 13960 45360 14020 45420
rect 13900 44180 13960 44240
rect 13960 43650 14020 43710
rect 13900 42470 13960 42530
rect 13960 41940 14020 42000
rect 13900 40760 13960 40820
rect 12430 39170 12490 39230
rect 13960 40230 14020 40290
rect 13960 39620 14020 39680
rect 14050 66320 14110 66380
rect 14050 64610 14110 64670
rect 14050 62900 14110 62960
rect 14050 61190 14110 61250
rect 14170 59480 14230 59540
rect 14170 57770 14230 57830
rect 14170 56060 14230 56120
rect 14170 54350 14230 54410
rect 14170 52640 14230 52700
rect 14170 50930 14230 50990
rect 14170 49220 14230 49280
rect 14170 47510 14230 47570
rect 14050 45800 14110 45860
rect 14050 44090 14110 44150
rect 14050 42380 14110 42440
rect 14050 40670 14110 40730
rect 17620 66320 17680 66380
rect 17620 64610 17680 64670
rect 17620 62900 17680 62960
rect 17620 61190 17680 61250
rect 17500 59480 17560 59540
rect 17500 57770 17560 57830
rect 17500 56060 17560 56120
rect 17500 54350 17560 54410
rect 17500 52640 17560 52700
rect 17500 50930 17560 50990
rect 17500 49220 17560 49280
rect 17500 47510 17560 47570
rect 17620 45800 17680 45860
rect 17620 44090 17680 44150
rect 17620 42380 17680 42440
rect 17620 40670 17680 40730
rect 14250 39170 14310 39230
rect 14430 39230 14490 39290
rect 17240 39230 17300 39290
rect 17830 66358 17890 66370
rect 18250 66380 18310 66440
rect 17830 66324 17858 66358
rect 17858 66324 17890 66358
rect 17830 66310 17890 66324
rect 18670 66358 18730 66370
rect 18670 66324 18675 66358
rect 18675 66324 18709 66358
rect 18709 66324 18730 66358
rect 18670 66310 18730 66324
rect 18250 66210 18310 66270
rect 18250 66100 18310 66160
rect 17830 66048 17890 66060
rect 17830 66014 17858 66048
rect 17858 66014 17890 66048
rect 17830 66000 17890 66014
rect 18250 65930 18310 65990
rect 18670 66048 18730 66060
rect 18670 66014 18675 66048
rect 18675 66014 18709 66048
rect 18709 66014 18730 66048
rect 18670 66000 18730 66014
rect 17830 64648 17890 64660
rect 18250 64670 18310 64730
rect 17830 64614 17858 64648
rect 17858 64614 17890 64648
rect 17830 64600 17890 64614
rect 18670 64648 18730 64660
rect 18670 64614 18675 64648
rect 18675 64614 18709 64648
rect 18709 64614 18730 64648
rect 18670 64600 18730 64614
rect 18250 64500 18310 64560
rect 18250 64390 18310 64450
rect 17830 64338 17890 64350
rect 17830 64304 17858 64338
rect 17858 64304 17890 64338
rect 17830 64290 17890 64304
rect 18250 64220 18310 64280
rect 18670 64338 18730 64350
rect 18670 64304 18675 64338
rect 18675 64304 18709 64338
rect 18709 64304 18730 64338
rect 18670 64290 18730 64304
rect 17830 62938 17890 62950
rect 18250 62960 18310 63020
rect 17830 62904 17858 62938
rect 17858 62904 17890 62938
rect 17830 62890 17890 62904
rect 18670 62938 18730 62950
rect 18670 62904 18675 62938
rect 18675 62904 18709 62938
rect 18709 62904 18730 62938
rect 18670 62890 18730 62904
rect 18250 62790 18310 62850
rect 18250 62680 18310 62740
rect 17830 62628 17890 62640
rect 17830 62594 17858 62628
rect 17858 62594 17890 62628
rect 17830 62580 17890 62594
rect 18250 62510 18310 62570
rect 18670 62628 18730 62640
rect 18670 62594 18675 62628
rect 18675 62594 18709 62628
rect 18709 62594 18730 62628
rect 18670 62580 18730 62594
rect 17830 61228 17890 61240
rect 18250 61250 18310 61310
rect 17830 61194 17858 61228
rect 17858 61194 17890 61228
rect 17830 61180 17890 61194
rect 18670 61228 18730 61240
rect 18670 61194 18675 61228
rect 18675 61194 18709 61228
rect 18709 61194 18730 61228
rect 18670 61180 18730 61194
rect 18250 61080 18310 61140
rect 18250 60970 18310 61030
rect 17830 60918 17890 60930
rect 17830 60884 17858 60918
rect 17858 60884 17890 60918
rect 17830 60870 17890 60884
rect 18250 60800 18310 60860
rect 18670 60918 18730 60930
rect 18670 60884 18675 60918
rect 18675 60884 18709 60918
rect 18709 60884 18730 60918
rect 18670 60870 18730 60884
rect 17830 59518 17890 59530
rect 18250 59540 18310 59600
rect 17830 59484 17858 59518
rect 17858 59484 17890 59518
rect 17830 59470 17890 59484
rect 18670 59518 18730 59530
rect 18670 59484 18675 59518
rect 18675 59484 18709 59518
rect 18709 59484 18730 59518
rect 18670 59470 18730 59484
rect 18250 59370 18310 59430
rect 18250 59260 18310 59320
rect 17830 59208 17890 59220
rect 17830 59174 17858 59208
rect 17858 59174 17890 59208
rect 17830 59160 17890 59174
rect 18250 59090 18310 59150
rect 18670 59208 18730 59220
rect 18670 59174 18675 59208
rect 18675 59174 18709 59208
rect 18709 59174 18730 59208
rect 18670 59160 18730 59174
rect 17830 57808 17890 57820
rect 18250 57830 18310 57890
rect 17830 57774 17858 57808
rect 17858 57774 17890 57808
rect 17830 57760 17890 57774
rect 18670 57808 18730 57820
rect 18670 57774 18675 57808
rect 18675 57774 18709 57808
rect 18709 57774 18730 57808
rect 18670 57760 18730 57774
rect 18250 57660 18310 57720
rect 18250 57550 18310 57610
rect 17830 57498 17890 57510
rect 17830 57464 17858 57498
rect 17858 57464 17890 57498
rect 17830 57450 17890 57464
rect 18250 57380 18310 57440
rect 18670 57498 18730 57510
rect 18670 57464 18675 57498
rect 18675 57464 18709 57498
rect 18709 57464 18730 57498
rect 18670 57450 18730 57464
rect 17830 56098 17890 56110
rect 18250 56120 18310 56180
rect 17830 56064 17858 56098
rect 17858 56064 17890 56098
rect 17830 56050 17890 56064
rect 18670 56098 18730 56110
rect 18670 56064 18675 56098
rect 18675 56064 18709 56098
rect 18709 56064 18730 56098
rect 18670 56050 18730 56064
rect 18250 55950 18310 56010
rect 18250 55840 18310 55900
rect 17830 55788 17890 55800
rect 17830 55754 17858 55788
rect 17858 55754 17890 55788
rect 17830 55740 17890 55754
rect 18250 55670 18310 55730
rect 18670 55788 18730 55800
rect 18670 55754 18675 55788
rect 18675 55754 18709 55788
rect 18709 55754 18730 55788
rect 18670 55740 18730 55754
rect 17830 54388 17890 54400
rect 18250 54410 18310 54470
rect 17830 54354 17858 54388
rect 17858 54354 17890 54388
rect 17830 54340 17890 54354
rect 18670 54388 18730 54400
rect 18670 54354 18675 54388
rect 18675 54354 18709 54388
rect 18709 54354 18730 54388
rect 18670 54340 18730 54354
rect 18250 54240 18310 54300
rect 18250 54130 18310 54190
rect 17830 54078 17890 54090
rect 17830 54044 17858 54078
rect 17858 54044 17890 54078
rect 17830 54030 17890 54044
rect 18250 53960 18310 54020
rect 18670 54078 18730 54090
rect 18670 54044 18675 54078
rect 18675 54044 18709 54078
rect 18709 54044 18730 54078
rect 18670 54030 18730 54044
rect 17830 52678 17890 52690
rect 18250 52700 18310 52760
rect 17830 52644 17858 52678
rect 17858 52644 17890 52678
rect 17830 52630 17890 52644
rect 18670 52678 18730 52690
rect 18670 52644 18675 52678
rect 18675 52644 18709 52678
rect 18709 52644 18730 52678
rect 18670 52630 18730 52644
rect 18250 52530 18310 52590
rect 18250 52420 18310 52480
rect 17830 52368 17890 52380
rect 17830 52334 17858 52368
rect 17858 52334 17890 52368
rect 17830 52320 17890 52334
rect 18250 52250 18310 52310
rect 18670 52368 18730 52380
rect 18670 52334 18675 52368
rect 18675 52334 18709 52368
rect 18709 52334 18730 52368
rect 18670 52320 18730 52334
rect 17830 50968 17890 50980
rect 18250 50990 18310 51050
rect 17830 50934 17858 50968
rect 17858 50934 17890 50968
rect 17830 50920 17890 50934
rect 18670 50968 18730 50980
rect 18670 50934 18675 50968
rect 18675 50934 18709 50968
rect 18709 50934 18730 50968
rect 18670 50920 18730 50934
rect 18250 50820 18310 50880
rect 18250 50710 18310 50770
rect 17830 50658 17890 50670
rect 17830 50624 17858 50658
rect 17858 50624 17890 50658
rect 17830 50610 17890 50624
rect 18250 50540 18310 50600
rect 18670 50658 18730 50670
rect 18670 50624 18675 50658
rect 18675 50624 18709 50658
rect 18709 50624 18730 50658
rect 18670 50610 18730 50624
rect 17830 49258 17890 49270
rect 18250 49280 18310 49340
rect 17830 49224 17858 49258
rect 17858 49224 17890 49258
rect 17830 49210 17890 49224
rect 18670 49258 18730 49270
rect 18670 49224 18675 49258
rect 18675 49224 18709 49258
rect 18709 49224 18730 49258
rect 18670 49210 18730 49224
rect 18250 49110 18310 49170
rect 18250 49000 18310 49060
rect 17830 48948 17890 48960
rect 17830 48914 17858 48948
rect 17858 48914 17890 48948
rect 17830 48900 17890 48914
rect 18250 48830 18310 48890
rect 18670 48948 18730 48960
rect 18670 48914 18675 48948
rect 18675 48914 18709 48948
rect 18709 48914 18730 48948
rect 18670 48900 18730 48914
rect 17830 47548 17890 47560
rect 18250 47570 18310 47630
rect 17830 47514 17858 47548
rect 17858 47514 17890 47548
rect 17830 47500 17890 47514
rect 18670 47548 18730 47560
rect 18670 47514 18675 47548
rect 18675 47514 18709 47548
rect 18709 47514 18730 47548
rect 18670 47500 18730 47514
rect 18250 47400 18310 47460
rect 18250 47290 18310 47350
rect 17830 47238 17890 47250
rect 17830 47204 17858 47238
rect 17858 47204 17890 47238
rect 17830 47190 17890 47204
rect 18250 47120 18310 47180
rect 18670 47238 18730 47250
rect 18670 47204 18675 47238
rect 18675 47204 18709 47238
rect 18709 47204 18730 47238
rect 18670 47190 18730 47204
rect 17830 45838 17890 45850
rect 18250 45860 18310 45920
rect 17830 45804 17858 45838
rect 17858 45804 17890 45838
rect 17830 45790 17890 45804
rect 18670 45838 18730 45850
rect 18670 45804 18675 45838
rect 18675 45804 18709 45838
rect 18709 45804 18730 45838
rect 18670 45790 18730 45804
rect 18250 45690 18310 45750
rect 18250 45580 18310 45640
rect 17830 45528 17890 45540
rect 17830 45494 17858 45528
rect 17858 45494 17890 45528
rect 17830 45480 17890 45494
rect 18250 45410 18310 45470
rect 18670 45528 18730 45540
rect 18670 45494 18675 45528
rect 18675 45494 18709 45528
rect 18709 45494 18730 45528
rect 18670 45480 18730 45494
rect 17830 44128 17890 44140
rect 18250 44150 18310 44210
rect 17830 44094 17858 44128
rect 17858 44094 17890 44128
rect 17830 44080 17890 44094
rect 18670 44128 18730 44140
rect 18670 44094 18675 44128
rect 18675 44094 18709 44128
rect 18709 44094 18730 44128
rect 18670 44080 18730 44094
rect 18250 43980 18310 44040
rect 18250 43870 18310 43930
rect 17830 43818 17890 43830
rect 17830 43784 17858 43818
rect 17858 43784 17890 43818
rect 17830 43770 17890 43784
rect 18250 43700 18310 43760
rect 18670 43818 18730 43830
rect 18670 43784 18675 43818
rect 18675 43784 18709 43818
rect 18709 43784 18730 43818
rect 18670 43770 18730 43784
rect 17830 42418 17890 42430
rect 18250 42440 18310 42500
rect 17830 42384 17858 42418
rect 17858 42384 17890 42418
rect 17830 42370 17890 42384
rect 18670 42418 18730 42430
rect 18670 42384 18675 42418
rect 18675 42384 18709 42418
rect 18709 42384 18730 42418
rect 18670 42370 18730 42384
rect 18250 42270 18310 42330
rect 18250 42160 18310 42220
rect 17830 42108 17890 42120
rect 17830 42074 17858 42108
rect 17858 42074 17890 42108
rect 17830 42060 17890 42074
rect 18250 41990 18310 42050
rect 18670 42108 18730 42120
rect 18670 42074 18675 42108
rect 18675 42074 18709 42108
rect 18709 42074 18730 42108
rect 18670 42060 18730 42074
rect 17830 40708 17890 40720
rect 18250 40730 18310 40790
rect 17830 40674 17858 40708
rect 17858 40674 17890 40708
rect 17830 40660 17890 40674
rect 18670 40708 18730 40720
rect 18670 40674 18675 40708
rect 18675 40674 18709 40708
rect 18709 40674 18730 40708
rect 18670 40660 18730 40674
rect 18250 40560 18310 40620
rect 18250 40450 18310 40510
rect 17830 40398 17890 40410
rect 17830 40364 17858 40398
rect 17858 40364 17890 40398
rect 17830 40350 17890 40364
rect 18250 40280 18310 40340
rect 18670 40398 18730 40410
rect 18670 40364 18675 40398
rect 18675 40364 18709 40398
rect 18709 40364 18730 40398
rect 18670 40350 18730 40364
rect 17720 39620 17780 39680
rect 18790 39620 18850 39680
rect 18890 66410 18950 66470
rect 18950 65880 19010 65940
rect 18890 64700 18950 64760
rect 18950 64170 19010 64230
rect 18890 62990 18950 63050
rect 18950 62460 19010 62520
rect 18890 61280 18950 61340
rect 18950 60750 19010 60810
rect 18890 59570 18950 59630
rect 18950 59040 19010 59100
rect 18890 57860 18950 57920
rect 18950 57330 19010 57390
rect 18890 56150 18950 56210
rect 18950 55620 19010 55680
rect 18890 54440 18950 54500
rect 18950 53910 19010 53970
rect 18890 52730 18950 52790
rect 18950 52200 19010 52260
rect 18890 51020 18950 51080
rect 18950 50490 19010 50550
rect 18890 49310 18950 49370
rect 18950 48780 19010 48840
rect 18890 47600 18950 47660
rect 18950 47070 19010 47130
rect 18890 45890 18950 45950
rect 18950 45360 19010 45420
rect 18890 44180 18950 44240
rect 18950 43650 19010 43710
rect 18890 42470 18950 42530
rect 18950 41940 19010 42000
rect 18890 40760 18950 40820
rect 17420 39170 17480 39230
rect 18950 40230 19010 40290
rect 18950 39620 19010 39680
rect 19040 66320 19100 66380
rect 19040 64610 19100 64670
rect 19040 62900 19100 62960
rect 19040 61190 19100 61250
rect 19160 59480 19220 59540
rect 19160 57770 19220 57830
rect 19160 56060 19220 56120
rect 19160 54350 19220 54410
rect 19160 52640 19220 52700
rect 19160 50930 19220 50990
rect 19160 49220 19220 49280
rect 19160 47510 19220 47570
rect 19040 45800 19100 45860
rect 19040 44090 19100 44150
rect 19040 42380 19100 42440
rect 19040 40670 19100 40730
rect 22610 66320 22670 66380
rect 22610 64610 22670 64670
rect 22490 62900 22550 62960
rect 22490 61180 22550 61240
rect 22370 59480 22430 59540
rect 22250 57770 22310 57830
rect 22250 56060 22310 56120
rect 22250 54350 22310 54410
rect 22250 52640 22310 52700
rect 22250 50930 22310 50990
rect 22250 49220 22310 49280
rect 22370 47510 22430 47570
rect 21870 39350 21930 39410
rect 22490 45800 22550 45860
rect 22490 44090 22550 44150
rect 19240 39170 19300 39230
rect 19420 39230 19480 39290
rect 22050 39290 22110 39350
rect 22610 42380 22670 42440
rect 22610 40670 22670 40730
rect 22230 39230 22290 39290
rect 22820 66358 22880 66370
rect 23240 66380 23300 66440
rect 22820 66324 22848 66358
rect 22848 66324 22880 66358
rect 22820 66310 22880 66324
rect 23660 66358 23720 66370
rect 23660 66324 23665 66358
rect 23665 66324 23699 66358
rect 23699 66324 23720 66358
rect 23660 66310 23720 66324
rect 23240 66210 23300 66270
rect 23240 66100 23300 66160
rect 22820 66048 22880 66060
rect 22820 66014 22848 66048
rect 22848 66014 22880 66048
rect 22820 66000 22880 66014
rect 23240 65930 23300 65990
rect 23660 66048 23720 66060
rect 23660 66014 23665 66048
rect 23665 66014 23699 66048
rect 23699 66014 23720 66048
rect 23660 66000 23720 66014
rect 22820 64648 22880 64660
rect 23240 64670 23300 64730
rect 22820 64614 22848 64648
rect 22848 64614 22880 64648
rect 22820 64600 22880 64614
rect 23660 64648 23720 64660
rect 23660 64614 23665 64648
rect 23665 64614 23699 64648
rect 23699 64614 23720 64648
rect 23660 64600 23720 64614
rect 23240 64500 23300 64560
rect 23240 64390 23300 64450
rect 22820 64338 22880 64350
rect 22820 64304 22848 64338
rect 22848 64304 22880 64338
rect 22820 64290 22880 64304
rect 23240 64220 23300 64280
rect 23660 64338 23720 64350
rect 23660 64304 23665 64338
rect 23665 64304 23699 64338
rect 23699 64304 23720 64338
rect 23660 64290 23720 64304
rect 22820 62938 22880 62950
rect 23240 62960 23300 63020
rect 22820 62904 22848 62938
rect 22848 62904 22880 62938
rect 22820 62890 22880 62904
rect 23660 62938 23720 62950
rect 23660 62904 23665 62938
rect 23665 62904 23699 62938
rect 23699 62904 23720 62938
rect 23660 62890 23720 62904
rect 23240 62790 23300 62850
rect 23240 62680 23300 62740
rect 22820 62628 22880 62640
rect 22820 62594 22848 62628
rect 22848 62594 22880 62628
rect 22820 62580 22880 62594
rect 23240 62510 23300 62570
rect 23660 62628 23720 62640
rect 23660 62594 23665 62628
rect 23665 62594 23699 62628
rect 23699 62594 23720 62628
rect 23660 62580 23720 62594
rect 22820 61228 22880 61240
rect 23240 61250 23300 61310
rect 22820 61194 22848 61228
rect 22848 61194 22880 61228
rect 22820 61180 22880 61194
rect 23660 61228 23720 61240
rect 23660 61194 23665 61228
rect 23665 61194 23699 61228
rect 23699 61194 23720 61228
rect 23660 61180 23720 61194
rect 23240 61080 23300 61140
rect 23240 60970 23300 61030
rect 22820 60918 22880 60930
rect 22820 60884 22848 60918
rect 22848 60884 22880 60918
rect 22820 60870 22880 60884
rect 23240 60800 23300 60860
rect 23660 60918 23720 60930
rect 23660 60884 23665 60918
rect 23665 60884 23699 60918
rect 23699 60884 23720 60918
rect 23660 60870 23720 60884
rect 22820 59518 22880 59530
rect 23240 59540 23300 59600
rect 22820 59484 22848 59518
rect 22848 59484 22880 59518
rect 22820 59470 22880 59484
rect 23660 59518 23720 59530
rect 23660 59484 23665 59518
rect 23665 59484 23699 59518
rect 23699 59484 23720 59518
rect 23660 59470 23720 59484
rect 23240 59370 23300 59430
rect 23240 59260 23300 59320
rect 22820 59208 22880 59220
rect 22820 59174 22848 59208
rect 22848 59174 22880 59208
rect 22820 59160 22880 59174
rect 23240 59090 23300 59150
rect 23660 59208 23720 59220
rect 23660 59174 23665 59208
rect 23665 59174 23699 59208
rect 23699 59174 23720 59208
rect 23660 59160 23720 59174
rect 22820 57808 22880 57820
rect 23240 57830 23300 57890
rect 22820 57774 22848 57808
rect 22848 57774 22880 57808
rect 22820 57760 22880 57774
rect 23660 57808 23720 57820
rect 23660 57774 23665 57808
rect 23665 57774 23699 57808
rect 23699 57774 23720 57808
rect 23660 57760 23720 57774
rect 23240 57660 23300 57720
rect 23240 57550 23300 57610
rect 22820 57498 22880 57510
rect 22820 57464 22848 57498
rect 22848 57464 22880 57498
rect 22820 57450 22880 57464
rect 23240 57380 23300 57440
rect 23660 57498 23720 57510
rect 23660 57464 23665 57498
rect 23665 57464 23699 57498
rect 23699 57464 23720 57498
rect 23660 57450 23720 57464
rect 22820 56098 22880 56110
rect 23240 56120 23300 56180
rect 22820 56064 22848 56098
rect 22848 56064 22880 56098
rect 22820 56050 22880 56064
rect 23660 56098 23720 56110
rect 23660 56064 23665 56098
rect 23665 56064 23699 56098
rect 23699 56064 23720 56098
rect 23660 56050 23720 56064
rect 23240 55950 23300 56010
rect 23240 55840 23300 55900
rect 22820 55788 22880 55800
rect 22820 55754 22848 55788
rect 22848 55754 22880 55788
rect 22820 55740 22880 55754
rect 23240 55670 23300 55730
rect 23660 55788 23720 55800
rect 23660 55754 23665 55788
rect 23665 55754 23699 55788
rect 23699 55754 23720 55788
rect 23660 55740 23720 55754
rect 22820 54388 22880 54400
rect 23240 54410 23300 54470
rect 22820 54354 22848 54388
rect 22848 54354 22880 54388
rect 22820 54340 22880 54354
rect 23660 54388 23720 54400
rect 23660 54354 23665 54388
rect 23665 54354 23699 54388
rect 23699 54354 23720 54388
rect 23660 54340 23720 54354
rect 23240 54240 23300 54300
rect 23240 54130 23300 54190
rect 22820 54078 22880 54090
rect 22820 54044 22848 54078
rect 22848 54044 22880 54078
rect 22820 54030 22880 54044
rect 23240 53960 23300 54020
rect 23660 54078 23720 54090
rect 23660 54044 23665 54078
rect 23665 54044 23699 54078
rect 23699 54044 23720 54078
rect 23660 54030 23720 54044
rect 22820 52678 22880 52690
rect 23240 52700 23300 52760
rect 22820 52644 22848 52678
rect 22848 52644 22880 52678
rect 22820 52630 22880 52644
rect 23660 52678 23720 52690
rect 23660 52644 23665 52678
rect 23665 52644 23699 52678
rect 23699 52644 23720 52678
rect 23660 52630 23720 52644
rect 23240 52530 23300 52590
rect 23240 52420 23300 52480
rect 22820 52368 22880 52380
rect 22820 52334 22848 52368
rect 22848 52334 22880 52368
rect 22820 52320 22880 52334
rect 23240 52250 23300 52310
rect 23660 52368 23720 52380
rect 23660 52334 23665 52368
rect 23665 52334 23699 52368
rect 23699 52334 23720 52368
rect 23660 52320 23720 52334
rect 22820 50968 22880 50980
rect 23240 50990 23300 51050
rect 22820 50934 22848 50968
rect 22848 50934 22880 50968
rect 22820 50920 22880 50934
rect 23660 50968 23720 50980
rect 23660 50934 23665 50968
rect 23665 50934 23699 50968
rect 23699 50934 23720 50968
rect 23660 50920 23720 50934
rect 23240 50820 23300 50880
rect 23240 50710 23300 50770
rect 22820 50658 22880 50670
rect 22820 50624 22848 50658
rect 22848 50624 22880 50658
rect 22820 50610 22880 50624
rect 23240 50540 23300 50600
rect 23660 50658 23720 50670
rect 23660 50624 23665 50658
rect 23665 50624 23699 50658
rect 23699 50624 23720 50658
rect 23660 50610 23720 50624
rect 22820 49258 22880 49270
rect 23240 49280 23300 49340
rect 22820 49224 22848 49258
rect 22848 49224 22880 49258
rect 22820 49210 22880 49224
rect 23660 49258 23720 49270
rect 23660 49224 23665 49258
rect 23665 49224 23699 49258
rect 23699 49224 23720 49258
rect 23660 49210 23720 49224
rect 23240 49110 23300 49170
rect 23240 49000 23300 49060
rect 22820 48948 22880 48960
rect 22820 48914 22848 48948
rect 22848 48914 22880 48948
rect 22820 48900 22880 48914
rect 23240 48830 23300 48890
rect 23660 48948 23720 48960
rect 23660 48914 23665 48948
rect 23665 48914 23699 48948
rect 23699 48914 23720 48948
rect 23660 48900 23720 48914
rect 22820 47548 22880 47560
rect 23240 47570 23300 47630
rect 22820 47514 22848 47548
rect 22848 47514 22880 47548
rect 22820 47500 22880 47514
rect 23660 47548 23720 47560
rect 23660 47514 23665 47548
rect 23665 47514 23699 47548
rect 23699 47514 23720 47548
rect 23660 47500 23720 47514
rect 23240 47400 23300 47460
rect 23240 47290 23300 47350
rect 22820 47238 22880 47250
rect 22820 47204 22848 47238
rect 22848 47204 22880 47238
rect 22820 47190 22880 47204
rect 23240 47120 23300 47180
rect 23660 47238 23720 47250
rect 23660 47204 23665 47238
rect 23665 47204 23699 47238
rect 23699 47204 23720 47238
rect 23660 47190 23720 47204
rect 22820 45838 22880 45850
rect 23240 45860 23300 45920
rect 22820 45804 22848 45838
rect 22848 45804 22880 45838
rect 22820 45790 22880 45804
rect 23660 45838 23720 45850
rect 23660 45804 23665 45838
rect 23665 45804 23699 45838
rect 23699 45804 23720 45838
rect 23660 45790 23720 45804
rect 23240 45690 23300 45750
rect 23240 45580 23300 45640
rect 22820 45528 22880 45540
rect 22820 45494 22848 45528
rect 22848 45494 22880 45528
rect 22820 45480 22880 45494
rect 23240 45410 23300 45470
rect 23660 45528 23720 45540
rect 23660 45494 23665 45528
rect 23665 45494 23699 45528
rect 23699 45494 23720 45528
rect 23660 45480 23720 45494
rect 22820 44128 22880 44140
rect 23240 44150 23300 44210
rect 22820 44094 22848 44128
rect 22848 44094 22880 44128
rect 22820 44080 22880 44094
rect 23660 44128 23720 44140
rect 23660 44094 23665 44128
rect 23665 44094 23699 44128
rect 23699 44094 23720 44128
rect 23660 44080 23720 44094
rect 23240 43980 23300 44040
rect 23240 43870 23300 43930
rect 22820 43818 22880 43830
rect 22820 43784 22848 43818
rect 22848 43784 22880 43818
rect 22820 43770 22880 43784
rect 23240 43700 23300 43760
rect 23660 43818 23720 43830
rect 23660 43784 23665 43818
rect 23665 43784 23699 43818
rect 23699 43784 23720 43818
rect 23660 43770 23720 43784
rect 22820 42418 22880 42430
rect 23240 42440 23300 42500
rect 22820 42384 22848 42418
rect 22848 42384 22880 42418
rect 22820 42370 22880 42384
rect 23660 42418 23720 42430
rect 23660 42384 23665 42418
rect 23665 42384 23699 42418
rect 23699 42384 23720 42418
rect 23660 42370 23720 42384
rect 23240 42270 23300 42330
rect 23240 42160 23300 42220
rect 22820 42108 22880 42120
rect 22820 42074 22848 42108
rect 22848 42074 22880 42108
rect 22820 42060 22880 42074
rect 23240 41990 23300 42050
rect 23660 42108 23720 42120
rect 23660 42074 23665 42108
rect 23665 42074 23699 42108
rect 23699 42074 23720 42108
rect 23660 42060 23720 42074
rect 22820 40708 22880 40720
rect 23240 40730 23300 40790
rect 22820 40674 22848 40708
rect 22848 40674 22880 40708
rect 22820 40660 22880 40674
rect 23660 40708 23720 40720
rect 23660 40674 23665 40708
rect 23665 40674 23699 40708
rect 23699 40674 23720 40708
rect 23660 40660 23720 40674
rect 23240 40560 23300 40620
rect 23240 40450 23300 40510
rect 22820 40398 22880 40410
rect 22820 40364 22848 40398
rect 22848 40364 22880 40398
rect 22820 40350 22880 40364
rect 23240 40280 23300 40340
rect 23660 40398 23720 40410
rect 23660 40364 23665 40398
rect 23665 40364 23699 40398
rect 23699 40364 23720 40398
rect 23660 40350 23720 40364
rect 22710 39620 22770 39680
rect 23780 39620 23840 39680
rect 23880 66410 23940 66470
rect 23940 65880 24000 65940
rect 23880 64700 23940 64760
rect 23940 64170 24000 64230
rect 23880 62990 23940 63050
rect 23940 62460 24000 62520
rect 23880 61280 23940 61340
rect 23940 60750 24000 60810
rect 23880 59570 23940 59630
rect 23940 59040 24000 59100
rect 23880 57860 23940 57920
rect 23940 57330 24000 57390
rect 23880 56150 23940 56210
rect 23940 55620 24000 55680
rect 23880 54440 23940 54500
rect 23940 53910 24000 53970
rect 23880 52730 23940 52790
rect 23940 52200 24000 52260
rect 23880 51020 23940 51080
rect 23940 50490 24000 50550
rect 23880 49310 23940 49370
rect 23940 48780 24000 48840
rect 23880 47600 23940 47660
rect 23940 47070 24000 47130
rect 23880 45890 23940 45950
rect 23940 45360 24000 45420
rect 23880 44180 23940 44240
rect 23940 43650 24000 43710
rect 23880 42470 23940 42530
rect 23940 41940 24000 42000
rect 23880 40760 23940 40820
rect 22410 39170 22470 39230
rect 23940 40230 24000 40290
rect 23940 39620 24000 39680
rect 24030 66320 24090 66380
rect 24030 64610 24090 64670
rect 24150 62900 24210 62960
rect 24150 61180 24210 61240
rect 24270 59480 24330 59540
rect 24390 57770 24450 57830
rect 24390 56060 24450 56120
rect 24390 54350 24450 54410
rect 24390 52640 24450 52700
rect 24390 50930 24450 50990
rect 24390 49220 24450 49280
rect 24270 47510 24330 47570
rect 24150 45800 24210 45860
rect 24150 44090 24210 44150
rect 24030 42380 24090 42440
rect 24030 40670 24090 40730
rect 27600 66320 27660 66380
rect 27600 64610 27660 64670
rect 27480 62900 27540 62960
rect 27480 61180 27540 61240
rect 27360 59480 27420 59540
rect 27240 57770 27300 57830
rect 27240 56060 27300 56120
rect 27240 54350 27300 54410
rect 27240 52640 27300 52700
rect 27240 50930 27300 50990
rect 27240 49220 27300 49280
rect 27360 47510 27420 47570
rect 24230 39170 24290 39230
rect 24410 39230 24470 39290
rect 24590 39290 24650 39350
rect 24770 39350 24830 39410
rect 26860 39350 26920 39410
rect 27480 45800 27540 45860
rect 27480 44090 27540 44150
rect 27040 39290 27100 39350
rect 27600 42380 27660 42440
rect 27600 40670 27660 40730
rect 27220 39230 27280 39290
rect 27810 66358 27870 66370
rect 28230 66380 28290 66440
rect 27810 66324 27838 66358
rect 27838 66324 27870 66358
rect 27810 66310 27870 66324
rect 28650 66358 28710 66370
rect 28650 66324 28655 66358
rect 28655 66324 28689 66358
rect 28689 66324 28710 66358
rect 28650 66310 28710 66324
rect 28230 66210 28290 66270
rect 28230 66100 28290 66160
rect 27810 66048 27870 66060
rect 27810 66014 27838 66048
rect 27838 66014 27870 66048
rect 27810 66000 27870 66014
rect 28230 65930 28290 65990
rect 28650 66048 28710 66060
rect 28650 66014 28655 66048
rect 28655 66014 28689 66048
rect 28689 66014 28710 66048
rect 28650 66000 28710 66014
rect 27810 64648 27870 64660
rect 28230 64670 28290 64730
rect 27810 64614 27838 64648
rect 27838 64614 27870 64648
rect 27810 64600 27870 64614
rect 28650 64648 28710 64660
rect 28650 64614 28655 64648
rect 28655 64614 28689 64648
rect 28689 64614 28710 64648
rect 28650 64600 28710 64614
rect 28230 64500 28290 64560
rect 28230 64390 28290 64450
rect 27810 64338 27870 64350
rect 27810 64304 27838 64338
rect 27838 64304 27870 64338
rect 27810 64290 27870 64304
rect 28230 64220 28290 64280
rect 28650 64338 28710 64350
rect 28650 64304 28655 64338
rect 28655 64304 28689 64338
rect 28689 64304 28710 64338
rect 28650 64290 28710 64304
rect 27810 62938 27870 62950
rect 28230 62960 28290 63020
rect 27810 62904 27838 62938
rect 27838 62904 27870 62938
rect 27810 62890 27870 62904
rect 28650 62938 28710 62950
rect 28650 62904 28655 62938
rect 28655 62904 28689 62938
rect 28689 62904 28710 62938
rect 28650 62890 28710 62904
rect 28230 62790 28290 62850
rect 28230 62680 28290 62740
rect 27810 62628 27870 62640
rect 27810 62594 27838 62628
rect 27838 62594 27870 62628
rect 27810 62580 27870 62594
rect 28230 62510 28290 62570
rect 28650 62628 28710 62640
rect 28650 62594 28655 62628
rect 28655 62594 28689 62628
rect 28689 62594 28710 62628
rect 28650 62580 28710 62594
rect 27810 61228 27870 61240
rect 28230 61250 28290 61310
rect 27810 61194 27838 61228
rect 27838 61194 27870 61228
rect 27810 61180 27870 61194
rect 28650 61228 28710 61240
rect 28650 61194 28655 61228
rect 28655 61194 28689 61228
rect 28689 61194 28710 61228
rect 28650 61180 28710 61194
rect 28230 61080 28290 61140
rect 28230 60970 28290 61030
rect 27810 60918 27870 60930
rect 27810 60884 27838 60918
rect 27838 60884 27870 60918
rect 27810 60870 27870 60884
rect 28230 60800 28290 60860
rect 28650 60918 28710 60930
rect 28650 60884 28655 60918
rect 28655 60884 28689 60918
rect 28689 60884 28710 60918
rect 28650 60870 28710 60884
rect 27810 59518 27870 59530
rect 28230 59540 28290 59600
rect 27810 59484 27838 59518
rect 27838 59484 27870 59518
rect 27810 59470 27870 59484
rect 28650 59518 28710 59530
rect 28650 59484 28655 59518
rect 28655 59484 28689 59518
rect 28689 59484 28710 59518
rect 28650 59470 28710 59484
rect 28230 59370 28290 59430
rect 28230 59260 28290 59320
rect 27810 59208 27870 59220
rect 27810 59174 27838 59208
rect 27838 59174 27870 59208
rect 27810 59160 27870 59174
rect 28230 59090 28290 59150
rect 28650 59208 28710 59220
rect 28650 59174 28655 59208
rect 28655 59174 28689 59208
rect 28689 59174 28710 59208
rect 28650 59160 28710 59174
rect 27810 57808 27870 57820
rect 28230 57830 28290 57890
rect 27810 57774 27838 57808
rect 27838 57774 27870 57808
rect 27810 57760 27870 57774
rect 28650 57808 28710 57820
rect 28650 57774 28655 57808
rect 28655 57774 28689 57808
rect 28689 57774 28710 57808
rect 28650 57760 28710 57774
rect 28230 57660 28290 57720
rect 28230 57550 28290 57610
rect 27810 57498 27870 57510
rect 27810 57464 27838 57498
rect 27838 57464 27870 57498
rect 27810 57450 27870 57464
rect 28230 57380 28290 57440
rect 28650 57498 28710 57510
rect 28650 57464 28655 57498
rect 28655 57464 28689 57498
rect 28689 57464 28710 57498
rect 28650 57450 28710 57464
rect 27810 56098 27870 56110
rect 28230 56120 28290 56180
rect 27810 56064 27838 56098
rect 27838 56064 27870 56098
rect 27810 56050 27870 56064
rect 28650 56098 28710 56110
rect 28650 56064 28655 56098
rect 28655 56064 28689 56098
rect 28689 56064 28710 56098
rect 28650 56050 28710 56064
rect 28230 55950 28290 56010
rect 28230 55840 28290 55900
rect 27810 55788 27870 55800
rect 27810 55754 27838 55788
rect 27838 55754 27870 55788
rect 27810 55740 27870 55754
rect 28230 55670 28290 55730
rect 28650 55788 28710 55800
rect 28650 55754 28655 55788
rect 28655 55754 28689 55788
rect 28689 55754 28710 55788
rect 28650 55740 28710 55754
rect 27810 54388 27870 54400
rect 28230 54410 28290 54470
rect 27810 54354 27838 54388
rect 27838 54354 27870 54388
rect 27810 54340 27870 54354
rect 28650 54388 28710 54400
rect 28650 54354 28655 54388
rect 28655 54354 28689 54388
rect 28689 54354 28710 54388
rect 28650 54340 28710 54354
rect 28230 54240 28290 54300
rect 28230 54130 28290 54190
rect 27810 54078 27870 54090
rect 27810 54044 27838 54078
rect 27838 54044 27870 54078
rect 27810 54030 27870 54044
rect 28230 53960 28290 54020
rect 28650 54078 28710 54090
rect 28650 54044 28655 54078
rect 28655 54044 28689 54078
rect 28689 54044 28710 54078
rect 28650 54030 28710 54044
rect 27810 52678 27870 52690
rect 28230 52700 28290 52760
rect 27810 52644 27838 52678
rect 27838 52644 27870 52678
rect 27810 52630 27870 52644
rect 28650 52678 28710 52690
rect 28650 52644 28655 52678
rect 28655 52644 28689 52678
rect 28689 52644 28710 52678
rect 28650 52630 28710 52644
rect 28230 52530 28290 52590
rect 28230 52420 28290 52480
rect 27810 52368 27870 52380
rect 27810 52334 27838 52368
rect 27838 52334 27870 52368
rect 27810 52320 27870 52334
rect 28230 52250 28290 52310
rect 28650 52368 28710 52380
rect 28650 52334 28655 52368
rect 28655 52334 28689 52368
rect 28689 52334 28710 52368
rect 28650 52320 28710 52334
rect 27810 50968 27870 50980
rect 28230 50990 28290 51050
rect 27810 50934 27838 50968
rect 27838 50934 27870 50968
rect 27810 50920 27870 50934
rect 28650 50968 28710 50980
rect 28650 50934 28655 50968
rect 28655 50934 28689 50968
rect 28689 50934 28710 50968
rect 28650 50920 28710 50934
rect 28230 50820 28290 50880
rect 28230 50710 28290 50770
rect 27810 50658 27870 50670
rect 27810 50624 27838 50658
rect 27838 50624 27870 50658
rect 27810 50610 27870 50624
rect 28230 50540 28290 50600
rect 28650 50658 28710 50670
rect 28650 50624 28655 50658
rect 28655 50624 28689 50658
rect 28689 50624 28710 50658
rect 28650 50610 28710 50624
rect 27810 49258 27870 49270
rect 28230 49280 28290 49340
rect 27810 49224 27838 49258
rect 27838 49224 27870 49258
rect 27810 49210 27870 49224
rect 28650 49258 28710 49270
rect 28650 49224 28655 49258
rect 28655 49224 28689 49258
rect 28689 49224 28710 49258
rect 28650 49210 28710 49224
rect 28230 49110 28290 49170
rect 28230 49000 28290 49060
rect 27810 48948 27870 48960
rect 27810 48914 27838 48948
rect 27838 48914 27870 48948
rect 27810 48900 27870 48914
rect 28230 48830 28290 48890
rect 28650 48948 28710 48960
rect 28650 48914 28655 48948
rect 28655 48914 28689 48948
rect 28689 48914 28710 48948
rect 28650 48900 28710 48914
rect 27810 47548 27870 47560
rect 28230 47570 28290 47630
rect 27810 47514 27838 47548
rect 27838 47514 27870 47548
rect 27810 47500 27870 47514
rect 28650 47548 28710 47560
rect 28650 47514 28655 47548
rect 28655 47514 28689 47548
rect 28689 47514 28710 47548
rect 28650 47500 28710 47514
rect 28230 47400 28290 47460
rect 28230 47290 28290 47350
rect 27810 47238 27870 47250
rect 27810 47204 27838 47238
rect 27838 47204 27870 47238
rect 27810 47190 27870 47204
rect 28230 47120 28290 47180
rect 28650 47238 28710 47250
rect 28650 47204 28655 47238
rect 28655 47204 28689 47238
rect 28689 47204 28710 47238
rect 28650 47190 28710 47204
rect 27810 45838 27870 45850
rect 28230 45860 28290 45920
rect 27810 45804 27838 45838
rect 27838 45804 27870 45838
rect 27810 45790 27870 45804
rect 28650 45838 28710 45850
rect 28650 45804 28655 45838
rect 28655 45804 28689 45838
rect 28689 45804 28710 45838
rect 28650 45790 28710 45804
rect 28230 45690 28290 45750
rect 28230 45580 28290 45640
rect 27810 45528 27870 45540
rect 27810 45494 27838 45528
rect 27838 45494 27870 45528
rect 27810 45480 27870 45494
rect 28230 45410 28290 45470
rect 28650 45528 28710 45540
rect 28650 45494 28655 45528
rect 28655 45494 28689 45528
rect 28689 45494 28710 45528
rect 28650 45480 28710 45494
rect 27810 44128 27870 44140
rect 28230 44150 28290 44210
rect 27810 44094 27838 44128
rect 27838 44094 27870 44128
rect 27810 44080 27870 44094
rect 28650 44128 28710 44140
rect 28650 44094 28655 44128
rect 28655 44094 28689 44128
rect 28689 44094 28710 44128
rect 28650 44080 28710 44094
rect 28230 43980 28290 44040
rect 28230 43870 28290 43930
rect 27810 43818 27870 43830
rect 27810 43784 27838 43818
rect 27838 43784 27870 43818
rect 27810 43770 27870 43784
rect 28230 43700 28290 43760
rect 28650 43818 28710 43830
rect 28650 43784 28655 43818
rect 28655 43784 28689 43818
rect 28689 43784 28710 43818
rect 28650 43770 28710 43784
rect 27810 42418 27870 42430
rect 28230 42440 28290 42500
rect 27810 42384 27838 42418
rect 27838 42384 27870 42418
rect 27810 42370 27870 42384
rect 28650 42418 28710 42430
rect 28650 42384 28655 42418
rect 28655 42384 28689 42418
rect 28689 42384 28710 42418
rect 28650 42370 28710 42384
rect 28230 42270 28290 42330
rect 28230 42160 28290 42220
rect 27810 42108 27870 42120
rect 27810 42074 27838 42108
rect 27838 42074 27870 42108
rect 27810 42060 27870 42074
rect 28230 41990 28290 42050
rect 28650 42108 28710 42120
rect 28650 42074 28655 42108
rect 28655 42074 28689 42108
rect 28689 42074 28710 42108
rect 28650 42060 28710 42074
rect 27810 40708 27870 40720
rect 28230 40730 28290 40790
rect 27810 40674 27838 40708
rect 27838 40674 27870 40708
rect 27810 40660 27870 40674
rect 28650 40708 28710 40720
rect 28650 40674 28655 40708
rect 28655 40674 28689 40708
rect 28689 40674 28710 40708
rect 28650 40660 28710 40674
rect 28230 40560 28290 40620
rect 28230 40450 28290 40510
rect 27810 40398 27870 40410
rect 27810 40364 27838 40398
rect 27838 40364 27870 40398
rect 27810 40350 27870 40364
rect 28230 40280 28290 40340
rect 28650 40398 28710 40410
rect 28650 40364 28655 40398
rect 28655 40364 28689 40398
rect 28689 40364 28710 40398
rect 28650 40350 28710 40364
rect 27700 39620 27760 39680
rect 28770 39620 28830 39680
rect 28870 66410 28930 66470
rect 28930 65880 28990 65940
rect 28870 64700 28930 64760
rect 28930 64170 28990 64230
rect 28870 62990 28930 63050
rect 28930 62460 28990 62520
rect 28870 61280 28930 61340
rect 28930 60750 28990 60810
rect 28870 59570 28930 59630
rect 28930 59040 28990 59100
rect 28870 57860 28930 57920
rect 28930 57330 28990 57390
rect 28870 56150 28930 56210
rect 28930 55620 28990 55680
rect 28870 54440 28930 54500
rect 28930 53910 28990 53970
rect 28870 52730 28930 52790
rect 28930 52200 28990 52260
rect 28870 51020 28930 51080
rect 28930 50490 28990 50550
rect 28870 49310 28930 49370
rect 28930 48780 28990 48840
rect 28870 47600 28930 47660
rect 28930 47070 28990 47130
rect 28870 45890 28930 45950
rect 28930 45360 28990 45420
rect 28870 44180 28930 44240
rect 28930 43650 28990 43710
rect 28870 42470 28930 42530
rect 28930 41940 28990 42000
rect 28870 40760 28930 40820
rect 27400 39170 27460 39230
rect 28930 40230 28990 40290
rect 28930 39620 28990 39680
rect 29020 66320 29080 66380
rect 29020 64610 29080 64670
rect 29140 62900 29200 62960
rect 29140 61180 29200 61240
rect 29260 59480 29320 59540
rect 29380 57770 29440 57830
rect 29380 56060 29440 56120
rect 29380 54350 29440 54410
rect 29380 52640 29440 52700
rect 29380 50930 29440 50990
rect 29380 49220 29440 49280
rect 29260 47510 29320 47570
rect 29140 45800 29200 45860
rect 29140 44090 29200 44150
rect 29020 42380 29080 42440
rect 29020 40670 29080 40730
rect 32590 66320 32650 66380
rect 32590 64610 32650 64670
rect 32470 62900 32530 62960
rect 32470 61190 32530 61250
rect 32350 59480 32410 59540
rect 32230 57770 32290 57830
rect 32110 56060 32170 56120
rect 31990 54350 32050 54410
rect 31990 52640 32050 52700
rect 32110 50930 32170 50990
rect 31490 39470 31550 39530
rect 32230 49220 32290 49280
rect 29220 39170 29280 39230
rect 29400 39230 29460 39290
rect 29580 39290 29640 39350
rect 29760 39350 29820 39410
rect 31670 39410 31730 39470
rect 32350 47510 32410 47570
rect 31850 39350 31910 39410
rect 32470 45800 32530 45860
rect 32470 44090 32530 44150
rect 32030 39290 32090 39350
rect 32590 42380 32650 42440
rect 32590 40670 32650 40730
rect 32210 39230 32270 39290
rect 32800 66358 32860 66370
rect 33220 66380 33280 66440
rect 32800 66324 32828 66358
rect 32828 66324 32860 66358
rect 32800 66310 32860 66324
rect 33640 66358 33700 66370
rect 33640 66324 33645 66358
rect 33645 66324 33679 66358
rect 33679 66324 33700 66358
rect 33640 66310 33700 66324
rect 33220 66210 33280 66270
rect 33220 66100 33280 66160
rect 32800 66048 32860 66060
rect 32800 66014 32828 66048
rect 32828 66014 32860 66048
rect 32800 66000 32860 66014
rect 33220 65930 33280 65990
rect 33640 66048 33700 66060
rect 33640 66014 33645 66048
rect 33645 66014 33679 66048
rect 33679 66014 33700 66048
rect 33640 66000 33700 66014
rect 32800 64648 32860 64660
rect 33220 64670 33280 64730
rect 32800 64614 32828 64648
rect 32828 64614 32860 64648
rect 32800 64600 32860 64614
rect 33640 64648 33700 64660
rect 33640 64614 33645 64648
rect 33645 64614 33679 64648
rect 33679 64614 33700 64648
rect 33640 64600 33700 64614
rect 33220 64500 33280 64560
rect 33220 64390 33280 64450
rect 32800 64338 32860 64350
rect 32800 64304 32828 64338
rect 32828 64304 32860 64338
rect 32800 64290 32860 64304
rect 33220 64220 33280 64280
rect 33640 64338 33700 64350
rect 33640 64304 33645 64338
rect 33645 64304 33679 64338
rect 33679 64304 33700 64338
rect 33640 64290 33700 64304
rect 32800 62938 32860 62950
rect 33220 62960 33280 63020
rect 32800 62904 32828 62938
rect 32828 62904 32860 62938
rect 32800 62890 32860 62904
rect 33640 62938 33700 62950
rect 33640 62904 33645 62938
rect 33645 62904 33679 62938
rect 33679 62904 33700 62938
rect 33640 62890 33700 62904
rect 33220 62790 33280 62850
rect 33220 62680 33280 62740
rect 32800 62628 32860 62640
rect 32800 62594 32828 62628
rect 32828 62594 32860 62628
rect 32800 62580 32860 62594
rect 33220 62510 33280 62570
rect 33640 62628 33700 62640
rect 33640 62594 33645 62628
rect 33645 62594 33679 62628
rect 33679 62594 33700 62628
rect 33640 62580 33700 62594
rect 32800 61228 32860 61240
rect 33220 61250 33280 61310
rect 32800 61194 32828 61228
rect 32828 61194 32860 61228
rect 32800 61180 32860 61194
rect 33640 61228 33700 61240
rect 33640 61194 33645 61228
rect 33645 61194 33679 61228
rect 33679 61194 33700 61228
rect 33640 61180 33700 61194
rect 33220 61080 33280 61140
rect 33220 60970 33280 61030
rect 32800 60918 32860 60930
rect 32800 60884 32828 60918
rect 32828 60884 32860 60918
rect 32800 60870 32860 60884
rect 33220 60800 33280 60860
rect 33640 60918 33700 60930
rect 33640 60884 33645 60918
rect 33645 60884 33679 60918
rect 33679 60884 33700 60918
rect 33640 60870 33700 60884
rect 32800 59518 32860 59530
rect 33220 59540 33280 59600
rect 32800 59484 32828 59518
rect 32828 59484 32860 59518
rect 32800 59470 32860 59484
rect 33640 59518 33700 59530
rect 33640 59484 33645 59518
rect 33645 59484 33679 59518
rect 33679 59484 33700 59518
rect 33640 59470 33700 59484
rect 33220 59370 33280 59430
rect 33220 59260 33280 59320
rect 32800 59208 32860 59220
rect 32800 59174 32828 59208
rect 32828 59174 32860 59208
rect 32800 59160 32860 59174
rect 33220 59090 33280 59150
rect 33640 59208 33700 59220
rect 33640 59174 33645 59208
rect 33645 59174 33679 59208
rect 33679 59174 33700 59208
rect 33640 59160 33700 59174
rect 32800 57808 32860 57820
rect 33220 57830 33280 57890
rect 32800 57774 32828 57808
rect 32828 57774 32860 57808
rect 32800 57760 32860 57774
rect 33640 57808 33700 57820
rect 33640 57774 33645 57808
rect 33645 57774 33679 57808
rect 33679 57774 33700 57808
rect 33640 57760 33700 57774
rect 33220 57660 33280 57720
rect 33220 57550 33280 57610
rect 32800 57498 32860 57510
rect 32800 57464 32828 57498
rect 32828 57464 32860 57498
rect 32800 57450 32860 57464
rect 33220 57380 33280 57440
rect 33640 57498 33700 57510
rect 33640 57464 33645 57498
rect 33645 57464 33679 57498
rect 33679 57464 33700 57498
rect 33640 57450 33700 57464
rect 32800 56098 32860 56110
rect 33220 56120 33280 56180
rect 32800 56064 32828 56098
rect 32828 56064 32860 56098
rect 32800 56050 32860 56064
rect 33640 56098 33700 56110
rect 33640 56064 33645 56098
rect 33645 56064 33679 56098
rect 33679 56064 33700 56098
rect 33640 56050 33700 56064
rect 33220 55950 33280 56010
rect 33220 55840 33280 55900
rect 32800 55788 32860 55800
rect 32800 55754 32828 55788
rect 32828 55754 32860 55788
rect 32800 55740 32860 55754
rect 33220 55670 33280 55730
rect 33640 55788 33700 55800
rect 33640 55754 33645 55788
rect 33645 55754 33679 55788
rect 33679 55754 33700 55788
rect 33640 55740 33700 55754
rect 32800 54388 32860 54400
rect 33220 54410 33280 54470
rect 32800 54354 32828 54388
rect 32828 54354 32860 54388
rect 32800 54340 32860 54354
rect 33640 54388 33700 54400
rect 33640 54354 33645 54388
rect 33645 54354 33679 54388
rect 33679 54354 33700 54388
rect 33640 54340 33700 54354
rect 33220 54240 33280 54300
rect 33220 54130 33280 54190
rect 32800 54078 32860 54090
rect 32800 54044 32828 54078
rect 32828 54044 32860 54078
rect 32800 54030 32860 54044
rect 33220 53960 33280 54020
rect 33640 54078 33700 54090
rect 33640 54044 33645 54078
rect 33645 54044 33679 54078
rect 33679 54044 33700 54078
rect 33640 54030 33700 54044
rect 32800 52678 32860 52690
rect 33220 52700 33280 52760
rect 32800 52644 32828 52678
rect 32828 52644 32860 52678
rect 32800 52630 32860 52644
rect 33640 52678 33700 52690
rect 33640 52644 33645 52678
rect 33645 52644 33679 52678
rect 33679 52644 33700 52678
rect 33640 52630 33700 52644
rect 33220 52530 33280 52590
rect 33220 52420 33280 52480
rect 32800 52368 32860 52380
rect 32800 52334 32828 52368
rect 32828 52334 32860 52368
rect 32800 52320 32860 52334
rect 33220 52250 33280 52310
rect 33640 52368 33700 52380
rect 33640 52334 33645 52368
rect 33645 52334 33679 52368
rect 33679 52334 33700 52368
rect 33640 52320 33700 52334
rect 32800 50968 32860 50980
rect 33220 50990 33280 51050
rect 32800 50934 32828 50968
rect 32828 50934 32860 50968
rect 32800 50920 32860 50934
rect 33640 50968 33700 50980
rect 33640 50934 33645 50968
rect 33645 50934 33679 50968
rect 33679 50934 33700 50968
rect 33640 50920 33700 50934
rect 33220 50820 33280 50880
rect 33220 50710 33280 50770
rect 32800 50658 32860 50670
rect 32800 50624 32828 50658
rect 32828 50624 32860 50658
rect 32800 50610 32860 50624
rect 33220 50540 33280 50600
rect 33640 50658 33700 50670
rect 33640 50624 33645 50658
rect 33645 50624 33679 50658
rect 33679 50624 33700 50658
rect 33640 50610 33700 50624
rect 32800 49258 32860 49270
rect 33220 49280 33280 49340
rect 32800 49224 32828 49258
rect 32828 49224 32860 49258
rect 32800 49210 32860 49224
rect 33640 49258 33700 49270
rect 33640 49224 33645 49258
rect 33645 49224 33679 49258
rect 33679 49224 33700 49258
rect 33640 49210 33700 49224
rect 33220 49110 33280 49170
rect 33220 49000 33280 49060
rect 32800 48948 32860 48960
rect 32800 48914 32828 48948
rect 32828 48914 32860 48948
rect 32800 48900 32860 48914
rect 33220 48830 33280 48890
rect 33640 48948 33700 48960
rect 33640 48914 33645 48948
rect 33645 48914 33679 48948
rect 33679 48914 33700 48948
rect 33640 48900 33700 48914
rect 32800 47548 32860 47560
rect 33220 47570 33280 47630
rect 32800 47514 32828 47548
rect 32828 47514 32860 47548
rect 32800 47500 32860 47514
rect 33640 47548 33700 47560
rect 33640 47514 33645 47548
rect 33645 47514 33679 47548
rect 33679 47514 33700 47548
rect 33640 47500 33700 47514
rect 33220 47400 33280 47460
rect 33220 47290 33280 47350
rect 32800 47238 32860 47250
rect 32800 47204 32828 47238
rect 32828 47204 32860 47238
rect 32800 47190 32860 47204
rect 33220 47120 33280 47180
rect 33640 47238 33700 47250
rect 33640 47204 33645 47238
rect 33645 47204 33679 47238
rect 33679 47204 33700 47238
rect 33640 47190 33700 47204
rect 32800 45838 32860 45850
rect 33220 45860 33280 45920
rect 32800 45804 32828 45838
rect 32828 45804 32860 45838
rect 32800 45790 32860 45804
rect 33640 45838 33700 45850
rect 33640 45804 33645 45838
rect 33645 45804 33679 45838
rect 33679 45804 33700 45838
rect 33640 45790 33700 45804
rect 33220 45690 33280 45750
rect 33220 45580 33280 45640
rect 32800 45528 32860 45540
rect 32800 45494 32828 45528
rect 32828 45494 32860 45528
rect 32800 45480 32860 45494
rect 33220 45410 33280 45470
rect 33640 45528 33700 45540
rect 33640 45494 33645 45528
rect 33645 45494 33679 45528
rect 33679 45494 33700 45528
rect 33640 45480 33700 45494
rect 32800 44128 32860 44140
rect 33220 44150 33280 44210
rect 32800 44094 32828 44128
rect 32828 44094 32860 44128
rect 32800 44080 32860 44094
rect 33640 44128 33700 44140
rect 33640 44094 33645 44128
rect 33645 44094 33679 44128
rect 33679 44094 33700 44128
rect 33640 44080 33700 44094
rect 33220 43980 33280 44040
rect 33220 43870 33280 43930
rect 32800 43818 32860 43830
rect 32800 43784 32828 43818
rect 32828 43784 32860 43818
rect 32800 43770 32860 43784
rect 33220 43700 33280 43760
rect 33640 43818 33700 43830
rect 33640 43784 33645 43818
rect 33645 43784 33679 43818
rect 33679 43784 33700 43818
rect 33640 43770 33700 43784
rect 32800 42418 32860 42430
rect 33220 42440 33280 42500
rect 32800 42384 32828 42418
rect 32828 42384 32860 42418
rect 32800 42370 32860 42384
rect 33640 42418 33700 42430
rect 33640 42384 33645 42418
rect 33645 42384 33679 42418
rect 33679 42384 33700 42418
rect 33640 42370 33700 42384
rect 33220 42270 33280 42330
rect 33220 42160 33280 42220
rect 32800 42108 32860 42120
rect 32800 42074 32828 42108
rect 32828 42074 32860 42108
rect 32800 42060 32860 42074
rect 33220 41990 33280 42050
rect 33640 42108 33700 42120
rect 33640 42074 33645 42108
rect 33645 42074 33679 42108
rect 33679 42074 33700 42108
rect 33640 42060 33700 42074
rect 32800 40708 32860 40720
rect 33220 40730 33280 40790
rect 32800 40674 32828 40708
rect 32828 40674 32860 40708
rect 32800 40660 32860 40674
rect 33640 40708 33700 40720
rect 33640 40674 33645 40708
rect 33645 40674 33679 40708
rect 33679 40674 33700 40708
rect 33640 40660 33700 40674
rect 33220 40560 33280 40620
rect 33220 40450 33280 40510
rect 32800 40398 32860 40410
rect 32800 40364 32828 40398
rect 32828 40364 32860 40398
rect 32800 40350 32860 40364
rect 33220 40280 33280 40340
rect 33640 40398 33700 40410
rect 33640 40364 33645 40398
rect 33645 40364 33679 40398
rect 33679 40364 33700 40398
rect 33640 40350 33700 40364
rect 32690 39620 32750 39680
rect 33760 39620 33820 39680
rect 33860 66410 33920 66470
rect 33920 65880 33980 65940
rect 33860 64700 33920 64760
rect 33920 64170 33980 64230
rect 33860 62990 33920 63050
rect 33920 62460 33980 62520
rect 33860 61280 33920 61340
rect 33920 60750 33980 60810
rect 33860 59570 33920 59630
rect 33920 59040 33980 59100
rect 33860 57860 33920 57920
rect 33920 57330 33980 57390
rect 33860 56150 33920 56210
rect 33920 55620 33980 55680
rect 33860 54440 33920 54500
rect 33920 53910 33980 53970
rect 33860 52730 33920 52790
rect 33920 52200 33980 52260
rect 33860 51020 33920 51080
rect 33920 50490 33980 50550
rect 33860 49310 33920 49370
rect 33920 48780 33980 48840
rect 33860 47600 33920 47660
rect 33920 47070 33980 47130
rect 33860 45890 33920 45950
rect 33920 45360 33980 45420
rect 33860 44180 33920 44240
rect 33920 43650 33980 43710
rect 33860 42470 33920 42530
rect 33920 41940 33980 42000
rect 33860 40760 33920 40820
rect 32390 39170 32450 39230
rect 33920 40230 33980 40290
rect 33920 39620 33980 39680
rect 34010 66320 34070 66380
rect 34010 64610 34070 64670
rect 34130 62900 34190 62960
rect 34130 61190 34190 61250
rect 34250 59480 34310 59540
rect 34370 57770 34430 57830
rect 34490 56060 34550 56120
rect 34610 54350 34670 54410
rect 34610 52640 34670 52700
rect 34490 50930 34550 50990
rect 34370 49220 34430 49280
rect 34250 47510 34310 47570
rect 34130 45800 34190 45860
rect 34130 44090 34190 44150
rect 34010 42380 34070 42440
rect 34010 40670 34070 40730
rect 36860 54340 36920 54400
rect 37580 66320 37640 66380
rect 37580 64610 37640 64670
rect 37460 62900 37520 62960
rect 37460 61190 37520 61250
rect 37340 59480 37400 59540
rect 37220 57770 37280 57830
rect 37100 56060 37160 56120
rect 36980 52640 37040 52700
rect 34210 39170 34270 39230
rect 34390 39230 34450 39290
rect 34570 39290 34630 39350
rect 34750 39350 34810 39410
rect 34930 39410 34990 39470
rect 35110 39470 35170 39530
rect 36300 39530 36360 39590
rect 37100 50930 37160 50990
rect 36480 39470 36540 39530
rect 37220 49220 37280 49280
rect 36660 39410 36720 39470
rect 37340 47510 37400 47570
rect 36840 39350 36900 39410
rect 37460 45800 37520 45860
rect 37460 44090 37520 44150
rect 37020 39290 37080 39350
rect 37580 42380 37640 42440
rect 37580 40670 37640 40730
rect 37200 39230 37260 39290
rect 37790 66358 37850 66370
rect 38210 66380 38270 66440
rect 37790 66324 37818 66358
rect 37818 66324 37850 66358
rect 37790 66310 37850 66324
rect 38630 66358 38690 66370
rect 38630 66324 38635 66358
rect 38635 66324 38669 66358
rect 38669 66324 38690 66358
rect 38630 66310 38690 66324
rect 38210 66210 38270 66270
rect 38210 66100 38270 66160
rect 37790 66048 37850 66060
rect 37790 66014 37818 66048
rect 37818 66014 37850 66048
rect 37790 66000 37850 66014
rect 38210 65930 38270 65990
rect 38630 66048 38690 66060
rect 38630 66014 38635 66048
rect 38635 66014 38669 66048
rect 38669 66014 38690 66048
rect 38630 66000 38690 66014
rect 37790 64648 37850 64660
rect 38210 64670 38270 64730
rect 37790 64614 37818 64648
rect 37818 64614 37850 64648
rect 37790 64600 37850 64614
rect 38630 64648 38690 64660
rect 38630 64614 38635 64648
rect 38635 64614 38669 64648
rect 38669 64614 38690 64648
rect 38630 64600 38690 64614
rect 38210 64500 38270 64560
rect 38210 64390 38270 64450
rect 37790 64338 37850 64350
rect 37790 64304 37818 64338
rect 37818 64304 37850 64338
rect 37790 64290 37850 64304
rect 38210 64220 38270 64280
rect 38630 64338 38690 64350
rect 38630 64304 38635 64338
rect 38635 64304 38669 64338
rect 38669 64304 38690 64338
rect 38630 64290 38690 64304
rect 37790 62938 37850 62950
rect 38210 62960 38270 63020
rect 37790 62904 37818 62938
rect 37818 62904 37850 62938
rect 37790 62890 37850 62904
rect 38630 62938 38690 62950
rect 38630 62904 38635 62938
rect 38635 62904 38669 62938
rect 38669 62904 38690 62938
rect 38630 62890 38690 62904
rect 38210 62790 38270 62850
rect 38210 62680 38270 62740
rect 37790 62628 37850 62640
rect 37790 62594 37818 62628
rect 37818 62594 37850 62628
rect 37790 62580 37850 62594
rect 38210 62510 38270 62570
rect 38630 62628 38690 62640
rect 38630 62594 38635 62628
rect 38635 62594 38669 62628
rect 38669 62594 38690 62628
rect 38630 62580 38690 62594
rect 37790 61228 37850 61240
rect 38210 61250 38270 61310
rect 37790 61194 37818 61228
rect 37818 61194 37850 61228
rect 37790 61180 37850 61194
rect 38630 61228 38690 61240
rect 38630 61194 38635 61228
rect 38635 61194 38669 61228
rect 38669 61194 38690 61228
rect 38630 61180 38690 61194
rect 38210 61080 38270 61140
rect 38210 60970 38270 61030
rect 37790 60918 37850 60930
rect 37790 60884 37818 60918
rect 37818 60884 37850 60918
rect 37790 60870 37850 60884
rect 38210 60800 38270 60860
rect 38630 60918 38690 60930
rect 38630 60884 38635 60918
rect 38635 60884 38669 60918
rect 38669 60884 38690 60918
rect 38630 60870 38690 60884
rect 37790 59518 37850 59530
rect 38210 59540 38270 59600
rect 37790 59484 37818 59518
rect 37818 59484 37850 59518
rect 37790 59470 37850 59484
rect 38630 59518 38690 59530
rect 38630 59484 38635 59518
rect 38635 59484 38669 59518
rect 38669 59484 38690 59518
rect 38630 59470 38690 59484
rect 38210 59370 38270 59430
rect 38210 59260 38270 59320
rect 37790 59208 37850 59220
rect 37790 59174 37818 59208
rect 37818 59174 37850 59208
rect 37790 59160 37850 59174
rect 38210 59090 38270 59150
rect 38630 59208 38690 59220
rect 38630 59174 38635 59208
rect 38635 59174 38669 59208
rect 38669 59174 38690 59208
rect 38630 59160 38690 59174
rect 37790 57808 37850 57820
rect 38210 57830 38270 57890
rect 37790 57774 37818 57808
rect 37818 57774 37850 57808
rect 37790 57760 37850 57774
rect 38630 57808 38690 57820
rect 38630 57774 38635 57808
rect 38635 57774 38669 57808
rect 38669 57774 38690 57808
rect 38630 57760 38690 57774
rect 38210 57660 38270 57720
rect 38210 57550 38270 57610
rect 37790 57498 37850 57510
rect 37790 57464 37818 57498
rect 37818 57464 37850 57498
rect 37790 57450 37850 57464
rect 38210 57380 38270 57440
rect 38630 57498 38690 57510
rect 38630 57464 38635 57498
rect 38635 57464 38669 57498
rect 38669 57464 38690 57498
rect 38630 57450 38690 57464
rect 37790 56098 37850 56110
rect 38210 56120 38270 56180
rect 37790 56064 37818 56098
rect 37818 56064 37850 56098
rect 37790 56050 37850 56064
rect 38630 56098 38690 56110
rect 38630 56064 38635 56098
rect 38635 56064 38669 56098
rect 38669 56064 38690 56098
rect 38630 56050 38690 56064
rect 38210 55950 38270 56010
rect 38210 55840 38270 55900
rect 37790 55788 37850 55800
rect 37790 55754 37818 55788
rect 37818 55754 37850 55788
rect 37790 55740 37850 55754
rect 38210 55670 38270 55730
rect 38630 55788 38690 55800
rect 38630 55754 38635 55788
rect 38635 55754 38669 55788
rect 38669 55754 38690 55788
rect 38630 55740 38690 55754
rect 37790 54388 37850 54400
rect 38210 54410 38270 54470
rect 37790 54354 37818 54388
rect 37818 54354 37850 54388
rect 37790 54340 37850 54354
rect 38630 54388 38690 54400
rect 38630 54354 38635 54388
rect 38635 54354 38669 54388
rect 38669 54354 38690 54388
rect 38630 54340 38690 54354
rect 38210 54240 38270 54300
rect 38210 54130 38270 54190
rect 37790 54078 37850 54090
rect 37790 54044 37818 54078
rect 37818 54044 37850 54078
rect 37790 54030 37850 54044
rect 38210 53960 38270 54020
rect 38630 54078 38690 54090
rect 38630 54044 38635 54078
rect 38635 54044 38669 54078
rect 38669 54044 38690 54078
rect 38630 54030 38690 54044
rect 37790 52678 37850 52690
rect 38210 52700 38270 52760
rect 37790 52644 37818 52678
rect 37818 52644 37850 52678
rect 37790 52630 37850 52644
rect 38630 52678 38690 52690
rect 38630 52644 38635 52678
rect 38635 52644 38669 52678
rect 38669 52644 38690 52678
rect 38630 52630 38690 52644
rect 38210 52530 38270 52590
rect 38210 52420 38270 52480
rect 37790 52368 37850 52380
rect 37790 52334 37818 52368
rect 37818 52334 37850 52368
rect 37790 52320 37850 52334
rect 38210 52250 38270 52310
rect 38630 52368 38690 52380
rect 38630 52334 38635 52368
rect 38635 52334 38669 52368
rect 38669 52334 38690 52368
rect 38630 52320 38690 52334
rect 37790 50968 37850 50980
rect 38210 50990 38270 51050
rect 37790 50934 37818 50968
rect 37818 50934 37850 50968
rect 37790 50920 37850 50934
rect 38630 50968 38690 50980
rect 38630 50934 38635 50968
rect 38635 50934 38669 50968
rect 38669 50934 38690 50968
rect 38630 50920 38690 50934
rect 38210 50820 38270 50880
rect 38210 50710 38270 50770
rect 37790 50658 37850 50670
rect 37790 50624 37818 50658
rect 37818 50624 37850 50658
rect 37790 50610 37850 50624
rect 38210 50540 38270 50600
rect 38630 50658 38690 50670
rect 38630 50624 38635 50658
rect 38635 50624 38669 50658
rect 38669 50624 38690 50658
rect 38630 50610 38690 50624
rect 37790 49258 37850 49270
rect 38210 49280 38270 49340
rect 37790 49224 37818 49258
rect 37818 49224 37850 49258
rect 37790 49210 37850 49224
rect 38630 49258 38690 49270
rect 38630 49224 38635 49258
rect 38635 49224 38669 49258
rect 38669 49224 38690 49258
rect 38630 49210 38690 49224
rect 38210 49110 38270 49170
rect 38210 49000 38270 49060
rect 37790 48948 37850 48960
rect 37790 48914 37818 48948
rect 37818 48914 37850 48948
rect 37790 48900 37850 48914
rect 38210 48830 38270 48890
rect 38630 48948 38690 48960
rect 38630 48914 38635 48948
rect 38635 48914 38669 48948
rect 38669 48914 38690 48948
rect 38630 48900 38690 48914
rect 37790 47548 37850 47560
rect 38210 47570 38270 47630
rect 37790 47514 37818 47548
rect 37818 47514 37850 47548
rect 37790 47500 37850 47514
rect 38630 47548 38690 47560
rect 38630 47514 38635 47548
rect 38635 47514 38669 47548
rect 38669 47514 38690 47548
rect 38630 47500 38690 47514
rect 38210 47400 38270 47460
rect 38210 47290 38270 47350
rect 37790 47238 37850 47250
rect 37790 47204 37818 47238
rect 37818 47204 37850 47238
rect 37790 47190 37850 47204
rect 38210 47120 38270 47180
rect 38630 47238 38690 47250
rect 38630 47204 38635 47238
rect 38635 47204 38669 47238
rect 38669 47204 38690 47238
rect 38630 47190 38690 47204
rect 37790 45838 37850 45850
rect 38210 45860 38270 45920
rect 37790 45804 37818 45838
rect 37818 45804 37850 45838
rect 37790 45790 37850 45804
rect 38630 45838 38690 45850
rect 38630 45804 38635 45838
rect 38635 45804 38669 45838
rect 38669 45804 38690 45838
rect 38630 45790 38690 45804
rect 38210 45690 38270 45750
rect 38210 45580 38270 45640
rect 37790 45528 37850 45540
rect 37790 45494 37818 45528
rect 37818 45494 37850 45528
rect 37790 45480 37850 45494
rect 38210 45410 38270 45470
rect 38630 45528 38690 45540
rect 38630 45494 38635 45528
rect 38635 45494 38669 45528
rect 38669 45494 38690 45528
rect 38630 45480 38690 45494
rect 37790 44128 37850 44140
rect 38210 44150 38270 44210
rect 37790 44094 37818 44128
rect 37818 44094 37850 44128
rect 37790 44080 37850 44094
rect 38630 44128 38690 44140
rect 38630 44094 38635 44128
rect 38635 44094 38669 44128
rect 38669 44094 38690 44128
rect 38630 44080 38690 44094
rect 38210 43980 38270 44040
rect 38210 43870 38270 43930
rect 37790 43818 37850 43830
rect 37790 43784 37818 43818
rect 37818 43784 37850 43818
rect 37790 43770 37850 43784
rect 38210 43700 38270 43760
rect 38630 43818 38690 43830
rect 38630 43784 38635 43818
rect 38635 43784 38669 43818
rect 38669 43784 38690 43818
rect 38630 43770 38690 43784
rect 37790 42418 37850 42430
rect 38210 42440 38270 42500
rect 37790 42384 37818 42418
rect 37818 42384 37850 42418
rect 37790 42370 37850 42384
rect 38630 42418 38690 42430
rect 38630 42384 38635 42418
rect 38635 42384 38669 42418
rect 38669 42384 38690 42418
rect 38630 42370 38690 42384
rect 38210 42270 38270 42330
rect 38210 42160 38270 42220
rect 37790 42108 37850 42120
rect 37790 42074 37818 42108
rect 37818 42074 37850 42108
rect 37790 42060 37850 42074
rect 38210 41990 38270 42050
rect 38630 42108 38690 42120
rect 38630 42074 38635 42108
rect 38635 42074 38669 42108
rect 38669 42074 38690 42108
rect 38630 42060 38690 42074
rect 37790 40708 37850 40720
rect 38210 40730 38270 40790
rect 37790 40674 37818 40708
rect 37818 40674 37850 40708
rect 37790 40660 37850 40674
rect 38630 40708 38690 40720
rect 38630 40674 38635 40708
rect 38635 40674 38669 40708
rect 38669 40674 38690 40708
rect 38630 40660 38690 40674
rect 38210 40560 38270 40620
rect 38210 40450 38270 40510
rect 37790 40398 37850 40410
rect 37790 40364 37818 40398
rect 37818 40364 37850 40398
rect 37790 40350 37850 40364
rect 38210 40280 38270 40340
rect 38630 40398 38690 40410
rect 38630 40364 38635 40398
rect 38635 40364 38669 40398
rect 38669 40364 38690 40398
rect 38630 40350 38690 40364
rect 37680 39620 37740 39680
rect 38750 39620 38810 39680
rect 38850 66410 38910 66470
rect 38910 65880 38970 65940
rect 38850 64700 38910 64760
rect 38910 64170 38970 64230
rect 38850 62990 38910 63050
rect 38910 62460 38970 62520
rect 38850 61280 38910 61340
rect 38910 60750 38970 60810
rect 38850 59570 38910 59630
rect 38910 59040 38970 59100
rect 38850 57860 38910 57920
rect 38910 57330 38970 57390
rect 38850 56150 38910 56210
rect 38910 55620 38970 55680
rect 38850 54440 38910 54500
rect 38910 53910 38970 53970
rect 38850 52730 38910 52790
rect 38910 52200 38970 52260
rect 38850 51020 38910 51080
rect 38910 50490 38970 50550
rect 38850 49310 38910 49370
rect 38910 48780 38970 48840
rect 38850 47600 38910 47660
rect 38910 47070 38970 47130
rect 38850 45890 38910 45950
rect 38910 45360 38970 45420
rect 38850 44180 38910 44240
rect 38910 43650 38970 43710
rect 38850 42470 38910 42530
rect 38910 41940 38970 42000
rect 38850 40760 38910 40820
rect 37380 39170 37440 39230
rect 38910 40230 38970 40290
rect 38910 39620 38970 39680
rect 39000 66320 39060 66380
rect 39000 64610 39060 64670
rect 39120 62900 39180 62960
rect 39120 61190 39180 61250
rect 39240 59480 39300 59540
rect 39360 57770 39420 57830
rect 39480 56060 39540 56120
rect 39720 54340 39780 54400
rect 41850 54340 41910 54400
rect 39600 52640 39660 52700
rect 39480 50930 39540 50990
rect 39360 49220 39420 49280
rect 39240 47510 39300 47570
rect 39120 45800 39180 45860
rect 39120 44080 39180 44140
rect 39000 42370 39060 42430
rect 39000 40670 39060 40730
rect 42570 66320 42630 66380
rect 42570 64610 42630 64670
rect 42450 62900 42510 62960
rect 42450 61190 42510 61250
rect 42330 59480 42390 59540
rect 42210 57770 42270 57830
rect 42090 56060 42150 56120
rect 41970 52640 42030 52700
rect 39200 39170 39260 39230
rect 39380 39230 39440 39290
rect 39560 39290 39620 39350
rect 39740 39350 39800 39410
rect 39920 39410 39980 39470
rect 40100 39470 40160 39530
rect 40280 39530 40340 39590
rect 41290 39530 41350 39590
rect 42090 50930 42150 50990
rect 41470 39470 41530 39530
rect 42210 49220 42270 49280
rect 41650 39410 41710 39470
rect 42330 47510 42390 47570
rect 41830 39350 41890 39410
rect 42450 45800 42510 45860
rect 42450 44090 42510 44150
rect 42010 39290 42070 39350
rect 42570 42380 42630 42440
rect 42570 40670 42630 40730
rect 42190 39230 42250 39290
rect 42780 66358 42840 66370
rect 43200 66380 43260 66440
rect 42780 66324 42808 66358
rect 42808 66324 42840 66358
rect 42780 66310 42840 66324
rect 43620 66358 43680 66370
rect 43620 66324 43625 66358
rect 43625 66324 43659 66358
rect 43659 66324 43680 66358
rect 43620 66310 43680 66324
rect 43200 66210 43260 66270
rect 43200 66100 43260 66160
rect 42780 66048 42840 66060
rect 42780 66014 42808 66048
rect 42808 66014 42840 66048
rect 42780 66000 42840 66014
rect 43200 65930 43260 65990
rect 43620 66048 43680 66060
rect 43620 66014 43625 66048
rect 43625 66014 43659 66048
rect 43659 66014 43680 66048
rect 43620 66000 43680 66014
rect 42780 64648 42840 64660
rect 43200 64670 43260 64730
rect 42780 64614 42808 64648
rect 42808 64614 42840 64648
rect 42780 64600 42840 64614
rect 43620 64648 43680 64660
rect 43620 64614 43625 64648
rect 43625 64614 43659 64648
rect 43659 64614 43680 64648
rect 43620 64600 43680 64614
rect 43200 64500 43260 64560
rect 43200 64390 43260 64450
rect 42780 64338 42840 64350
rect 42780 64304 42808 64338
rect 42808 64304 42840 64338
rect 42780 64290 42840 64304
rect 43200 64220 43260 64280
rect 43620 64338 43680 64350
rect 43620 64304 43625 64338
rect 43625 64304 43659 64338
rect 43659 64304 43680 64338
rect 43620 64290 43680 64304
rect 42780 62938 42840 62950
rect 43200 62960 43260 63020
rect 42780 62904 42808 62938
rect 42808 62904 42840 62938
rect 42780 62890 42840 62904
rect 43620 62938 43680 62950
rect 43620 62904 43625 62938
rect 43625 62904 43659 62938
rect 43659 62904 43680 62938
rect 43620 62890 43680 62904
rect 43200 62790 43260 62850
rect 43200 62680 43260 62740
rect 42780 62628 42840 62640
rect 42780 62594 42808 62628
rect 42808 62594 42840 62628
rect 42780 62580 42840 62594
rect 43200 62510 43260 62570
rect 43620 62628 43680 62640
rect 43620 62594 43625 62628
rect 43625 62594 43659 62628
rect 43659 62594 43680 62628
rect 43620 62580 43680 62594
rect 42780 61228 42840 61240
rect 43200 61250 43260 61310
rect 42780 61194 42808 61228
rect 42808 61194 42840 61228
rect 42780 61180 42840 61194
rect 43620 61228 43680 61240
rect 43620 61194 43625 61228
rect 43625 61194 43659 61228
rect 43659 61194 43680 61228
rect 43620 61180 43680 61194
rect 43200 61080 43260 61140
rect 43200 60970 43260 61030
rect 42780 60918 42840 60930
rect 42780 60884 42808 60918
rect 42808 60884 42840 60918
rect 42780 60870 42840 60884
rect 43200 60800 43260 60860
rect 43620 60918 43680 60930
rect 43620 60884 43625 60918
rect 43625 60884 43659 60918
rect 43659 60884 43680 60918
rect 43620 60870 43680 60884
rect 42780 59518 42840 59530
rect 43200 59540 43260 59600
rect 42780 59484 42808 59518
rect 42808 59484 42840 59518
rect 42780 59470 42840 59484
rect 43620 59518 43680 59530
rect 43620 59484 43625 59518
rect 43625 59484 43659 59518
rect 43659 59484 43680 59518
rect 43620 59470 43680 59484
rect 43200 59370 43260 59430
rect 43200 59260 43260 59320
rect 42780 59208 42840 59220
rect 42780 59174 42808 59208
rect 42808 59174 42840 59208
rect 42780 59160 42840 59174
rect 43200 59090 43260 59150
rect 43620 59208 43680 59220
rect 43620 59174 43625 59208
rect 43625 59174 43659 59208
rect 43659 59174 43680 59208
rect 43620 59160 43680 59174
rect 42780 57808 42840 57820
rect 43200 57830 43260 57890
rect 42780 57774 42808 57808
rect 42808 57774 42840 57808
rect 42780 57760 42840 57774
rect 43620 57808 43680 57820
rect 43620 57774 43625 57808
rect 43625 57774 43659 57808
rect 43659 57774 43680 57808
rect 43620 57760 43680 57774
rect 43200 57660 43260 57720
rect 43200 57550 43260 57610
rect 42780 57498 42840 57510
rect 42780 57464 42808 57498
rect 42808 57464 42840 57498
rect 42780 57450 42840 57464
rect 43200 57380 43260 57440
rect 43620 57498 43680 57510
rect 43620 57464 43625 57498
rect 43625 57464 43659 57498
rect 43659 57464 43680 57498
rect 43620 57450 43680 57464
rect 42780 56098 42840 56110
rect 43200 56120 43260 56180
rect 42780 56064 42808 56098
rect 42808 56064 42840 56098
rect 42780 56050 42840 56064
rect 43620 56098 43680 56110
rect 43620 56064 43625 56098
rect 43625 56064 43659 56098
rect 43659 56064 43680 56098
rect 43620 56050 43680 56064
rect 43200 55950 43260 56010
rect 43200 55840 43260 55900
rect 42780 55788 42840 55800
rect 42780 55754 42808 55788
rect 42808 55754 42840 55788
rect 42780 55740 42840 55754
rect 43200 55670 43260 55730
rect 43620 55788 43680 55800
rect 43620 55754 43625 55788
rect 43625 55754 43659 55788
rect 43659 55754 43680 55788
rect 43620 55740 43680 55754
rect 42780 54388 42840 54400
rect 43200 54410 43260 54470
rect 42780 54354 42808 54388
rect 42808 54354 42840 54388
rect 42780 54340 42840 54354
rect 43620 54388 43680 54400
rect 43620 54354 43625 54388
rect 43625 54354 43659 54388
rect 43659 54354 43680 54388
rect 43620 54340 43680 54354
rect 43200 54240 43260 54300
rect 43200 54130 43260 54190
rect 42780 54078 42840 54090
rect 42780 54044 42808 54078
rect 42808 54044 42840 54078
rect 42780 54030 42840 54044
rect 43200 53960 43260 54020
rect 43620 54078 43680 54090
rect 43620 54044 43625 54078
rect 43625 54044 43659 54078
rect 43659 54044 43680 54078
rect 43620 54030 43680 54044
rect 42780 52678 42840 52690
rect 43200 52700 43260 52760
rect 42780 52644 42808 52678
rect 42808 52644 42840 52678
rect 42780 52630 42840 52644
rect 43620 52678 43680 52690
rect 43620 52644 43625 52678
rect 43625 52644 43659 52678
rect 43659 52644 43680 52678
rect 43620 52630 43680 52644
rect 43200 52530 43260 52590
rect 43200 52420 43260 52480
rect 42780 52368 42840 52380
rect 42780 52334 42808 52368
rect 42808 52334 42840 52368
rect 42780 52320 42840 52334
rect 43200 52250 43260 52310
rect 43620 52368 43680 52380
rect 43620 52334 43625 52368
rect 43625 52334 43659 52368
rect 43659 52334 43680 52368
rect 43620 52320 43680 52334
rect 42780 50968 42840 50980
rect 43200 50990 43260 51050
rect 42780 50934 42808 50968
rect 42808 50934 42840 50968
rect 42780 50920 42840 50934
rect 43620 50968 43680 50980
rect 43620 50934 43625 50968
rect 43625 50934 43659 50968
rect 43659 50934 43680 50968
rect 43620 50920 43680 50934
rect 43200 50820 43260 50880
rect 43200 50710 43260 50770
rect 42780 50658 42840 50670
rect 42780 50624 42808 50658
rect 42808 50624 42840 50658
rect 42780 50610 42840 50624
rect 43200 50540 43260 50600
rect 43620 50658 43680 50670
rect 43620 50624 43625 50658
rect 43625 50624 43659 50658
rect 43659 50624 43680 50658
rect 43620 50610 43680 50624
rect 42780 49258 42840 49270
rect 43200 49280 43260 49340
rect 42780 49224 42808 49258
rect 42808 49224 42840 49258
rect 42780 49210 42840 49224
rect 43620 49258 43680 49270
rect 43620 49224 43625 49258
rect 43625 49224 43659 49258
rect 43659 49224 43680 49258
rect 43620 49210 43680 49224
rect 43200 49110 43260 49170
rect 43200 49000 43260 49060
rect 42780 48948 42840 48960
rect 42780 48914 42808 48948
rect 42808 48914 42840 48948
rect 42780 48900 42840 48914
rect 43200 48830 43260 48890
rect 43620 48948 43680 48960
rect 43620 48914 43625 48948
rect 43625 48914 43659 48948
rect 43659 48914 43680 48948
rect 43620 48900 43680 48914
rect 42780 47548 42840 47560
rect 43200 47570 43260 47630
rect 42780 47514 42808 47548
rect 42808 47514 42840 47548
rect 42780 47500 42840 47514
rect 43620 47548 43680 47560
rect 43620 47514 43625 47548
rect 43625 47514 43659 47548
rect 43659 47514 43680 47548
rect 43620 47500 43680 47514
rect 43200 47400 43260 47460
rect 43200 47290 43260 47350
rect 42780 47238 42840 47250
rect 42780 47204 42808 47238
rect 42808 47204 42840 47238
rect 42780 47190 42840 47204
rect 43200 47120 43260 47180
rect 43620 47238 43680 47250
rect 43620 47204 43625 47238
rect 43625 47204 43659 47238
rect 43659 47204 43680 47238
rect 43620 47190 43680 47204
rect 42780 45838 42840 45850
rect 43200 45860 43260 45920
rect 42780 45804 42808 45838
rect 42808 45804 42840 45838
rect 42780 45790 42840 45804
rect 43620 45838 43680 45850
rect 43620 45804 43625 45838
rect 43625 45804 43659 45838
rect 43659 45804 43680 45838
rect 43620 45790 43680 45804
rect 43200 45690 43260 45750
rect 43200 45580 43260 45640
rect 42780 45528 42840 45540
rect 42780 45494 42808 45528
rect 42808 45494 42840 45528
rect 42780 45480 42840 45494
rect 43200 45410 43260 45470
rect 43620 45528 43680 45540
rect 43620 45494 43625 45528
rect 43625 45494 43659 45528
rect 43659 45494 43680 45528
rect 43620 45480 43680 45494
rect 42780 44128 42840 44140
rect 43200 44150 43260 44210
rect 42780 44094 42808 44128
rect 42808 44094 42840 44128
rect 42780 44080 42840 44094
rect 43620 44128 43680 44140
rect 43620 44094 43625 44128
rect 43625 44094 43659 44128
rect 43659 44094 43680 44128
rect 43620 44080 43680 44094
rect 43200 43980 43260 44040
rect 43200 43870 43260 43930
rect 42780 43818 42840 43830
rect 42780 43784 42808 43818
rect 42808 43784 42840 43818
rect 42780 43770 42840 43784
rect 43200 43700 43260 43760
rect 43620 43818 43680 43830
rect 43620 43784 43625 43818
rect 43625 43784 43659 43818
rect 43659 43784 43680 43818
rect 43620 43770 43680 43784
rect 42780 42418 42840 42430
rect 43200 42440 43260 42500
rect 42780 42384 42808 42418
rect 42808 42384 42840 42418
rect 42780 42370 42840 42384
rect 43620 42418 43680 42430
rect 43620 42384 43625 42418
rect 43625 42384 43659 42418
rect 43659 42384 43680 42418
rect 43620 42370 43680 42384
rect 43200 42270 43260 42330
rect 43200 42160 43260 42220
rect 42780 42108 42840 42120
rect 42780 42074 42808 42108
rect 42808 42074 42840 42108
rect 42780 42060 42840 42074
rect 43200 41990 43260 42050
rect 43620 42108 43680 42120
rect 43620 42074 43625 42108
rect 43625 42074 43659 42108
rect 43659 42074 43680 42108
rect 43620 42060 43680 42074
rect 42780 40708 42840 40720
rect 43200 40730 43260 40790
rect 42780 40674 42808 40708
rect 42808 40674 42840 40708
rect 42780 40660 42840 40674
rect 43620 40708 43680 40720
rect 43620 40674 43625 40708
rect 43625 40674 43659 40708
rect 43659 40674 43680 40708
rect 43620 40660 43680 40674
rect 43200 40560 43260 40620
rect 43200 40450 43260 40510
rect 42780 40398 42840 40410
rect 42780 40364 42808 40398
rect 42808 40364 42840 40398
rect 42780 40350 42840 40364
rect 43200 40280 43260 40340
rect 43620 40398 43680 40410
rect 43620 40364 43625 40398
rect 43625 40364 43659 40398
rect 43659 40364 43680 40398
rect 43620 40350 43680 40364
rect 42670 39620 42730 39680
rect 43740 39620 43800 39680
rect 43840 66410 43900 66470
rect 43900 65880 43960 65940
rect 43840 64700 43900 64760
rect 43900 64170 43960 64230
rect 43840 62990 43900 63050
rect 43900 62460 43960 62520
rect 43840 61280 43900 61340
rect 43900 60750 43960 60810
rect 43840 59570 43900 59630
rect 43900 59040 43960 59100
rect 43840 57860 43900 57920
rect 43900 57330 43960 57390
rect 43840 56150 43900 56210
rect 43900 55620 43960 55680
rect 43840 54440 43900 54500
rect 43900 53910 43960 53970
rect 43840 52730 43900 52790
rect 43900 52200 43960 52260
rect 43840 51020 43900 51080
rect 43900 50490 43960 50550
rect 43840 49310 43900 49370
rect 43900 48780 43960 48840
rect 43840 47600 43900 47660
rect 43900 47070 43960 47130
rect 43840 45890 43900 45950
rect 43900 45360 43960 45420
rect 43840 44180 43900 44240
rect 43900 43650 43960 43710
rect 43840 42470 43900 42530
rect 43900 41940 43960 42000
rect 43840 40760 43900 40820
rect 42370 39170 42430 39230
rect 43900 40230 43960 40290
rect 43900 39620 43960 39680
rect 43990 66320 44050 66380
rect 43990 64610 44050 64670
rect 44110 62900 44170 62960
rect 44110 61190 44170 61250
rect 44230 59480 44290 59540
rect 44350 57770 44410 57830
rect 44470 56060 44530 56120
rect 44710 54340 44770 54400
rect 44590 52640 44650 52700
rect 44470 50930 44530 50990
rect 44350 49220 44410 49280
rect 44230 47510 44290 47570
rect 44110 45800 44170 45860
rect 44110 44080 44170 44140
rect 43990 42370 44050 42430
rect 43990 40670 44050 40730
rect 47560 66320 47620 66380
rect 47560 64610 47620 64670
rect 47440 62900 47500 62960
rect 47440 61190 47500 61250
rect 47320 59480 47380 59540
rect 47200 57770 47260 57830
rect 47080 56060 47140 56120
rect 46960 54350 47020 54410
rect 46960 52640 47020 52700
rect 44190 39170 44250 39230
rect 44370 39230 44430 39290
rect 44550 39290 44610 39350
rect 44730 39350 44790 39410
rect 44910 39410 44970 39470
rect 45090 39470 45150 39530
rect 45270 39530 45330 39590
rect 47080 50930 47140 50990
rect 46460 39470 46520 39530
rect 47200 49220 47260 49280
rect 46640 39410 46700 39470
rect 47320 47510 47380 47570
rect 46820 39350 46880 39410
rect 47440 45800 47500 45860
rect 47440 44090 47500 44150
rect 47000 39290 47060 39350
rect 47560 42380 47620 42440
rect 47560 40670 47620 40730
rect 47180 39230 47240 39290
rect 47770 66358 47830 66370
rect 48190 66380 48250 66440
rect 47770 66324 47798 66358
rect 47798 66324 47830 66358
rect 47770 66310 47830 66324
rect 48610 66358 48670 66370
rect 48610 66324 48615 66358
rect 48615 66324 48649 66358
rect 48649 66324 48670 66358
rect 48610 66310 48670 66324
rect 48190 66210 48250 66270
rect 48190 66100 48250 66160
rect 47770 66048 47830 66060
rect 47770 66014 47798 66048
rect 47798 66014 47830 66048
rect 47770 66000 47830 66014
rect 48190 65930 48250 65990
rect 48610 66048 48670 66060
rect 48610 66014 48615 66048
rect 48615 66014 48649 66048
rect 48649 66014 48670 66048
rect 48610 66000 48670 66014
rect 47770 64648 47830 64660
rect 48190 64670 48250 64730
rect 47770 64614 47798 64648
rect 47798 64614 47830 64648
rect 47770 64600 47830 64614
rect 48610 64648 48670 64660
rect 48610 64614 48615 64648
rect 48615 64614 48649 64648
rect 48649 64614 48670 64648
rect 48610 64600 48670 64614
rect 48190 64500 48250 64560
rect 48190 64390 48250 64450
rect 47770 64338 47830 64350
rect 47770 64304 47798 64338
rect 47798 64304 47830 64338
rect 47770 64290 47830 64304
rect 48190 64220 48250 64280
rect 48610 64338 48670 64350
rect 48610 64304 48615 64338
rect 48615 64304 48649 64338
rect 48649 64304 48670 64338
rect 48610 64290 48670 64304
rect 47770 62938 47830 62950
rect 48190 62960 48250 63020
rect 47770 62904 47798 62938
rect 47798 62904 47830 62938
rect 47770 62890 47830 62904
rect 48610 62938 48670 62950
rect 48610 62904 48615 62938
rect 48615 62904 48649 62938
rect 48649 62904 48670 62938
rect 48610 62890 48670 62904
rect 48190 62790 48250 62850
rect 48190 62680 48250 62740
rect 47770 62628 47830 62640
rect 47770 62594 47798 62628
rect 47798 62594 47830 62628
rect 47770 62580 47830 62594
rect 48190 62510 48250 62570
rect 48610 62628 48670 62640
rect 48610 62594 48615 62628
rect 48615 62594 48649 62628
rect 48649 62594 48670 62628
rect 48610 62580 48670 62594
rect 47770 61228 47830 61240
rect 48190 61250 48250 61310
rect 47770 61194 47798 61228
rect 47798 61194 47830 61228
rect 47770 61180 47830 61194
rect 48610 61228 48670 61240
rect 48610 61194 48615 61228
rect 48615 61194 48649 61228
rect 48649 61194 48670 61228
rect 48610 61180 48670 61194
rect 48190 61080 48250 61140
rect 48190 60970 48250 61030
rect 47770 60918 47830 60930
rect 47770 60884 47798 60918
rect 47798 60884 47830 60918
rect 47770 60870 47830 60884
rect 48190 60800 48250 60860
rect 48610 60918 48670 60930
rect 48610 60884 48615 60918
rect 48615 60884 48649 60918
rect 48649 60884 48670 60918
rect 48610 60870 48670 60884
rect 47770 59518 47830 59530
rect 48190 59540 48250 59600
rect 47770 59484 47798 59518
rect 47798 59484 47830 59518
rect 47770 59470 47830 59484
rect 48610 59518 48670 59530
rect 48610 59484 48615 59518
rect 48615 59484 48649 59518
rect 48649 59484 48670 59518
rect 48610 59470 48670 59484
rect 48190 59370 48250 59430
rect 48190 59260 48250 59320
rect 47770 59208 47830 59220
rect 47770 59174 47798 59208
rect 47798 59174 47830 59208
rect 47770 59160 47830 59174
rect 48190 59090 48250 59150
rect 48610 59208 48670 59220
rect 48610 59174 48615 59208
rect 48615 59174 48649 59208
rect 48649 59174 48670 59208
rect 48610 59160 48670 59174
rect 47770 57808 47830 57820
rect 48190 57830 48250 57890
rect 47770 57774 47798 57808
rect 47798 57774 47830 57808
rect 47770 57760 47830 57774
rect 48610 57808 48670 57820
rect 48610 57774 48615 57808
rect 48615 57774 48649 57808
rect 48649 57774 48670 57808
rect 48610 57760 48670 57774
rect 48190 57660 48250 57720
rect 48190 57550 48250 57610
rect 47770 57498 47830 57510
rect 47770 57464 47798 57498
rect 47798 57464 47830 57498
rect 47770 57450 47830 57464
rect 48190 57380 48250 57440
rect 48610 57498 48670 57510
rect 48610 57464 48615 57498
rect 48615 57464 48649 57498
rect 48649 57464 48670 57498
rect 48610 57450 48670 57464
rect 47770 56098 47830 56110
rect 48190 56120 48250 56180
rect 47770 56064 47798 56098
rect 47798 56064 47830 56098
rect 47770 56050 47830 56064
rect 48610 56098 48670 56110
rect 48610 56064 48615 56098
rect 48615 56064 48649 56098
rect 48649 56064 48670 56098
rect 48610 56050 48670 56064
rect 48190 55950 48250 56010
rect 48190 55840 48250 55900
rect 47770 55788 47830 55800
rect 47770 55754 47798 55788
rect 47798 55754 47830 55788
rect 47770 55740 47830 55754
rect 48190 55670 48250 55730
rect 48610 55788 48670 55800
rect 48610 55754 48615 55788
rect 48615 55754 48649 55788
rect 48649 55754 48670 55788
rect 48610 55740 48670 55754
rect 47770 54388 47830 54400
rect 48190 54410 48250 54470
rect 47770 54354 47798 54388
rect 47798 54354 47830 54388
rect 47770 54340 47830 54354
rect 48610 54388 48670 54400
rect 48610 54354 48615 54388
rect 48615 54354 48649 54388
rect 48649 54354 48670 54388
rect 48610 54340 48670 54354
rect 48190 54240 48250 54300
rect 48190 54130 48250 54190
rect 47770 54078 47830 54090
rect 47770 54044 47798 54078
rect 47798 54044 47830 54078
rect 47770 54030 47830 54044
rect 48190 53960 48250 54020
rect 48610 54078 48670 54090
rect 48610 54044 48615 54078
rect 48615 54044 48649 54078
rect 48649 54044 48670 54078
rect 48610 54030 48670 54044
rect 47770 52678 47830 52690
rect 48190 52700 48250 52760
rect 47770 52644 47798 52678
rect 47798 52644 47830 52678
rect 47770 52630 47830 52644
rect 48610 52678 48670 52690
rect 48610 52644 48615 52678
rect 48615 52644 48649 52678
rect 48649 52644 48670 52678
rect 48610 52630 48670 52644
rect 48190 52530 48250 52590
rect 48190 52420 48250 52480
rect 47770 52368 47830 52380
rect 47770 52334 47798 52368
rect 47798 52334 47830 52368
rect 47770 52320 47830 52334
rect 48190 52250 48250 52310
rect 48610 52368 48670 52380
rect 48610 52334 48615 52368
rect 48615 52334 48649 52368
rect 48649 52334 48670 52368
rect 48610 52320 48670 52334
rect 47770 50968 47830 50980
rect 48190 50990 48250 51050
rect 47770 50934 47798 50968
rect 47798 50934 47830 50968
rect 47770 50920 47830 50934
rect 48610 50968 48670 50980
rect 48610 50934 48615 50968
rect 48615 50934 48649 50968
rect 48649 50934 48670 50968
rect 48610 50920 48670 50934
rect 48190 50820 48250 50880
rect 48190 50710 48250 50770
rect 47770 50658 47830 50670
rect 47770 50624 47798 50658
rect 47798 50624 47830 50658
rect 47770 50610 47830 50624
rect 48190 50540 48250 50600
rect 48610 50658 48670 50670
rect 48610 50624 48615 50658
rect 48615 50624 48649 50658
rect 48649 50624 48670 50658
rect 48610 50610 48670 50624
rect 47770 49258 47830 49270
rect 48190 49280 48250 49340
rect 47770 49224 47798 49258
rect 47798 49224 47830 49258
rect 47770 49210 47830 49224
rect 48610 49258 48670 49270
rect 48610 49224 48615 49258
rect 48615 49224 48649 49258
rect 48649 49224 48670 49258
rect 48610 49210 48670 49224
rect 48190 49110 48250 49170
rect 48190 49000 48250 49060
rect 47770 48948 47830 48960
rect 47770 48914 47798 48948
rect 47798 48914 47830 48948
rect 47770 48900 47830 48914
rect 48190 48830 48250 48890
rect 48610 48948 48670 48960
rect 48610 48914 48615 48948
rect 48615 48914 48649 48948
rect 48649 48914 48670 48948
rect 48610 48900 48670 48914
rect 47770 47548 47830 47560
rect 48190 47570 48250 47630
rect 47770 47514 47798 47548
rect 47798 47514 47830 47548
rect 47770 47500 47830 47514
rect 48610 47548 48670 47560
rect 48610 47514 48615 47548
rect 48615 47514 48649 47548
rect 48649 47514 48670 47548
rect 48610 47500 48670 47514
rect 48190 47400 48250 47460
rect 48190 47290 48250 47350
rect 47770 47238 47830 47250
rect 47770 47204 47798 47238
rect 47798 47204 47830 47238
rect 47770 47190 47830 47204
rect 48190 47120 48250 47180
rect 48610 47238 48670 47250
rect 48610 47204 48615 47238
rect 48615 47204 48649 47238
rect 48649 47204 48670 47238
rect 48610 47190 48670 47204
rect 47770 45838 47830 45850
rect 48190 45860 48250 45920
rect 47770 45804 47798 45838
rect 47798 45804 47830 45838
rect 47770 45790 47830 45804
rect 48610 45838 48670 45850
rect 48610 45804 48615 45838
rect 48615 45804 48649 45838
rect 48649 45804 48670 45838
rect 48610 45790 48670 45804
rect 48190 45690 48250 45750
rect 48190 45580 48250 45640
rect 47770 45528 47830 45540
rect 47770 45494 47798 45528
rect 47798 45494 47830 45528
rect 47770 45480 47830 45494
rect 48190 45410 48250 45470
rect 48610 45528 48670 45540
rect 48610 45494 48615 45528
rect 48615 45494 48649 45528
rect 48649 45494 48670 45528
rect 48610 45480 48670 45494
rect 47770 44128 47830 44140
rect 48190 44150 48250 44210
rect 47770 44094 47798 44128
rect 47798 44094 47830 44128
rect 47770 44080 47830 44094
rect 48610 44128 48670 44140
rect 48610 44094 48615 44128
rect 48615 44094 48649 44128
rect 48649 44094 48670 44128
rect 48610 44080 48670 44094
rect 48190 43980 48250 44040
rect 48190 43870 48250 43930
rect 47770 43818 47830 43830
rect 47770 43784 47798 43818
rect 47798 43784 47830 43818
rect 47770 43770 47830 43784
rect 48190 43700 48250 43760
rect 48610 43818 48670 43830
rect 48610 43784 48615 43818
rect 48615 43784 48649 43818
rect 48649 43784 48670 43818
rect 48610 43770 48670 43784
rect 47770 42418 47830 42430
rect 48190 42440 48250 42500
rect 47770 42384 47798 42418
rect 47798 42384 47830 42418
rect 47770 42370 47830 42384
rect 48610 42418 48670 42430
rect 48610 42384 48615 42418
rect 48615 42384 48649 42418
rect 48649 42384 48670 42418
rect 48610 42370 48670 42384
rect 48190 42270 48250 42330
rect 48190 42160 48250 42220
rect 47770 42108 47830 42120
rect 47770 42074 47798 42108
rect 47798 42074 47830 42108
rect 47770 42060 47830 42074
rect 48190 41990 48250 42050
rect 48610 42108 48670 42120
rect 48610 42074 48615 42108
rect 48615 42074 48649 42108
rect 48649 42074 48670 42108
rect 48610 42060 48670 42074
rect 47770 40708 47830 40720
rect 48190 40730 48250 40790
rect 47770 40674 47798 40708
rect 47798 40674 47830 40708
rect 47770 40660 47830 40674
rect 48610 40708 48670 40720
rect 48610 40674 48615 40708
rect 48615 40674 48649 40708
rect 48649 40674 48670 40708
rect 48610 40660 48670 40674
rect 48190 40560 48250 40620
rect 48190 40450 48250 40510
rect 47770 40398 47830 40410
rect 47770 40364 47798 40398
rect 47798 40364 47830 40398
rect 47770 40350 47830 40364
rect 48190 40280 48250 40340
rect 48610 40398 48670 40410
rect 48610 40364 48615 40398
rect 48615 40364 48649 40398
rect 48649 40364 48670 40398
rect 48610 40350 48670 40364
rect 47660 39620 47720 39680
rect 48730 39620 48790 39680
rect 48830 66410 48890 66470
rect 48890 65880 48950 65940
rect 48830 64700 48890 64760
rect 48890 64170 48950 64230
rect 48830 62990 48890 63050
rect 48890 62460 48950 62520
rect 48830 61280 48890 61340
rect 48890 60750 48950 60810
rect 48830 59570 48890 59630
rect 48890 59040 48950 59100
rect 48830 57860 48890 57920
rect 48890 57330 48950 57390
rect 48830 56150 48890 56210
rect 48890 55620 48950 55680
rect 48830 54440 48890 54500
rect 48890 53910 48950 53970
rect 48830 52730 48890 52790
rect 48890 52200 48950 52260
rect 48830 51020 48890 51080
rect 48890 50490 48950 50550
rect 48830 49310 48890 49370
rect 48890 48780 48950 48840
rect 48830 47600 48890 47660
rect 48890 47070 48950 47130
rect 48830 45890 48890 45950
rect 48890 45360 48950 45420
rect 48830 44180 48890 44240
rect 48890 43650 48950 43710
rect 48830 42470 48890 42530
rect 48890 41940 48950 42000
rect 48830 40760 48890 40820
rect 47360 39170 47420 39230
rect 48890 40230 48950 40290
rect 48890 39620 48950 39680
rect 48980 66320 49040 66380
rect 48980 64610 49040 64670
rect 49100 62900 49160 62960
rect 49100 61190 49160 61250
rect 49220 59480 49280 59540
rect 49340 57770 49400 57830
rect 49460 56060 49520 56120
rect 49580 54350 49640 54410
rect 49580 52640 49640 52700
rect 49460 50930 49520 50990
rect 49340 49220 49400 49280
rect 49220 47510 49280 47570
rect 49100 45800 49160 45860
rect 49100 44090 49160 44150
rect 48980 42380 49040 42440
rect 48980 40670 49040 40730
rect 52550 66320 52610 66380
rect 52550 64610 52610 64670
rect 52430 62900 52490 62960
rect 52430 61180 52490 61240
rect 52310 59480 52370 59540
rect 52190 57770 52250 57830
rect 52190 56060 52250 56120
rect 52190 54350 52250 54410
rect 52190 52640 52250 52700
rect 52190 50930 52250 50990
rect 52190 49220 52250 49280
rect 49180 39170 49240 39230
rect 49360 39230 49420 39290
rect 49540 39290 49600 39350
rect 49720 39350 49780 39410
rect 49900 39410 49960 39470
rect 50080 39470 50140 39530
rect 52310 47510 52370 47570
rect 51810 39350 51870 39410
rect 52430 45800 52490 45860
rect 52430 44090 52490 44150
rect 51990 39290 52050 39350
rect 52550 42380 52610 42440
rect 52550 40670 52610 40730
rect 52170 39230 52230 39290
rect 52760 66358 52820 66370
rect 53180 66380 53240 66440
rect 52760 66324 52788 66358
rect 52788 66324 52820 66358
rect 52760 66310 52820 66324
rect 53600 66358 53660 66370
rect 53600 66324 53605 66358
rect 53605 66324 53639 66358
rect 53639 66324 53660 66358
rect 53600 66310 53660 66324
rect 53180 66210 53240 66270
rect 53180 66100 53240 66160
rect 52760 66048 52820 66060
rect 52760 66014 52788 66048
rect 52788 66014 52820 66048
rect 52760 66000 52820 66014
rect 53180 65930 53240 65990
rect 53600 66048 53660 66060
rect 53600 66014 53605 66048
rect 53605 66014 53639 66048
rect 53639 66014 53660 66048
rect 53600 66000 53660 66014
rect 52760 64648 52820 64660
rect 53180 64670 53240 64730
rect 52760 64614 52788 64648
rect 52788 64614 52820 64648
rect 52760 64600 52820 64614
rect 53600 64648 53660 64660
rect 53600 64614 53605 64648
rect 53605 64614 53639 64648
rect 53639 64614 53660 64648
rect 53600 64600 53660 64614
rect 53180 64500 53240 64560
rect 53180 64390 53240 64450
rect 52760 64338 52820 64350
rect 52760 64304 52788 64338
rect 52788 64304 52820 64338
rect 52760 64290 52820 64304
rect 53180 64220 53240 64280
rect 53600 64338 53660 64350
rect 53600 64304 53605 64338
rect 53605 64304 53639 64338
rect 53639 64304 53660 64338
rect 53600 64290 53660 64304
rect 52760 62938 52820 62950
rect 53180 62960 53240 63020
rect 52760 62904 52788 62938
rect 52788 62904 52820 62938
rect 52760 62890 52820 62904
rect 53600 62938 53660 62950
rect 53600 62904 53605 62938
rect 53605 62904 53639 62938
rect 53639 62904 53660 62938
rect 53600 62890 53660 62904
rect 53180 62790 53240 62850
rect 53180 62680 53240 62740
rect 52760 62628 52820 62640
rect 52760 62594 52788 62628
rect 52788 62594 52820 62628
rect 52760 62580 52820 62594
rect 53180 62510 53240 62570
rect 53600 62628 53660 62640
rect 53600 62594 53605 62628
rect 53605 62594 53639 62628
rect 53639 62594 53660 62628
rect 53600 62580 53660 62594
rect 52760 61228 52820 61240
rect 53180 61250 53240 61310
rect 52760 61194 52788 61228
rect 52788 61194 52820 61228
rect 52760 61180 52820 61194
rect 53600 61228 53660 61240
rect 53600 61194 53605 61228
rect 53605 61194 53639 61228
rect 53639 61194 53660 61228
rect 53600 61180 53660 61194
rect 53180 61080 53240 61140
rect 53180 60970 53240 61030
rect 52760 60918 52820 60930
rect 52760 60884 52788 60918
rect 52788 60884 52820 60918
rect 52760 60870 52820 60884
rect 53180 60800 53240 60860
rect 53600 60918 53660 60930
rect 53600 60884 53605 60918
rect 53605 60884 53639 60918
rect 53639 60884 53660 60918
rect 53600 60870 53660 60884
rect 52760 59518 52820 59530
rect 53180 59540 53240 59600
rect 52760 59484 52788 59518
rect 52788 59484 52820 59518
rect 52760 59470 52820 59484
rect 53600 59518 53660 59530
rect 53600 59484 53605 59518
rect 53605 59484 53639 59518
rect 53639 59484 53660 59518
rect 53600 59470 53660 59484
rect 53180 59370 53240 59430
rect 53180 59260 53240 59320
rect 52760 59208 52820 59220
rect 52760 59174 52788 59208
rect 52788 59174 52820 59208
rect 52760 59160 52820 59174
rect 53180 59090 53240 59150
rect 53600 59208 53660 59220
rect 53600 59174 53605 59208
rect 53605 59174 53639 59208
rect 53639 59174 53660 59208
rect 53600 59160 53660 59174
rect 52760 57808 52820 57820
rect 53180 57830 53240 57890
rect 52760 57774 52788 57808
rect 52788 57774 52820 57808
rect 52760 57760 52820 57774
rect 53600 57808 53660 57820
rect 53600 57774 53605 57808
rect 53605 57774 53639 57808
rect 53639 57774 53660 57808
rect 53600 57760 53660 57774
rect 53180 57660 53240 57720
rect 53180 57550 53240 57610
rect 52760 57498 52820 57510
rect 52760 57464 52788 57498
rect 52788 57464 52820 57498
rect 52760 57450 52820 57464
rect 53180 57380 53240 57440
rect 53600 57498 53660 57510
rect 53600 57464 53605 57498
rect 53605 57464 53639 57498
rect 53639 57464 53660 57498
rect 53600 57450 53660 57464
rect 52760 56098 52820 56110
rect 53180 56120 53240 56180
rect 52760 56064 52788 56098
rect 52788 56064 52820 56098
rect 52760 56050 52820 56064
rect 53600 56098 53660 56110
rect 53600 56064 53605 56098
rect 53605 56064 53639 56098
rect 53639 56064 53660 56098
rect 53600 56050 53660 56064
rect 53180 55950 53240 56010
rect 53180 55840 53240 55900
rect 52760 55788 52820 55800
rect 52760 55754 52788 55788
rect 52788 55754 52820 55788
rect 52760 55740 52820 55754
rect 53180 55670 53240 55730
rect 53600 55788 53660 55800
rect 53600 55754 53605 55788
rect 53605 55754 53639 55788
rect 53639 55754 53660 55788
rect 53600 55740 53660 55754
rect 52760 54388 52820 54400
rect 53180 54410 53240 54470
rect 52760 54354 52788 54388
rect 52788 54354 52820 54388
rect 52760 54340 52820 54354
rect 53600 54388 53660 54400
rect 53600 54354 53605 54388
rect 53605 54354 53639 54388
rect 53639 54354 53660 54388
rect 53600 54340 53660 54354
rect 53180 54240 53240 54300
rect 53180 54130 53240 54190
rect 52760 54078 52820 54090
rect 52760 54044 52788 54078
rect 52788 54044 52820 54078
rect 52760 54030 52820 54044
rect 53180 53960 53240 54020
rect 53600 54078 53660 54090
rect 53600 54044 53605 54078
rect 53605 54044 53639 54078
rect 53639 54044 53660 54078
rect 53600 54030 53660 54044
rect 52760 52678 52820 52690
rect 53180 52700 53240 52760
rect 52760 52644 52788 52678
rect 52788 52644 52820 52678
rect 52760 52630 52820 52644
rect 53600 52678 53660 52690
rect 53600 52644 53605 52678
rect 53605 52644 53639 52678
rect 53639 52644 53660 52678
rect 53600 52630 53660 52644
rect 53180 52530 53240 52590
rect 53180 52420 53240 52480
rect 52760 52368 52820 52380
rect 52760 52334 52788 52368
rect 52788 52334 52820 52368
rect 52760 52320 52820 52334
rect 53180 52250 53240 52310
rect 53600 52368 53660 52380
rect 53600 52334 53605 52368
rect 53605 52334 53639 52368
rect 53639 52334 53660 52368
rect 53600 52320 53660 52334
rect 52760 50968 52820 50980
rect 53180 50990 53240 51050
rect 52760 50934 52788 50968
rect 52788 50934 52820 50968
rect 52760 50920 52820 50934
rect 53600 50968 53660 50980
rect 53600 50934 53605 50968
rect 53605 50934 53639 50968
rect 53639 50934 53660 50968
rect 53600 50920 53660 50934
rect 53180 50820 53240 50880
rect 53180 50710 53240 50770
rect 52760 50658 52820 50670
rect 52760 50624 52788 50658
rect 52788 50624 52820 50658
rect 52760 50610 52820 50624
rect 53180 50540 53240 50600
rect 53600 50658 53660 50670
rect 53600 50624 53605 50658
rect 53605 50624 53639 50658
rect 53639 50624 53660 50658
rect 53600 50610 53660 50624
rect 52760 49258 52820 49270
rect 53180 49280 53240 49340
rect 52760 49224 52788 49258
rect 52788 49224 52820 49258
rect 52760 49210 52820 49224
rect 53600 49258 53660 49270
rect 53600 49224 53605 49258
rect 53605 49224 53639 49258
rect 53639 49224 53660 49258
rect 53600 49210 53660 49224
rect 53180 49110 53240 49170
rect 53180 49000 53240 49060
rect 52760 48948 52820 48960
rect 52760 48914 52788 48948
rect 52788 48914 52820 48948
rect 52760 48900 52820 48914
rect 53180 48830 53240 48890
rect 53600 48948 53660 48960
rect 53600 48914 53605 48948
rect 53605 48914 53639 48948
rect 53639 48914 53660 48948
rect 53600 48900 53660 48914
rect 52760 47548 52820 47560
rect 53180 47570 53240 47630
rect 52760 47514 52788 47548
rect 52788 47514 52820 47548
rect 52760 47500 52820 47514
rect 53600 47548 53660 47560
rect 53600 47514 53605 47548
rect 53605 47514 53639 47548
rect 53639 47514 53660 47548
rect 53600 47500 53660 47514
rect 53180 47400 53240 47460
rect 53180 47290 53240 47350
rect 52760 47238 52820 47250
rect 52760 47204 52788 47238
rect 52788 47204 52820 47238
rect 52760 47190 52820 47204
rect 53180 47120 53240 47180
rect 53600 47238 53660 47250
rect 53600 47204 53605 47238
rect 53605 47204 53639 47238
rect 53639 47204 53660 47238
rect 53600 47190 53660 47204
rect 52760 45838 52820 45850
rect 53180 45860 53240 45920
rect 52760 45804 52788 45838
rect 52788 45804 52820 45838
rect 52760 45790 52820 45804
rect 53600 45838 53660 45850
rect 53600 45804 53605 45838
rect 53605 45804 53639 45838
rect 53639 45804 53660 45838
rect 53600 45790 53660 45804
rect 53180 45690 53240 45750
rect 53180 45580 53240 45640
rect 52760 45528 52820 45540
rect 52760 45494 52788 45528
rect 52788 45494 52820 45528
rect 52760 45480 52820 45494
rect 53180 45410 53240 45470
rect 53600 45528 53660 45540
rect 53600 45494 53605 45528
rect 53605 45494 53639 45528
rect 53639 45494 53660 45528
rect 53600 45480 53660 45494
rect 52760 44128 52820 44140
rect 53180 44150 53240 44210
rect 52760 44094 52788 44128
rect 52788 44094 52820 44128
rect 52760 44080 52820 44094
rect 53600 44128 53660 44140
rect 53600 44094 53605 44128
rect 53605 44094 53639 44128
rect 53639 44094 53660 44128
rect 53600 44080 53660 44094
rect 53180 43980 53240 44040
rect 53180 43870 53240 43930
rect 52760 43818 52820 43830
rect 52760 43784 52788 43818
rect 52788 43784 52820 43818
rect 52760 43770 52820 43784
rect 53180 43700 53240 43760
rect 53600 43818 53660 43830
rect 53600 43784 53605 43818
rect 53605 43784 53639 43818
rect 53639 43784 53660 43818
rect 53600 43770 53660 43784
rect 52760 42418 52820 42430
rect 53180 42440 53240 42500
rect 52760 42384 52788 42418
rect 52788 42384 52820 42418
rect 52760 42370 52820 42384
rect 53600 42418 53660 42430
rect 53600 42384 53605 42418
rect 53605 42384 53639 42418
rect 53639 42384 53660 42418
rect 53600 42370 53660 42384
rect 53180 42270 53240 42330
rect 53180 42160 53240 42220
rect 52760 42108 52820 42120
rect 52760 42074 52788 42108
rect 52788 42074 52820 42108
rect 52760 42060 52820 42074
rect 53180 41990 53240 42050
rect 53600 42108 53660 42120
rect 53600 42074 53605 42108
rect 53605 42074 53639 42108
rect 53639 42074 53660 42108
rect 53600 42060 53660 42074
rect 52760 40708 52820 40720
rect 53180 40730 53240 40790
rect 52760 40674 52788 40708
rect 52788 40674 52820 40708
rect 52760 40660 52820 40674
rect 53600 40708 53660 40720
rect 53600 40674 53605 40708
rect 53605 40674 53639 40708
rect 53639 40674 53660 40708
rect 53600 40660 53660 40674
rect 53180 40560 53240 40620
rect 53180 40450 53240 40510
rect 52760 40398 52820 40410
rect 52760 40364 52788 40398
rect 52788 40364 52820 40398
rect 52760 40350 52820 40364
rect 53180 40280 53240 40340
rect 53600 40398 53660 40410
rect 53600 40364 53605 40398
rect 53605 40364 53639 40398
rect 53639 40364 53660 40398
rect 53600 40350 53660 40364
rect 52650 39620 52710 39680
rect 53720 39620 53780 39680
rect 53820 66410 53880 66470
rect 53880 65880 53940 65940
rect 53820 64700 53880 64760
rect 53880 64170 53940 64230
rect 53820 62990 53880 63050
rect 53880 62460 53940 62520
rect 53820 61280 53880 61340
rect 53880 60750 53940 60810
rect 53820 59570 53880 59630
rect 53880 59040 53940 59100
rect 53820 57860 53880 57920
rect 53880 57330 53940 57390
rect 53820 56150 53880 56210
rect 53880 55620 53940 55680
rect 53820 54440 53880 54500
rect 53880 53910 53940 53970
rect 53820 52730 53880 52790
rect 53880 52200 53940 52260
rect 53820 51020 53880 51080
rect 53880 50490 53940 50550
rect 53820 49310 53880 49370
rect 53880 48780 53940 48840
rect 53820 47600 53880 47660
rect 53880 47070 53940 47130
rect 53820 45890 53880 45950
rect 53880 45360 53940 45420
rect 53820 44180 53880 44240
rect 53880 43650 53940 43710
rect 53820 42470 53880 42530
rect 53880 41940 53940 42000
rect 53820 40760 53880 40820
rect 52350 39170 52410 39230
rect 53880 40230 53940 40290
rect 53880 39620 53940 39680
rect 53970 66320 54030 66380
rect 53970 64610 54030 64670
rect 54090 62900 54150 62960
rect 54090 61180 54150 61240
rect 54210 59480 54270 59540
rect 54330 57770 54390 57830
rect 54330 56060 54390 56120
rect 54330 54350 54390 54410
rect 54330 52640 54390 52700
rect 54330 50930 54390 50990
rect 54330 49220 54390 49280
rect 54210 47510 54270 47570
rect 54090 45800 54150 45860
rect 54090 44090 54150 44150
rect 53970 42380 54030 42440
rect 53970 40670 54030 40730
rect 57540 66320 57600 66380
rect 57540 64610 57600 64670
rect 57420 62900 57480 62960
rect 57420 61180 57480 61240
rect 57300 59480 57360 59540
rect 57180 57770 57240 57830
rect 57180 56060 57240 56120
rect 57180 54350 57240 54410
rect 57180 52640 57240 52700
rect 57180 50930 57240 50990
rect 57180 49220 57240 49280
rect 57300 47510 57360 47570
rect 54170 39170 54230 39230
rect 54350 39230 54410 39290
rect 54530 39290 54590 39350
rect 54710 39350 54770 39410
rect 56800 39350 56860 39410
rect 57420 45800 57480 45860
rect 57420 44090 57480 44150
rect 56980 39290 57040 39350
rect 57540 42380 57600 42440
rect 57540 40670 57600 40730
rect 57160 39230 57220 39290
rect 57750 66358 57810 66370
rect 58170 66380 58230 66440
rect 57750 66324 57778 66358
rect 57778 66324 57810 66358
rect 57750 66310 57810 66324
rect 58590 66358 58650 66370
rect 58590 66324 58595 66358
rect 58595 66324 58629 66358
rect 58629 66324 58650 66358
rect 58590 66310 58650 66324
rect 58170 66210 58230 66270
rect 58170 66100 58230 66160
rect 57750 66048 57810 66060
rect 57750 66014 57778 66048
rect 57778 66014 57810 66048
rect 57750 66000 57810 66014
rect 58170 65930 58230 65990
rect 58590 66048 58650 66060
rect 58590 66014 58595 66048
rect 58595 66014 58629 66048
rect 58629 66014 58650 66048
rect 58590 66000 58650 66014
rect 57750 64648 57810 64660
rect 58170 64670 58230 64730
rect 57750 64614 57778 64648
rect 57778 64614 57810 64648
rect 57750 64600 57810 64614
rect 58590 64648 58650 64660
rect 58590 64614 58595 64648
rect 58595 64614 58629 64648
rect 58629 64614 58650 64648
rect 58590 64600 58650 64614
rect 58170 64500 58230 64560
rect 58170 64390 58230 64450
rect 57750 64338 57810 64350
rect 57750 64304 57778 64338
rect 57778 64304 57810 64338
rect 57750 64290 57810 64304
rect 58170 64220 58230 64280
rect 58590 64338 58650 64350
rect 58590 64304 58595 64338
rect 58595 64304 58629 64338
rect 58629 64304 58650 64338
rect 58590 64290 58650 64304
rect 57750 62938 57810 62950
rect 58170 62960 58230 63020
rect 57750 62904 57778 62938
rect 57778 62904 57810 62938
rect 57750 62890 57810 62904
rect 58590 62938 58650 62950
rect 58590 62904 58595 62938
rect 58595 62904 58629 62938
rect 58629 62904 58650 62938
rect 58590 62890 58650 62904
rect 58170 62790 58230 62850
rect 58170 62680 58230 62740
rect 57750 62628 57810 62640
rect 57750 62594 57778 62628
rect 57778 62594 57810 62628
rect 57750 62580 57810 62594
rect 58170 62510 58230 62570
rect 58590 62628 58650 62640
rect 58590 62594 58595 62628
rect 58595 62594 58629 62628
rect 58629 62594 58650 62628
rect 58590 62580 58650 62594
rect 57750 61228 57810 61240
rect 58170 61250 58230 61310
rect 57750 61194 57778 61228
rect 57778 61194 57810 61228
rect 57750 61180 57810 61194
rect 58590 61228 58650 61240
rect 58590 61194 58595 61228
rect 58595 61194 58629 61228
rect 58629 61194 58650 61228
rect 58590 61180 58650 61194
rect 58170 61080 58230 61140
rect 58170 60970 58230 61030
rect 57750 60918 57810 60930
rect 57750 60884 57778 60918
rect 57778 60884 57810 60918
rect 57750 60870 57810 60884
rect 58170 60800 58230 60860
rect 58590 60918 58650 60930
rect 58590 60884 58595 60918
rect 58595 60884 58629 60918
rect 58629 60884 58650 60918
rect 58590 60870 58650 60884
rect 57750 59518 57810 59530
rect 58170 59540 58230 59600
rect 57750 59484 57778 59518
rect 57778 59484 57810 59518
rect 57750 59470 57810 59484
rect 58590 59518 58650 59530
rect 58590 59484 58595 59518
rect 58595 59484 58629 59518
rect 58629 59484 58650 59518
rect 58590 59470 58650 59484
rect 58170 59370 58230 59430
rect 58170 59260 58230 59320
rect 57750 59208 57810 59220
rect 57750 59174 57778 59208
rect 57778 59174 57810 59208
rect 57750 59160 57810 59174
rect 58170 59090 58230 59150
rect 58590 59208 58650 59220
rect 58590 59174 58595 59208
rect 58595 59174 58629 59208
rect 58629 59174 58650 59208
rect 58590 59160 58650 59174
rect 57750 57808 57810 57820
rect 58170 57830 58230 57890
rect 57750 57774 57778 57808
rect 57778 57774 57810 57808
rect 57750 57760 57810 57774
rect 58590 57808 58650 57820
rect 58590 57774 58595 57808
rect 58595 57774 58629 57808
rect 58629 57774 58650 57808
rect 58590 57760 58650 57774
rect 58170 57660 58230 57720
rect 58170 57550 58230 57610
rect 57750 57498 57810 57510
rect 57750 57464 57778 57498
rect 57778 57464 57810 57498
rect 57750 57450 57810 57464
rect 58170 57380 58230 57440
rect 58590 57498 58650 57510
rect 58590 57464 58595 57498
rect 58595 57464 58629 57498
rect 58629 57464 58650 57498
rect 58590 57450 58650 57464
rect 57750 56098 57810 56110
rect 58170 56120 58230 56180
rect 57750 56064 57778 56098
rect 57778 56064 57810 56098
rect 57750 56050 57810 56064
rect 58590 56098 58650 56110
rect 58590 56064 58595 56098
rect 58595 56064 58629 56098
rect 58629 56064 58650 56098
rect 58590 56050 58650 56064
rect 58170 55950 58230 56010
rect 58170 55840 58230 55900
rect 57750 55788 57810 55800
rect 57750 55754 57778 55788
rect 57778 55754 57810 55788
rect 57750 55740 57810 55754
rect 58170 55670 58230 55730
rect 58590 55788 58650 55800
rect 58590 55754 58595 55788
rect 58595 55754 58629 55788
rect 58629 55754 58650 55788
rect 58590 55740 58650 55754
rect 57750 54388 57810 54400
rect 58170 54410 58230 54470
rect 57750 54354 57778 54388
rect 57778 54354 57810 54388
rect 57750 54340 57810 54354
rect 58590 54388 58650 54400
rect 58590 54354 58595 54388
rect 58595 54354 58629 54388
rect 58629 54354 58650 54388
rect 58590 54340 58650 54354
rect 58170 54240 58230 54300
rect 58170 54130 58230 54190
rect 57750 54078 57810 54090
rect 57750 54044 57778 54078
rect 57778 54044 57810 54078
rect 57750 54030 57810 54044
rect 58170 53960 58230 54020
rect 58590 54078 58650 54090
rect 58590 54044 58595 54078
rect 58595 54044 58629 54078
rect 58629 54044 58650 54078
rect 58590 54030 58650 54044
rect 57750 52678 57810 52690
rect 58170 52700 58230 52760
rect 57750 52644 57778 52678
rect 57778 52644 57810 52678
rect 57750 52630 57810 52644
rect 58590 52678 58650 52690
rect 58590 52644 58595 52678
rect 58595 52644 58629 52678
rect 58629 52644 58650 52678
rect 58590 52630 58650 52644
rect 58170 52530 58230 52590
rect 58170 52420 58230 52480
rect 57750 52368 57810 52380
rect 57750 52334 57778 52368
rect 57778 52334 57810 52368
rect 57750 52320 57810 52334
rect 58170 52250 58230 52310
rect 58590 52368 58650 52380
rect 58590 52334 58595 52368
rect 58595 52334 58629 52368
rect 58629 52334 58650 52368
rect 58590 52320 58650 52334
rect 57750 50968 57810 50980
rect 58170 50990 58230 51050
rect 57750 50934 57778 50968
rect 57778 50934 57810 50968
rect 57750 50920 57810 50934
rect 58590 50968 58650 50980
rect 58590 50934 58595 50968
rect 58595 50934 58629 50968
rect 58629 50934 58650 50968
rect 58590 50920 58650 50934
rect 58170 50820 58230 50880
rect 58170 50710 58230 50770
rect 57750 50658 57810 50670
rect 57750 50624 57778 50658
rect 57778 50624 57810 50658
rect 57750 50610 57810 50624
rect 58170 50540 58230 50600
rect 58590 50658 58650 50670
rect 58590 50624 58595 50658
rect 58595 50624 58629 50658
rect 58629 50624 58650 50658
rect 58590 50610 58650 50624
rect 57750 49258 57810 49270
rect 58170 49280 58230 49340
rect 57750 49224 57778 49258
rect 57778 49224 57810 49258
rect 57750 49210 57810 49224
rect 58590 49258 58650 49270
rect 58590 49224 58595 49258
rect 58595 49224 58629 49258
rect 58629 49224 58650 49258
rect 58590 49210 58650 49224
rect 58170 49110 58230 49170
rect 58170 49000 58230 49060
rect 57750 48948 57810 48960
rect 57750 48914 57778 48948
rect 57778 48914 57810 48948
rect 57750 48900 57810 48914
rect 58170 48830 58230 48890
rect 58590 48948 58650 48960
rect 58590 48914 58595 48948
rect 58595 48914 58629 48948
rect 58629 48914 58650 48948
rect 58590 48900 58650 48914
rect 57750 47548 57810 47560
rect 58170 47570 58230 47630
rect 57750 47514 57778 47548
rect 57778 47514 57810 47548
rect 57750 47500 57810 47514
rect 58590 47548 58650 47560
rect 58590 47514 58595 47548
rect 58595 47514 58629 47548
rect 58629 47514 58650 47548
rect 58590 47500 58650 47514
rect 58170 47400 58230 47460
rect 58170 47290 58230 47350
rect 57750 47238 57810 47250
rect 57750 47204 57778 47238
rect 57778 47204 57810 47238
rect 57750 47190 57810 47204
rect 58170 47120 58230 47180
rect 58590 47238 58650 47250
rect 58590 47204 58595 47238
rect 58595 47204 58629 47238
rect 58629 47204 58650 47238
rect 58590 47190 58650 47204
rect 57750 45838 57810 45850
rect 58170 45860 58230 45920
rect 57750 45804 57778 45838
rect 57778 45804 57810 45838
rect 57750 45790 57810 45804
rect 58590 45838 58650 45850
rect 58590 45804 58595 45838
rect 58595 45804 58629 45838
rect 58629 45804 58650 45838
rect 58590 45790 58650 45804
rect 58170 45690 58230 45750
rect 58170 45580 58230 45640
rect 57750 45528 57810 45540
rect 57750 45494 57778 45528
rect 57778 45494 57810 45528
rect 57750 45480 57810 45494
rect 58170 45410 58230 45470
rect 58590 45528 58650 45540
rect 58590 45494 58595 45528
rect 58595 45494 58629 45528
rect 58629 45494 58650 45528
rect 58590 45480 58650 45494
rect 57750 44128 57810 44140
rect 58170 44150 58230 44210
rect 57750 44094 57778 44128
rect 57778 44094 57810 44128
rect 57750 44080 57810 44094
rect 58590 44128 58650 44140
rect 58590 44094 58595 44128
rect 58595 44094 58629 44128
rect 58629 44094 58650 44128
rect 58590 44080 58650 44094
rect 58170 43980 58230 44040
rect 58170 43870 58230 43930
rect 57750 43818 57810 43830
rect 57750 43784 57778 43818
rect 57778 43784 57810 43818
rect 57750 43770 57810 43784
rect 58170 43700 58230 43760
rect 58590 43818 58650 43830
rect 58590 43784 58595 43818
rect 58595 43784 58629 43818
rect 58629 43784 58650 43818
rect 58590 43770 58650 43784
rect 57750 42418 57810 42430
rect 58170 42440 58230 42500
rect 57750 42384 57778 42418
rect 57778 42384 57810 42418
rect 57750 42370 57810 42384
rect 58590 42418 58650 42430
rect 58590 42384 58595 42418
rect 58595 42384 58629 42418
rect 58629 42384 58650 42418
rect 58590 42370 58650 42384
rect 58170 42270 58230 42330
rect 58170 42160 58230 42220
rect 57750 42108 57810 42120
rect 57750 42074 57778 42108
rect 57778 42074 57810 42108
rect 57750 42060 57810 42074
rect 58170 41990 58230 42050
rect 58590 42108 58650 42120
rect 58590 42074 58595 42108
rect 58595 42074 58629 42108
rect 58629 42074 58650 42108
rect 58590 42060 58650 42074
rect 57750 40708 57810 40720
rect 58170 40730 58230 40790
rect 57750 40674 57778 40708
rect 57778 40674 57810 40708
rect 57750 40660 57810 40674
rect 58590 40708 58650 40720
rect 58590 40674 58595 40708
rect 58595 40674 58629 40708
rect 58629 40674 58650 40708
rect 58590 40660 58650 40674
rect 58170 40560 58230 40620
rect 58170 40450 58230 40510
rect 57750 40398 57810 40410
rect 57750 40364 57778 40398
rect 57778 40364 57810 40398
rect 57750 40350 57810 40364
rect 58170 40280 58230 40340
rect 58590 40398 58650 40410
rect 58590 40364 58595 40398
rect 58595 40364 58629 40398
rect 58629 40364 58650 40398
rect 58590 40350 58650 40364
rect 57640 39620 57700 39680
rect 58710 39620 58770 39680
rect 58810 66410 58870 66470
rect 58870 65880 58930 65940
rect 58810 64700 58870 64760
rect 58870 64170 58930 64230
rect 58810 62990 58870 63050
rect 58870 62460 58930 62520
rect 58810 61280 58870 61340
rect 58870 60750 58930 60810
rect 58810 59570 58870 59630
rect 58870 59040 58930 59100
rect 58810 57860 58870 57920
rect 58870 57330 58930 57390
rect 58810 56150 58870 56210
rect 58870 55620 58930 55680
rect 58810 54440 58870 54500
rect 58870 53910 58930 53970
rect 58810 52730 58870 52790
rect 58870 52200 58930 52260
rect 58810 51020 58870 51080
rect 58870 50490 58930 50550
rect 58810 49310 58870 49370
rect 58870 48780 58930 48840
rect 58810 47600 58870 47660
rect 58870 47070 58930 47130
rect 58810 45890 58870 45950
rect 58870 45360 58930 45420
rect 58810 44180 58870 44240
rect 58870 43650 58930 43710
rect 58810 42470 58870 42530
rect 58870 41940 58930 42000
rect 58810 40760 58870 40820
rect 57340 39170 57400 39230
rect 58870 40230 58930 40290
rect 58870 39620 58930 39680
rect 58960 66320 59020 66380
rect 58960 64610 59020 64670
rect 59080 62900 59140 62960
rect 59080 61180 59140 61240
rect 59200 59480 59260 59540
rect 59320 57770 59380 57830
rect 59320 56060 59380 56120
rect 59320 54350 59380 54410
rect 59320 52640 59380 52700
rect 59320 50930 59380 50990
rect 59320 49220 59380 49280
rect 59200 47510 59260 47570
rect 59080 45800 59140 45860
rect 59080 44090 59140 44150
rect 58960 42380 59020 42440
rect 58960 40670 59020 40730
rect 62530 66320 62590 66380
rect 62530 64610 62590 64670
rect 62530 62900 62590 62960
rect 62530 61190 62590 61250
rect 62410 59480 62470 59540
rect 62410 57770 62470 57830
rect 62410 56060 62470 56120
rect 62410 54350 62470 54410
rect 62410 52640 62470 52700
rect 62410 50930 62470 50990
rect 62410 49220 62470 49280
rect 62410 47510 62470 47570
rect 59160 39170 59220 39230
rect 59340 39230 59400 39290
rect 59520 39290 59580 39350
rect 59700 39350 59760 39410
rect 62530 45800 62590 45860
rect 62530 44090 62590 44150
rect 62530 42380 62590 42440
rect 62530 40670 62590 40730
rect 62150 39230 62210 39290
rect 62740 66358 62800 66370
rect 63160 66380 63220 66440
rect 62740 66324 62768 66358
rect 62768 66324 62800 66358
rect 62740 66310 62800 66324
rect 63580 66358 63640 66370
rect 63580 66324 63585 66358
rect 63585 66324 63619 66358
rect 63619 66324 63640 66358
rect 63580 66310 63640 66324
rect 63160 66210 63220 66270
rect 63160 66100 63220 66160
rect 62740 66048 62800 66060
rect 62740 66014 62768 66048
rect 62768 66014 62800 66048
rect 62740 66000 62800 66014
rect 63160 65930 63220 65990
rect 63580 66048 63640 66060
rect 63580 66014 63585 66048
rect 63585 66014 63619 66048
rect 63619 66014 63640 66048
rect 63580 66000 63640 66014
rect 62740 64648 62800 64660
rect 63160 64670 63220 64730
rect 62740 64614 62768 64648
rect 62768 64614 62800 64648
rect 62740 64600 62800 64614
rect 63580 64648 63640 64660
rect 63580 64614 63585 64648
rect 63585 64614 63619 64648
rect 63619 64614 63640 64648
rect 63580 64600 63640 64614
rect 63160 64500 63220 64560
rect 63160 64390 63220 64450
rect 62740 64338 62800 64350
rect 62740 64304 62768 64338
rect 62768 64304 62800 64338
rect 62740 64290 62800 64304
rect 63160 64220 63220 64280
rect 63580 64338 63640 64350
rect 63580 64304 63585 64338
rect 63585 64304 63619 64338
rect 63619 64304 63640 64338
rect 63580 64290 63640 64304
rect 62740 62938 62800 62950
rect 63160 62960 63220 63020
rect 62740 62904 62768 62938
rect 62768 62904 62800 62938
rect 62740 62890 62800 62904
rect 63580 62938 63640 62950
rect 63580 62904 63585 62938
rect 63585 62904 63619 62938
rect 63619 62904 63640 62938
rect 63580 62890 63640 62904
rect 63160 62790 63220 62850
rect 63160 62680 63220 62740
rect 62740 62628 62800 62640
rect 62740 62594 62768 62628
rect 62768 62594 62800 62628
rect 62740 62580 62800 62594
rect 63160 62510 63220 62570
rect 63580 62628 63640 62640
rect 63580 62594 63585 62628
rect 63585 62594 63619 62628
rect 63619 62594 63640 62628
rect 63580 62580 63640 62594
rect 62740 61228 62800 61240
rect 63160 61250 63220 61310
rect 62740 61194 62768 61228
rect 62768 61194 62800 61228
rect 62740 61180 62800 61194
rect 63580 61228 63640 61240
rect 63580 61194 63585 61228
rect 63585 61194 63619 61228
rect 63619 61194 63640 61228
rect 63580 61180 63640 61194
rect 63160 61080 63220 61140
rect 63160 60970 63220 61030
rect 62740 60918 62800 60930
rect 62740 60884 62768 60918
rect 62768 60884 62800 60918
rect 62740 60870 62800 60884
rect 63160 60800 63220 60860
rect 63580 60918 63640 60930
rect 63580 60884 63585 60918
rect 63585 60884 63619 60918
rect 63619 60884 63640 60918
rect 63580 60870 63640 60884
rect 62740 59518 62800 59530
rect 63160 59540 63220 59600
rect 62740 59484 62768 59518
rect 62768 59484 62800 59518
rect 62740 59470 62800 59484
rect 63580 59518 63640 59530
rect 63580 59484 63585 59518
rect 63585 59484 63619 59518
rect 63619 59484 63640 59518
rect 63580 59470 63640 59484
rect 63160 59370 63220 59430
rect 63160 59260 63220 59320
rect 62740 59208 62800 59220
rect 62740 59174 62768 59208
rect 62768 59174 62800 59208
rect 62740 59160 62800 59174
rect 63160 59090 63220 59150
rect 63580 59208 63640 59220
rect 63580 59174 63585 59208
rect 63585 59174 63619 59208
rect 63619 59174 63640 59208
rect 63580 59160 63640 59174
rect 62740 57808 62800 57820
rect 63160 57830 63220 57890
rect 62740 57774 62768 57808
rect 62768 57774 62800 57808
rect 62740 57760 62800 57774
rect 63580 57808 63640 57820
rect 63580 57774 63585 57808
rect 63585 57774 63619 57808
rect 63619 57774 63640 57808
rect 63580 57760 63640 57774
rect 63160 57660 63220 57720
rect 63160 57550 63220 57610
rect 62740 57498 62800 57510
rect 62740 57464 62768 57498
rect 62768 57464 62800 57498
rect 62740 57450 62800 57464
rect 63160 57380 63220 57440
rect 63580 57498 63640 57510
rect 63580 57464 63585 57498
rect 63585 57464 63619 57498
rect 63619 57464 63640 57498
rect 63580 57450 63640 57464
rect 62740 56098 62800 56110
rect 63160 56120 63220 56180
rect 62740 56064 62768 56098
rect 62768 56064 62800 56098
rect 62740 56050 62800 56064
rect 63580 56098 63640 56110
rect 63580 56064 63585 56098
rect 63585 56064 63619 56098
rect 63619 56064 63640 56098
rect 63580 56050 63640 56064
rect 63160 55950 63220 56010
rect 63160 55840 63220 55900
rect 62740 55788 62800 55800
rect 62740 55754 62768 55788
rect 62768 55754 62800 55788
rect 62740 55740 62800 55754
rect 63160 55670 63220 55730
rect 63580 55788 63640 55800
rect 63580 55754 63585 55788
rect 63585 55754 63619 55788
rect 63619 55754 63640 55788
rect 63580 55740 63640 55754
rect 62740 54388 62800 54400
rect 63160 54410 63220 54470
rect 62740 54354 62768 54388
rect 62768 54354 62800 54388
rect 62740 54340 62800 54354
rect 63580 54388 63640 54400
rect 63580 54354 63585 54388
rect 63585 54354 63619 54388
rect 63619 54354 63640 54388
rect 63580 54340 63640 54354
rect 63160 54240 63220 54300
rect 63160 54130 63220 54190
rect 62740 54078 62800 54090
rect 62740 54044 62768 54078
rect 62768 54044 62800 54078
rect 62740 54030 62800 54044
rect 63160 53960 63220 54020
rect 63580 54078 63640 54090
rect 63580 54044 63585 54078
rect 63585 54044 63619 54078
rect 63619 54044 63640 54078
rect 63580 54030 63640 54044
rect 62740 52678 62800 52690
rect 63160 52700 63220 52760
rect 62740 52644 62768 52678
rect 62768 52644 62800 52678
rect 62740 52630 62800 52644
rect 63580 52678 63640 52690
rect 63580 52644 63585 52678
rect 63585 52644 63619 52678
rect 63619 52644 63640 52678
rect 63580 52630 63640 52644
rect 63160 52530 63220 52590
rect 63160 52420 63220 52480
rect 62740 52368 62800 52380
rect 62740 52334 62768 52368
rect 62768 52334 62800 52368
rect 62740 52320 62800 52334
rect 63160 52250 63220 52310
rect 63580 52368 63640 52380
rect 63580 52334 63585 52368
rect 63585 52334 63619 52368
rect 63619 52334 63640 52368
rect 63580 52320 63640 52334
rect 62740 50968 62800 50980
rect 63160 50990 63220 51050
rect 62740 50934 62768 50968
rect 62768 50934 62800 50968
rect 62740 50920 62800 50934
rect 63580 50968 63640 50980
rect 63580 50934 63585 50968
rect 63585 50934 63619 50968
rect 63619 50934 63640 50968
rect 63580 50920 63640 50934
rect 63160 50820 63220 50880
rect 63160 50710 63220 50770
rect 62740 50658 62800 50670
rect 62740 50624 62768 50658
rect 62768 50624 62800 50658
rect 62740 50610 62800 50624
rect 63160 50540 63220 50600
rect 63580 50658 63640 50670
rect 63580 50624 63585 50658
rect 63585 50624 63619 50658
rect 63619 50624 63640 50658
rect 63580 50610 63640 50624
rect 62740 49258 62800 49270
rect 63160 49280 63220 49340
rect 62740 49224 62768 49258
rect 62768 49224 62800 49258
rect 62740 49210 62800 49224
rect 63580 49258 63640 49270
rect 63580 49224 63585 49258
rect 63585 49224 63619 49258
rect 63619 49224 63640 49258
rect 63580 49210 63640 49224
rect 63160 49110 63220 49170
rect 63160 49000 63220 49060
rect 62740 48948 62800 48960
rect 62740 48914 62768 48948
rect 62768 48914 62800 48948
rect 62740 48900 62800 48914
rect 63160 48830 63220 48890
rect 63580 48948 63640 48960
rect 63580 48914 63585 48948
rect 63585 48914 63619 48948
rect 63619 48914 63640 48948
rect 63580 48900 63640 48914
rect 62740 47548 62800 47560
rect 63160 47570 63220 47630
rect 62740 47514 62768 47548
rect 62768 47514 62800 47548
rect 62740 47500 62800 47514
rect 63580 47548 63640 47560
rect 63580 47514 63585 47548
rect 63585 47514 63619 47548
rect 63619 47514 63640 47548
rect 63580 47500 63640 47514
rect 63160 47400 63220 47460
rect 63160 47290 63220 47350
rect 62740 47238 62800 47250
rect 62740 47204 62768 47238
rect 62768 47204 62800 47238
rect 62740 47190 62800 47204
rect 63160 47120 63220 47180
rect 63580 47238 63640 47250
rect 63580 47204 63585 47238
rect 63585 47204 63619 47238
rect 63619 47204 63640 47238
rect 63580 47190 63640 47204
rect 62740 45838 62800 45850
rect 63160 45860 63220 45920
rect 62740 45804 62768 45838
rect 62768 45804 62800 45838
rect 62740 45790 62800 45804
rect 63580 45838 63640 45850
rect 63580 45804 63585 45838
rect 63585 45804 63619 45838
rect 63619 45804 63640 45838
rect 63580 45790 63640 45804
rect 63160 45690 63220 45750
rect 63160 45580 63220 45640
rect 62740 45528 62800 45540
rect 62740 45494 62768 45528
rect 62768 45494 62800 45528
rect 62740 45480 62800 45494
rect 63160 45410 63220 45470
rect 63580 45528 63640 45540
rect 63580 45494 63585 45528
rect 63585 45494 63619 45528
rect 63619 45494 63640 45528
rect 63580 45480 63640 45494
rect 62740 44128 62800 44140
rect 63160 44150 63220 44210
rect 62740 44094 62768 44128
rect 62768 44094 62800 44128
rect 62740 44080 62800 44094
rect 63580 44128 63640 44140
rect 63580 44094 63585 44128
rect 63585 44094 63619 44128
rect 63619 44094 63640 44128
rect 63580 44080 63640 44094
rect 63160 43980 63220 44040
rect 63160 43870 63220 43930
rect 62740 43818 62800 43830
rect 62740 43784 62768 43818
rect 62768 43784 62800 43818
rect 62740 43770 62800 43784
rect 63160 43700 63220 43760
rect 63580 43818 63640 43830
rect 63580 43784 63585 43818
rect 63585 43784 63619 43818
rect 63619 43784 63640 43818
rect 63580 43770 63640 43784
rect 62740 42418 62800 42430
rect 63160 42440 63220 42500
rect 62740 42384 62768 42418
rect 62768 42384 62800 42418
rect 62740 42370 62800 42384
rect 63580 42418 63640 42430
rect 63580 42384 63585 42418
rect 63585 42384 63619 42418
rect 63619 42384 63640 42418
rect 63580 42370 63640 42384
rect 63160 42270 63220 42330
rect 63160 42160 63220 42220
rect 62740 42108 62800 42120
rect 62740 42074 62768 42108
rect 62768 42074 62800 42108
rect 62740 42060 62800 42074
rect 63160 41990 63220 42050
rect 63580 42108 63640 42120
rect 63580 42074 63585 42108
rect 63585 42074 63619 42108
rect 63619 42074 63640 42108
rect 63580 42060 63640 42074
rect 62740 40708 62800 40720
rect 63160 40730 63220 40790
rect 62740 40674 62768 40708
rect 62768 40674 62800 40708
rect 62740 40660 62800 40674
rect 63580 40708 63640 40720
rect 63580 40674 63585 40708
rect 63585 40674 63619 40708
rect 63619 40674 63640 40708
rect 63580 40660 63640 40674
rect 63160 40560 63220 40620
rect 63160 40450 63220 40510
rect 62740 40398 62800 40410
rect 62740 40364 62768 40398
rect 62768 40364 62800 40398
rect 62740 40350 62800 40364
rect 63160 40280 63220 40340
rect 63580 40398 63640 40410
rect 63580 40364 63585 40398
rect 63585 40364 63619 40398
rect 63619 40364 63640 40398
rect 63580 40350 63640 40364
rect 62630 39620 62690 39680
rect 63700 39620 63760 39680
rect 63800 66410 63860 66470
rect 63860 65880 63920 65940
rect 63800 64700 63860 64760
rect 63860 64170 63920 64230
rect 63800 62990 63860 63050
rect 63860 62460 63920 62520
rect 63800 61280 63860 61340
rect 63860 60750 63920 60810
rect 63800 59570 63860 59630
rect 63860 59040 63920 59100
rect 63800 57860 63860 57920
rect 63860 57330 63920 57390
rect 63800 56150 63860 56210
rect 63860 55620 63920 55680
rect 63800 54440 63860 54500
rect 63860 53910 63920 53970
rect 63800 52730 63860 52790
rect 63860 52200 63920 52260
rect 63800 51020 63860 51080
rect 63860 50490 63920 50550
rect 63800 49310 63860 49370
rect 63860 48780 63920 48840
rect 63800 47600 63860 47660
rect 63860 47070 63920 47130
rect 63800 45890 63860 45950
rect 63860 45360 63920 45420
rect 63800 44180 63860 44240
rect 63860 43650 63920 43710
rect 63800 42470 63860 42530
rect 63860 41940 63920 42000
rect 63800 40760 63860 40820
rect 62330 39170 62390 39230
rect 63860 40230 63920 40290
rect 63860 39620 63920 39680
rect 63950 66320 64010 66380
rect 63950 64610 64010 64670
rect 63950 62900 64010 62960
rect 63950 61190 64010 61250
rect 64070 59480 64130 59540
rect 64070 57770 64130 57830
rect 64070 56060 64130 56120
rect 64070 54350 64130 54410
rect 64070 52640 64130 52700
rect 64070 50930 64130 50990
rect 64070 49220 64130 49280
rect 64070 47510 64130 47570
rect 63950 45800 64010 45860
rect 63950 44090 64010 44150
rect 63950 42380 64010 42440
rect 63950 40670 64010 40730
rect 67520 66320 67580 66380
rect 67520 64610 67580 64670
rect 67520 62900 67580 62960
rect 67520 61190 67580 61250
rect 67400 59480 67460 59540
rect 67400 57770 67460 57830
rect 67400 56060 67460 56120
rect 67400 54350 67460 54410
rect 67400 52640 67460 52700
rect 67400 50930 67460 50990
rect 67400 49220 67460 49280
rect 67400 47510 67460 47570
rect 67520 45800 67580 45860
rect 67520 44090 67580 44150
rect 67520 42380 67580 42440
rect 67520 40670 67580 40730
rect 64150 39170 64210 39230
rect 64330 39230 64390 39290
rect 67140 39230 67200 39290
rect 67730 66358 67790 66370
rect 68150 66380 68210 66440
rect 67730 66324 67758 66358
rect 67758 66324 67790 66358
rect 67730 66310 67790 66324
rect 68570 66358 68630 66370
rect 68570 66324 68575 66358
rect 68575 66324 68609 66358
rect 68609 66324 68630 66358
rect 68570 66310 68630 66324
rect 68150 66210 68210 66270
rect 68150 66100 68210 66160
rect 67730 66048 67790 66060
rect 67730 66014 67758 66048
rect 67758 66014 67790 66048
rect 67730 66000 67790 66014
rect 68150 65930 68210 65990
rect 68570 66048 68630 66060
rect 68570 66014 68575 66048
rect 68575 66014 68609 66048
rect 68609 66014 68630 66048
rect 68570 66000 68630 66014
rect 67730 64648 67790 64660
rect 68150 64670 68210 64730
rect 67730 64614 67758 64648
rect 67758 64614 67790 64648
rect 67730 64600 67790 64614
rect 68570 64648 68630 64660
rect 68570 64614 68575 64648
rect 68575 64614 68609 64648
rect 68609 64614 68630 64648
rect 68570 64600 68630 64614
rect 68150 64500 68210 64560
rect 68150 64390 68210 64450
rect 67730 64338 67790 64350
rect 67730 64304 67758 64338
rect 67758 64304 67790 64338
rect 67730 64290 67790 64304
rect 68150 64220 68210 64280
rect 68570 64338 68630 64350
rect 68570 64304 68575 64338
rect 68575 64304 68609 64338
rect 68609 64304 68630 64338
rect 68570 64290 68630 64304
rect 67730 62938 67790 62950
rect 68150 62960 68210 63020
rect 67730 62904 67758 62938
rect 67758 62904 67790 62938
rect 67730 62890 67790 62904
rect 68570 62938 68630 62950
rect 68570 62904 68575 62938
rect 68575 62904 68609 62938
rect 68609 62904 68630 62938
rect 68570 62890 68630 62904
rect 68150 62790 68210 62850
rect 68150 62680 68210 62740
rect 67730 62628 67790 62640
rect 67730 62594 67758 62628
rect 67758 62594 67790 62628
rect 67730 62580 67790 62594
rect 68150 62510 68210 62570
rect 68570 62628 68630 62640
rect 68570 62594 68575 62628
rect 68575 62594 68609 62628
rect 68609 62594 68630 62628
rect 68570 62580 68630 62594
rect 67730 61228 67790 61240
rect 68150 61250 68210 61310
rect 67730 61194 67758 61228
rect 67758 61194 67790 61228
rect 67730 61180 67790 61194
rect 68570 61228 68630 61240
rect 68570 61194 68575 61228
rect 68575 61194 68609 61228
rect 68609 61194 68630 61228
rect 68570 61180 68630 61194
rect 68150 61080 68210 61140
rect 68150 60970 68210 61030
rect 67730 60918 67790 60930
rect 67730 60884 67758 60918
rect 67758 60884 67790 60918
rect 67730 60870 67790 60884
rect 68150 60800 68210 60860
rect 68570 60918 68630 60930
rect 68570 60884 68575 60918
rect 68575 60884 68609 60918
rect 68609 60884 68630 60918
rect 68570 60870 68630 60884
rect 67730 59518 67790 59530
rect 68150 59540 68210 59600
rect 67730 59484 67758 59518
rect 67758 59484 67790 59518
rect 67730 59470 67790 59484
rect 68570 59518 68630 59530
rect 68570 59484 68575 59518
rect 68575 59484 68609 59518
rect 68609 59484 68630 59518
rect 68570 59470 68630 59484
rect 68150 59370 68210 59430
rect 68150 59260 68210 59320
rect 67730 59208 67790 59220
rect 67730 59174 67758 59208
rect 67758 59174 67790 59208
rect 67730 59160 67790 59174
rect 68150 59090 68210 59150
rect 68570 59208 68630 59220
rect 68570 59174 68575 59208
rect 68575 59174 68609 59208
rect 68609 59174 68630 59208
rect 68570 59160 68630 59174
rect 67730 57808 67790 57820
rect 68150 57830 68210 57890
rect 67730 57774 67758 57808
rect 67758 57774 67790 57808
rect 67730 57760 67790 57774
rect 68570 57808 68630 57820
rect 68570 57774 68575 57808
rect 68575 57774 68609 57808
rect 68609 57774 68630 57808
rect 68570 57760 68630 57774
rect 68150 57660 68210 57720
rect 68150 57550 68210 57610
rect 67730 57498 67790 57510
rect 67730 57464 67758 57498
rect 67758 57464 67790 57498
rect 67730 57450 67790 57464
rect 68150 57380 68210 57440
rect 68570 57498 68630 57510
rect 68570 57464 68575 57498
rect 68575 57464 68609 57498
rect 68609 57464 68630 57498
rect 68570 57450 68630 57464
rect 67730 56098 67790 56110
rect 68150 56120 68210 56180
rect 67730 56064 67758 56098
rect 67758 56064 67790 56098
rect 67730 56050 67790 56064
rect 68570 56098 68630 56110
rect 68570 56064 68575 56098
rect 68575 56064 68609 56098
rect 68609 56064 68630 56098
rect 68570 56050 68630 56064
rect 68150 55950 68210 56010
rect 68150 55840 68210 55900
rect 67730 55788 67790 55800
rect 67730 55754 67758 55788
rect 67758 55754 67790 55788
rect 67730 55740 67790 55754
rect 68150 55670 68210 55730
rect 68570 55788 68630 55800
rect 68570 55754 68575 55788
rect 68575 55754 68609 55788
rect 68609 55754 68630 55788
rect 68570 55740 68630 55754
rect 67730 54388 67790 54400
rect 68150 54410 68210 54470
rect 67730 54354 67758 54388
rect 67758 54354 67790 54388
rect 67730 54340 67790 54354
rect 68570 54388 68630 54400
rect 68570 54354 68575 54388
rect 68575 54354 68609 54388
rect 68609 54354 68630 54388
rect 68570 54340 68630 54354
rect 68150 54240 68210 54300
rect 68150 54130 68210 54190
rect 67730 54078 67790 54090
rect 67730 54044 67758 54078
rect 67758 54044 67790 54078
rect 67730 54030 67790 54044
rect 68150 53960 68210 54020
rect 68570 54078 68630 54090
rect 68570 54044 68575 54078
rect 68575 54044 68609 54078
rect 68609 54044 68630 54078
rect 68570 54030 68630 54044
rect 67730 52678 67790 52690
rect 68150 52700 68210 52760
rect 67730 52644 67758 52678
rect 67758 52644 67790 52678
rect 67730 52630 67790 52644
rect 68570 52678 68630 52690
rect 68570 52644 68575 52678
rect 68575 52644 68609 52678
rect 68609 52644 68630 52678
rect 68570 52630 68630 52644
rect 68150 52530 68210 52590
rect 68150 52420 68210 52480
rect 67730 52368 67790 52380
rect 67730 52334 67758 52368
rect 67758 52334 67790 52368
rect 67730 52320 67790 52334
rect 68150 52250 68210 52310
rect 68570 52368 68630 52380
rect 68570 52334 68575 52368
rect 68575 52334 68609 52368
rect 68609 52334 68630 52368
rect 68570 52320 68630 52334
rect 67730 50968 67790 50980
rect 68150 50990 68210 51050
rect 67730 50934 67758 50968
rect 67758 50934 67790 50968
rect 67730 50920 67790 50934
rect 68570 50968 68630 50980
rect 68570 50934 68575 50968
rect 68575 50934 68609 50968
rect 68609 50934 68630 50968
rect 68570 50920 68630 50934
rect 68150 50820 68210 50880
rect 68150 50710 68210 50770
rect 67730 50658 67790 50670
rect 67730 50624 67758 50658
rect 67758 50624 67790 50658
rect 67730 50610 67790 50624
rect 68150 50540 68210 50600
rect 68570 50658 68630 50670
rect 68570 50624 68575 50658
rect 68575 50624 68609 50658
rect 68609 50624 68630 50658
rect 68570 50610 68630 50624
rect 67730 49258 67790 49270
rect 68150 49280 68210 49340
rect 67730 49224 67758 49258
rect 67758 49224 67790 49258
rect 67730 49210 67790 49224
rect 68570 49258 68630 49270
rect 68570 49224 68575 49258
rect 68575 49224 68609 49258
rect 68609 49224 68630 49258
rect 68570 49210 68630 49224
rect 68150 49110 68210 49170
rect 68150 49000 68210 49060
rect 67730 48948 67790 48960
rect 67730 48914 67758 48948
rect 67758 48914 67790 48948
rect 67730 48900 67790 48914
rect 68150 48830 68210 48890
rect 68570 48948 68630 48960
rect 68570 48914 68575 48948
rect 68575 48914 68609 48948
rect 68609 48914 68630 48948
rect 68570 48900 68630 48914
rect 67730 47548 67790 47560
rect 68150 47570 68210 47630
rect 67730 47514 67758 47548
rect 67758 47514 67790 47548
rect 67730 47500 67790 47514
rect 68570 47548 68630 47560
rect 68570 47514 68575 47548
rect 68575 47514 68609 47548
rect 68609 47514 68630 47548
rect 68570 47500 68630 47514
rect 68150 47400 68210 47460
rect 68150 47290 68210 47350
rect 67730 47238 67790 47250
rect 67730 47204 67758 47238
rect 67758 47204 67790 47238
rect 67730 47190 67790 47204
rect 68150 47120 68210 47180
rect 68570 47238 68630 47250
rect 68570 47204 68575 47238
rect 68575 47204 68609 47238
rect 68609 47204 68630 47238
rect 68570 47190 68630 47204
rect 67730 45838 67790 45850
rect 68150 45860 68210 45920
rect 67730 45804 67758 45838
rect 67758 45804 67790 45838
rect 67730 45790 67790 45804
rect 68570 45838 68630 45850
rect 68570 45804 68575 45838
rect 68575 45804 68609 45838
rect 68609 45804 68630 45838
rect 68570 45790 68630 45804
rect 68150 45690 68210 45750
rect 68150 45580 68210 45640
rect 67730 45528 67790 45540
rect 67730 45494 67758 45528
rect 67758 45494 67790 45528
rect 67730 45480 67790 45494
rect 68150 45410 68210 45470
rect 68570 45528 68630 45540
rect 68570 45494 68575 45528
rect 68575 45494 68609 45528
rect 68609 45494 68630 45528
rect 68570 45480 68630 45494
rect 67730 44128 67790 44140
rect 68150 44150 68210 44210
rect 67730 44094 67758 44128
rect 67758 44094 67790 44128
rect 67730 44080 67790 44094
rect 68570 44128 68630 44140
rect 68570 44094 68575 44128
rect 68575 44094 68609 44128
rect 68609 44094 68630 44128
rect 68570 44080 68630 44094
rect 68150 43980 68210 44040
rect 68150 43870 68210 43930
rect 67730 43818 67790 43830
rect 67730 43784 67758 43818
rect 67758 43784 67790 43818
rect 67730 43770 67790 43784
rect 68150 43700 68210 43760
rect 68570 43818 68630 43830
rect 68570 43784 68575 43818
rect 68575 43784 68609 43818
rect 68609 43784 68630 43818
rect 68570 43770 68630 43784
rect 67730 42418 67790 42430
rect 68150 42440 68210 42500
rect 67730 42384 67758 42418
rect 67758 42384 67790 42418
rect 67730 42370 67790 42384
rect 68570 42418 68630 42430
rect 68570 42384 68575 42418
rect 68575 42384 68609 42418
rect 68609 42384 68630 42418
rect 68570 42370 68630 42384
rect 68150 42270 68210 42330
rect 68150 42160 68210 42220
rect 67730 42108 67790 42120
rect 67730 42074 67758 42108
rect 67758 42074 67790 42108
rect 67730 42060 67790 42074
rect 68150 41990 68210 42050
rect 68570 42108 68630 42120
rect 68570 42074 68575 42108
rect 68575 42074 68609 42108
rect 68609 42074 68630 42108
rect 68570 42060 68630 42074
rect 67730 40708 67790 40720
rect 68150 40730 68210 40790
rect 67730 40674 67758 40708
rect 67758 40674 67790 40708
rect 67730 40660 67790 40674
rect 68570 40708 68630 40720
rect 68570 40674 68575 40708
rect 68575 40674 68609 40708
rect 68609 40674 68630 40708
rect 68570 40660 68630 40674
rect 68150 40560 68210 40620
rect 68150 40450 68210 40510
rect 67730 40398 67790 40410
rect 67730 40364 67758 40398
rect 67758 40364 67790 40398
rect 67730 40350 67790 40364
rect 68150 40280 68210 40340
rect 68570 40398 68630 40410
rect 68570 40364 68575 40398
rect 68575 40364 68609 40398
rect 68609 40364 68630 40398
rect 68570 40350 68630 40364
rect 67620 39620 67680 39680
rect 68690 39620 68750 39680
rect 68790 66410 68850 66470
rect 68850 65880 68910 65940
rect 68790 64700 68850 64760
rect 68850 64170 68910 64230
rect 68790 62990 68850 63050
rect 68850 62460 68910 62520
rect 68790 61280 68850 61340
rect 68850 60750 68910 60810
rect 68790 59570 68850 59630
rect 68850 59040 68910 59100
rect 68790 57860 68850 57920
rect 68850 57330 68910 57390
rect 68790 56150 68850 56210
rect 68850 55620 68910 55680
rect 68790 54440 68850 54500
rect 68850 53910 68910 53970
rect 68790 52730 68850 52790
rect 68850 52200 68910 52260
rect 68790 51020 68850 51080
rect 68850 50490 68910 50550
rect 68790 49310 68850 49370
rect 68850 48780 68910 48840
rect 68790 47600 68850 47660
rect 68850 47070 68910 47130
rect 68790 45890 68850 45950
rect 68850 45360 68910 45420
rect 68790 44180 68850 44240
rect 68850 43650 68910 43710
rect 68790 42470 68850 42530
rect 68850 41940 68910 42000
rect 68790 40760 68850 40820
rect 67320 39170 67380 39230
rect 68850 40230 68910 40290
rect 68850 39620 68910 39680
rect 68940 66320 69000 66380
rect 68940 64610 69000 64670
rect 68940 62900 69000 62960
rect 68940 61190 69000 61250
rect 69060 59480 69120 59540
rect 69060 57770 69120 57830
rect 69060 56060 69120 56120
rect 69060 54350 69120 54410
rect 69060 52640 69120 52700
rect 69060 50930 69120 50990
rect 69060 49220 69120 49280
rect 69060 47510 69120 47570
rect 68940 45800 69000 45860
rect 68940 44090 69000 44150
rect 68940 42380 69000 42440
rect 68940 40670 69000 40730
rect 72510 66320 72570 66380
rect 72510 64610 72570 64670
rect 72510 62900 72570 62960
rect 72510 61190 72570 61250
rect 72510 59480 72570 59540
rect 72510 57770 72570 57830
rect 72510 56060 72570 56120
rect 72510 54350 72570 54410
rect 72510 52640 72570 52700
rect 72510 50930 72570 50990
rect 72510 49220 72570 49280
rect 72510 47510 72570 47570
rect 72510 45800 72570 45860
rect 72510 44090 72570 44150
rect 72510 42380 72570 42440
rect 72510 40670 72570 40730
rect 69140 39170 69200 39230
rect 69320 39230 69380 39290
rect 72720 66358 72780 66370
rect 73140 66380 73200 66440
rect 72720 66324 72748 66358
rect 72748 66324 72780 66358
rect 72720 66310 72780 66324
rect 73560 66358 73620 66370
rect 73560 66324 73565 66358
rect 73565 66324 73599 66358
rect 73599 66324 73620 66358
rect 73560 66310 73620 66324
rect 73140 66210 73200 66270
rect 73140 66100 73200 66160
rect 72720 66048 72780 66060
rect 72720 66014 72748 66048
rect 72748 66014 72780 66048
rect 72720 66000 72780 66014
rect 73140 65930 73200 65990
rect 73560 66048 73620 66060
rect 73560 66014 73565 66048
rect 73565 66014 73599 66048
rect 73599 66014 73620 66048
rect 73560 66000 73620 66014
rect 72720 64648 72780 64660
rect 73140 64670 73200 64730
rect 72720 64614 72748 64648
rect 72748 64614 72780 64648
rect 72720 64600 72780 64614
rect 73560 64648 73620 64660
rect 73560 64614 73565 64648
rect 73565 64614 73599 64648
rect 73599 64614 73620 64648
rect 73560 64600 73620 64614
rect 73140 64500 73200 64560
rect 73140 64390 73200 64450
rect 72720 64338 72780 64350
rect 72720 64304 72748 64338
rect 72748 64304 72780 64338
rect 72720 64290 72780 64304
rect 73140 64220 73200 64280
rect 73560 64338 73620 64350
rect 73560 64304 73565 64338
rect 73565 64304 73599 64338
rect 73599 64304 73620 64338
rect 73560 64290 73620 64304
rect 72720 62938 72780 62950
rect 73140 62960 73200 63020
rect 72720 62904 72748 62938
rect 72748 62904 72780 62938
rect 72720 62890 72780 62904
rect 73560 62938 73620 62950
rect 73560 62904 73565 62938
rect 73565 62904 73599 62938
rect 73599 62904 73620 62938
rect 73560 62890 73620 62904
rect 73140 62790 73200 62850
rect 73140 62680 73200 62740
rect 72720 62628 72780 62640
rect 72720 62594 72748 62628
rect 72748 62594 72780 62628
rect 72720 62580 72780 62594
rect 73140 62510 73200 62570
rect 73560 62628 73620 62640
rect 73560 62594 73565 62628
rect 73565 62594 73599 62628
rect 73599 62594 73620 62628
rect 73560 62580 73620 62594
rect 72720 61228 72780 61240
rect 73140 61250 73200 61310
rect 72720 61194 72748 61228
rect 72748 61194 72780 61228
rect 72720 61180 72780 61194
rect 73560 61228 73620 61240
rect 73560 61194 73565 61228
rect 73565 61194 73599 61228
rect 73599 61194 73620 61228
rect 73560 61180 73620 61194
rect 73140 61080 73200 61140
rect 73140 60970 73200 61030
rect 72720 60918 72780 60930
rect 72720 60884 72748 60918
rect 72748 60884 72780 60918
rect 72720 60870 72780 60884
rect 73140 60800 73200 60860
rect 73560 60918 73620 60930
rect 73560 60884 73565 60918
rect 73565 60884 73599 60918
rect 73599 60884 73620 60918
rect 73560 60870 73620 60884
rect 72720 59518 72780 59530
rect 73140 59540 73200 59600
rect 72720 59484 72748 59518
rect 72748 59484 72780 59518
rect 72720 59470 72780 59484
rect 73560 59518 73620 59530
rect 73560 59484 73565 59518
rect 73565 59484 73599 59518
rect 73599 59484 73620 59518
rect 73560 59470 73620 59484
rect 73140 59370 73200 59430
rect 73140 59260 73200 59320
rect 72720 59208 72780 59220
rect 72720 59174 72748 59208
rect 72748 59174 72780 59208
rect 72720 59160 72780 59174
rect 73140 59090 73200 59150
rect 73560 59208 73620 59220
rect 73560 59174 73565 59208
rect 73565 59174 73599 59208
rect 73599 59174 73620 59208
rect 73560 59160 73620 59174
rect 72720 57808 72780 57820
rect 73140 57830 73200 57890
rect 72720 57774 72748 57808
rect 72748 57774 72780 57808
rect 72720 57760 72780 57774
rect 73560 57808 73620 57820
rect 73560 57774 73565 57808
rect 73565 57774 73599 57808
rect 73599 57774 73620 57808
rect 73560 57760 73620 57774
rect 73140 57660 73200 57720
rect 73140 57550 73200 57610
rect 72720 57498 72780 57510
rect 72720 57464 72748 57498
rect 72748 57464 72780 57498
rect 72720 57450 72780 57464
rect 73140 57380 73200 57440
rect 73560 57498 73620 57510
rect 73560 57464 73565 57498
rect 73565 57464 73599 57498
rect 73599 57464 73620 57498
rect 73560 57450 73620 57464
rect 72720 56098 72780 56110
rect 73140 56120 73200 56180
rect 72720 56064 72748 56098
rect 72748 56064 72780 56098
rect 72720 56050 72780 56064
rect 73560 56098 73620 56110
rect 73560 56064 73565 56098
rect 73565 56064 73599 56098
rect 73599 56064 73620 56098
rect 73560 56050 73620 56064
rect 73140 55950 73200 56010
rect 73140 55840 73200 55900
rect 72720 55788 72780 55800
rect 72720 55754 72748 55788
rect 72748 55754 72780 55788
rect 72720 55740 72780 55754
rect 73140 55670 73200 55730
rect 73560 55788 73620 55800
rect 73560 55754 73565 55788
rect 73565 55754 73599 55788
rect 73599 55754 73620 55788
rect 73560 55740 73620 55754
rect 72720 54388 72780 54400
rect 73140 54410 73200 54470
rect 72720 54354 72748 54388
rect 72748 54354 72780 54388
rect 72720 54340 72780 54354
rect 73560 54388 73620 54400
rect 73560 54354 73565 54388
rect 73565 54354 73599 54388
rect 73599 54354 73620 54388
rect 73560 54340 73620 54354
rect 73140 54240 73200 54300
rect 73140 54130 73200 54190
rect 72720 54078 72780 54090
rect 72720 54044 72748 54078
rect 72748 54044 72780 54078
rect 72720 54030 72780 54044
rect 73140 53960 73200 54020
rect 73560 54078 73620 54090
rect 73560 54044 73565 54078
rect 73565 54044 73599 54078
rect 73599 54044 73620 54078
rect 73560 54030 73620 54044
rect 72720 52678 72780 52690
rect 73140 52700 73200 52760
rect 72720 52644 72748 52678
rect 72748 52644 72780 52678
rect 72720 52630 72780 52644
rect 73560 52678 73620 52690
rect 73560 52644 73565 52678
rect 73565 52644 73599 52678
rect 73599 52644 73620 52678
rect 73560 52630 73620 52644
rect 73140 52530 73200 52590
rect 73140 52420 73200 52480
rect 72720 52368 72780 52380
rect 72720 52334 72748 52368
rect 72748 52334 72780 52368
rect 72720 52320 72780 52334
rect 73140 52250 73200 52310
rect 73560 52368 73620 52380
rect 73560 52334 73565 52368
rect 73565 52334 73599 52368
rect 73599 52334 73620 52368
rect 73560 52320 73620 52334
rect 72720 50968 72780 50980
rect 73140 50990 73200 51050
rect 72720 50934 72748 50968
rect 72748 50934 72780 50968
rect 72720 50920 72780 50934
rect 73560 50968 73620 50980
rect 73560 50934 73565 50968
rect 73565 50934 73599 50968
rect 73599 50934 73620 50968
rect 73560 50920 73620 50934
rect 73140 50820 73200 50880
rect 73140 50710 73200 50770
rect 72720 50658 72780 50670
rect 72720 50624 72748 50658
rect 72748 50624 72780 50658
rect 72720 50610 72780 50624
rect 73140 50540 73200 50600
rect 73560 50658 73620 50670
rect 73560 50624 73565 50658
rect 73565 50624 73599 50658
rect 73599 50624 73620 50658
rect 73560 50610 73620 50624
rect 72720 49258 72780 49270
rect 73140 49280 73200 49340
rect 72720 49224 72748 49258
rect 72748 49224 72780 49258
rect 72720 49210 72780 49224
rect 73560 49258 73620 49270
rect 73560 49224 73565 49258
rect 73565 49224 73599 49258
rect 73599 49224 73620 49258
rect 73560 49210 73620 49224
rect 73140 49110 73200 49170
rect 73140 49000 73200 49060
rect 72720 48948 72780 48960
rect 72720 48914 72748 48948
rect 72748 48914 72780 48948
rect 72720 48900 72780 48914
rect 73140 48830 73200 48890
rect 73560 48948 73620 48960
rect 73560 48914 73565 48948
rect 73565 48914 73599 48948
rect 73599 48914 73620 48948
rect 73560 48900 73620 48914
rect 72720 47548 72780 47560
rect 73140 47570 73200 47630
rect 72720 47514 72748 47548
rect 72748 47514 72780 47548
rect 72720 47500 72780 47514
rect 73560 47548 73620 47560
rect 73560 47514 73565 47548
rect 73565 47514 73599 47548
rect 73599 47514 73620 47548
rect 73560 47500 73620 47514
rect 73140 47400 73200 47460
rect 73140 47290 73200 47350
rect 72720 47238 72780 47250
rect 72720 47204 72748 47238
rect 72748 47204 72780 47238
rect 72720 47190 72780 47204
rect 73140 47120 73200 47180
rect 73560 47238 73620 47250
rect 73560 47204 73565 47238
rect 73565 47204 73599 47238
rect 73599 47204 73620 47238
rect 73560 47190 73620 47204
rect 72720 45838 72780 45850
rect 73140 45860 73200 45920
rect 72720 45804 72748 45838
rect 72748 45804 72780 45838
rect 72720 45790 72780 45804
rect 73560 45838 73620 45850
rect 73560 45804 73565 45838
rect 73565 45804 73599 45838
rect 73599 45804 73620 45838
rect 73560 45790 73620 45804
rect 73140 45690 73200 45750
rect 73140 45580 73200 45640
rect 72720 45528 72780 45540
rect 72720 45494 72748 45528
rect 72748 45494 72780 45528
rect 72720 45480 72780 45494
rect 73140 45410 73200 45470
rect 73560 45528 73620 45540
rect 73560 45494 73565 45528
rect 73565 45494 73599 45528
rect 73599 45494 73620 45528
rect 73560 45480 73620 45494
rect 72720 44128 72780 44140
rect 73140 44150 73200 44210
rect 72720 44094 72748 44128
rect 72748 44094 72780 44128
rect 72720 44080 72780 44094
rect 73560 44128 73620 44140
rect 73560 44094 73565 44128
rect 73565 44094 73599 44128
rect 73599 44094 73620 44128
rect 73560 44080 73620 44094
rect 73140 43980 73200 44040
rect 73140 43870 73200 43930
rect 72720 43818 72780 43830
rect 72720 43784 72748 43818
rect 72748 43784 72780 43818
rect 72720 43770 72780 43784
rect 73140 43700 73200 43760
rect 73560 43818 73620 43830
rect 73560 43784 73565 43818
rect 73565 43784 73599 43818
rect 73599 43784 73620 43818
rect 73560 43770 73620 43784
rect 72720 42418 72780 42430
rect 73140 42440 73200 42500
rect 72720 42384 72748 42418
rect 72748 42384 72780 42418
rect 72720 42370 72780 42384
rect 73560 42418 73620 42430
rect 73560 42384 73565 42418
rect 73565 42384 73599 42418
rect 73599 42384 73620 42418
rect 73560 42370 73620 42384
rect 73140 42270 73200 42330
rect 73140 42160 73200 42220
rect 72720 42108 72780 42120
rect 72720 42074 72748 42108
rect 72748 42074 72780 42108
rect 72720 42060 72780 42074
rect 73140 41990 73200 42050
rect 73560 42108 73620 42120
rect 73560 42074 73565 42108
rect 73565 42074 73599 42108
rect 73599 42074 73620 42108
rect 73560 42060 73620 42074
rect 72720 40708 72780 40720
rect 73140 40730 73200 40790
rect 72720 40674 72748 40708
rect 72748 40674 72780 40708
rect 72720 40660 72780 40674
rect 73560 40708 73620 40720
rect 73560 40674 73565 40708
rect 73565 40674 73599 40708
rect 73599 40674 73620 40708
rect 73560 40660 73620 40674
rect 73140 40560 73200 40620
rect 73140 40450 73200 40510
rect 72720 40398 72780 40410
rect 72720 40364 72748 40398
rect 72748 40364 72780 40398
rect 72720 40350 72780 40364
rect 73140 40280 73200 40340
rect 73560 40398 73620 40410
rect 73560 40364 73565 40398
rect 73565 40364 73599 40398
rect 73599 40364 73620 40398
rect 73560 40350 73620 40364
rect 72610 39620 72670 39680
rect 73680 39620 73740 39680
rect 73780 66410 73840 66470
rect 73840 65880 73900 65940
rect 73780 64700 73840 64760
rect 73840 64170 73900 64230
rect 73780 62990 73840 63050
rect 73840 62460 73900 62520
rect 73780 61280 73840 61340
rect 73840 60750 73900 60810
rect 73780 59570 73840 59630
rect 73840 59040 73900 59100
rect 73780 57860 73840 57920
rect 73840 57330 73900 57390
rect 73780 56150 73840 56210
rect 73840 55620 73900 55680
rect 73780 54440 73840 54500
rect 73840 53910 73900 53970
rect 73780 52730 73840 52790
rect 73840 52200 73900 52260
rect 73780 51020 73840 51080
rect 73840 50490 73900 50550
rect 73780 49310 73840 49370
rect 73840 48780 73900 48840
rect 73780 47600 73840 47660
rect 73840 47070 73900 47130
rect 73780 45890 73840 45950
rect 73840 45360 73900 45420
rect 73780 44180 73840 44240
rect 73840 43650 73900 43710
rect 73780 42470 73840 42530
rect 73840 41940 73900 42000
rect 73780 40760 73840 40820
rect 72310 39170 72370 39230
rect 73840 40230 73900 40290
rect 73840 39620 73900 39680
rect 73930 66320 73990 66380
rect 73930 64610 73990 64670
rect 73930 62900 73990 62960
rect 73930 61190 73990 61250
rect 73930 59480 73990 59540
rect 73930 57770 73990 57830
rect 73930 56060 73990 56120
rect 73930 54350 73990 54410
rect 73930 52640 73990 52700
rect 73930 50930 73990 50990
rect 73930 49220 73990 49280
rect 73930 47510 73990 47570
rect 73930 45800 73990 45860
rect 73930 44090 73990 44150
rect 73930 42380 73990 42440
rect 73930 40670 73990 40730
rect 77500 66320 77560 66380
rect 77500 64610 77560 64670
rect 77500 62900 77560 62960
rect 77500 61190 77560 61250
rect 77500 59480 77560 59540
rect 77500 57770 77560 57830
rect 77500 56060 77560 56120
rect 77500 54350 77560 54410
rect 77500 52640 77560 52700
rect 77500 50930 77560 50990
rect 77500 49220 77560 49280
rect 77500 47510 77560 47570
rect 77500 45800 77560 45860
rect 77500 44090 77560 44150
rect 77500 42380 77560 42440
rect 77500 40670 77560 40730
rect 77710 66358 77770 66370
rect 78130 66380 78190 66440
rect 77710 66324 77738 66358
rect 77738 66324 77770 66358
rect 77710 66310 77770 66324
rect 78550 66358 78610 66370
rect 78550 66324 78555 66358
rect 78555 66324 78589 66358
rect 78589 66324 78610 66358
rect 78550 66310 78610 66324
rect 78130 66210 78190 66270
rect 78130 66100 78190 66160
rect 77710 66048 77770 66060
rect 77710 66014 77738 66048
rect 77738 66014 77770 66048
rect 77710 66000 77770 66014
rect 78130 65930 78190 65990
rect 78550 66048 78610 66060
rect 78550 66014 78555 66048
rect 78555 66014 78589 66048
rect 78589 66014 78610 66048
rect 78550 66000 78610 66014
rect 77710 64648 77770 64660
rect 78130 64670 78190 64730
rect 77710 64614 77738 64648
rect 77738 64614 77770 64648
rect 77710 64600 77770 64614
rect 78550 64648 78610 64660
rect 78550 64614 78555 64648
rect 78555 64614 78589 64648
rect 78589 64614 78610 64648
rect 78550 64600 78610 64614
rect 78130 64500 78190 64560
rect 78130 64390 78190 64450
rect 77710 64338 77770 64350
rect 77710 64304 77738 64338
rect 77738 64304 77770 64338
rect 77710 64290 77770 64304
rect 78130 64220 78190 64280
rect 78550 64338 78610 64350
rect 78550 64304 78555 64338
rect 78555 64304 78589 64338
rect 78589 64304 78610 64338
rect 78550 64290 78610 64304
rect 77710 62938 77770 62950
rect 78130 62960 78190 63020
rect 77710 62904 77738 62938
rect 77738 62904 77770 62938
rect 77710 62890 77770 62904
rect 78550 62938 78610 62950
rect 78550 62904 78555 62938
rect 78555 62904 78589 62938
rect 78589 62904 78610 62938
rect 78550 62890 78610 62904
rect 78130 62790 78190 62850
rect 78130 62680 78190 62740
rect 77710 62628 77770 62640
rect 77710 62594 77738 62628
rect 77738 62594 77770 62628
rect 77710 62580 77770 62594
rect 78130 62510 78190 62570
rect 78550 62628 78610 62640
rect 78550 62594 78555 62628
rect 78555 62594 78589 62628
rect 78589 62594 78610 62628
rect 78550 62580 78610 62594
rect 77710 61228 77770 61240
rect 78130 61250 78190 61310
rect 77710 61194 77738 61228
rect 77738 61194 77770 61228
rect 77710 61180 77770 61194
rect 78550 61228 78610 61240
rect 78550 61194 78555 61228
rect 78555 61194 78589 61228
rect 78589 61194 78610 61228
rect 78550 61180 78610 61194
rect 78130 61080 78190 61140
rect 78130 60970 78190 61030
rect 77710 60918 77770 60930
rect 77710 60884 77738 60918
rect 77738 60884 77770 60918
rect 77710 60870 77770 60884
rect 78130 60800 78190 60860
rect 78550 60918 78610 60930
rect 78550 60884 78555 60918
rect 78555 60884 78589 60918
rect 78589 60884 78610 60918
rect 78550 60870 78610 60884
rect 77710 59518 77770 59530
rect 78130 59540 78190 59600
rect 77710 59484 77738 59518
rect 77738 59484 77770 59518
rect 77710 59470 77770 59484
rect 78550 59518 78610 59530
rect 78550 59484 78555 59518
rect 78555 59484 78589 59518
rect 78589 59484 78610 59518
rect 78550 59470 78610 59484
rect 78130 59370 78190 59430
rect 78130 59260 78190 59320
rect 77710 59208 77770 59220
rect 77710 59174 77738 59208
rect 77738 59174 77770 59208
rect 77710 59160 77770 59174
rect 78130 59090 78190 59150
rect 78550 59208 78610 59220
rect 78550 59174 78555 59208
rect 78555 59174 78589 59208
rect 78589 59174 78610 59208
rect 78550 59160 78610 59174
rect 77710 57808 77770 57820
rect 78130 57830 78190 57890
rect 77710 57774 77738 57808
rect 77738 57774 77770 57808
rect 77710 57760 77770 57774
rect 78550 57808 78610 57820
rect 78550 57774 78555 57808
rect 78555 57774 78589 57808
rect 78589 57774 78610 57808
rect 78550 57760 78610 57774
rect 78130 57660 78190 57720
rect 78130 57550 78190 57610
rect 77710 57498 77770 57510
rect 77710 57464 77738 57498
rect 77738 57464 77770 57498
rect 77710 57450 77770 57464
rect 78130 57380 78190 57440
rect 78550 57498 78610 57510
rect 78550 57464 78555 57498
rect 78555 57464 78589 57498
rect 78589 57464 78610 57498
rect 78550 57450 78610 57464
rect 77710 56098 77770 56110
rect 78130 56120 78190 56180
rect 77710 56064 77738 56098
rect 77738 56064 77770 56098
rect 77710 56050 77770 56064
rect 78550 56098 78610 56110
rect 78550 56064 78555 56098
rect 78555 56064 78589 56098
rect 78589 56064 78610 56098
rect 78550 56050 78610 56064
rect 78130 55950 78190 56010
rect 78130 55840 78190 55900
rect 77710 55788 77770 55800
rect 77710 55754 77738 55788
rect 77738 55754 77770 55788
rect 77710 55740 77770 55754
rect 78130 55670 78190 55730
rect 78550 55788 78610 55800
rect 78550 55754 78555 55788
rect 78555 55754 78589 55788
rect 78589 55754 78610 55788
rect 78550 55740 78610 55754
rect 77710 54388 77770 54400
rect 78130 54410 78190 54470
rect 77710 54354 77738 54388
rect 77738 54354 77770 54388
rect 77710 54340 77770 54354
rect 78550 54388 78610 54400
rect 78550 54354 78555 54388
rect 78555 54354 78589 54388
rect 78589 54354 78610 54388
rect 78550 54340 78610 54354
rect 78130 54240 78190 54300
rect 78130 54130 78190 54190
rect 77710 54078 77770 54090
rect 77710 54044 77738 54078
rect 77738 54044 77770 54078
rect 77710 54030 77770 54044
rect 78130 53960 78190 54020
rect 78550 54078 78610 54090
rect 78550 54044 78555 54078
rect 78555 54044 78589 54078
rect 78589 54044 78610 54078
rect 78550 54030 78610 54044
rect 77710 52678 77770 52690
rect 78130 52700 78190 52760
rect 77710 52644 77738 52678
rect 77738 52644 77770 52678
rect 77710 52630 77770 52644
rect 78550 52678 78610 52690
rect 78550 52644 78555 52678
rect 78555 52644 78589 52678
rect 78589 52644 78610 52678
rect 78550 52630 78610 52644
rect 78130 52530 78190 52590
rect 78130 52420 78190 52480
rect 77710 52368 77770 52380
rect 77710 52334 77738 52368
rect 77738 52334 77770 52368
rect 77710 52320 77770 52334
rect 78130 52250 78190 52310
rect 78550 52368 78610 52380
rect 78550 52334 78555 52368
rect 78555 52334 78589 52368
rect 78589 52334 78610 52368
rect 78550 52320 78610 52334
rect 77710 50968 77770 50980
rect 78130 50990 78190 51050
rect 77710 50934 77738 50968
rect 77738 50934 77770 50968
rect 77710 50920 77770 50934
rect 78550 50968 78610 50980
rect 78550 50934 78555 50968
rect 78555 50934 78589 50968
rect 78589 50934 78610 50968
rect 78550 50920 78610 50934
rect 78130 50820 78190 50880
rect 78130 50710 78190 50770
rect 77710 50658 77770 50670
rect 77710 50624 77738 50658
rect 77738 50624 77770 50658
rect 77710 50610 77770 50624
rect 78130 50540 78190 50600
rect 78550 50658 78610 50670
rect 78550 50624 78555 50658
rect 78555 50624 78589 50658
rect 78589 50624 78610 50658
rect 78550 50610 78610 50624
rect 77710 49258 77770 49270
rect 78130 49280 78190 49340
rect 77710 49224 77738 49258
rect 77738 49224 77770 49258
rect 77710 49210 77770 49224
rect 78550 49258 78610 49270
rect 78550 49224 78555 49258
rect 78555 49224 78589 49258
rect 78589 49224 78610 49258
rect 78550 49210 78610 49224
rect 78130 49110 78190 49170
rect 78130 49000 78190 49060
rect 77710 48948 77770 48960
rect 77710 48914 77738 48948
rect 77738 48914 77770 48948
rect 77710 48900 77770 48914
rect 78130 48830 78190 48890
rect 78550 48948 78610 48960
rect 78550 48914 78555 48948
rect 78555 48914 78589 48948
rect 78589 48914 78610 48948
rect 78550 48900 78610 48914
rect 77710 47548 77770 47560
rect 78130 47570 78190 47630
rect 77710 47514 77738 47548
rect 77738 47514 77770 47548
rect 77710 47500 77770 47514
rect 78550 47548 78610 47560
rect 78550 47514 78555 47548
rect 78555 47514 78589 47548
rect 78589 47514 78610 47548
rect 78550 47500 78610 47514
rect 78130 47400 78190 47460
rect 78130 47290 78190 47350
rect 77710 47238 77770 47250
rect 77710 47204 77738 47238
rect 77738 47204 77770 47238
rect 77710 47190 77770 47204
rect 78130 47120 78190 47180
rect 78550 47238 78610 47250
rect 78550 47204 78555 47238
rect 78555 47204 78589 47238
rect 78589 47204 78610 47238
rect 78550 47190 78610 47204
rect 77710 45838 77770 45850
rect 78130 45860 78190 45920
rect 77710 45804 77738 45838
rect 77738 45804 77770 45838
rect 77710 45790 77770 45804
rect 78550 45838 78610 45850
rect 78550 45804 78555 45838
rect 78555 45804 78589 45838
rect 78589 45804 78610 45838
rect 78550 45790 78610 45804
rect 78130 45690 78190 45750
rect 78130 45580 78190 45640
rect 77710 45528 77770 45540
rect 77710 45494 77738 45528
rect 77738 45494 77770 45528
rect 77710 45480 77770 45494
rect 78130 45410 78190 45470
rect 78550 45528 78610 45540
rect 78550 45494 78555 45528
rect 78555 45494 78589 45528
rect 78589 45494 78610 45528
rect 78550 45480 78610 45494
rect 77710 44128 77770 44140
rect 78130 44150 78190 44210
rect 77710 44094 77738 44128
rect 77738 44094 77770 44128
rect 77710 44080 77770 44094
rect 78550 44128 78610 44140
rect 78550 44094 78555 44128
rect 78555 44094 78589 44128
rect 78589 44094 78610 44128
rect 78550 44080 78610 44094
rect 78130 43980 78190 44040
rect 78130 43870 78190 43930
rect 77710 43818 77770 43830
rect 77710 43784 77738 43818
rect 77738 43784 77770 43818
rect 77710 43770 77770 43784
rect 78130 43700 78190 43760
rect 78550 43818 78610 43830
rect 78550 43784 78555 43818
rect 78555 43784 78589 43818
rect 78589 43784 78610 43818
rect 78550 43770 78610 43784
rect 77710 42418 77770 42430
rect 78130 42440 78190 42500
rect 77710 42384 77738 42418
rect 77738 42384 77770 42418
rect 77710 42370 77770 42384
rect 78550 42418 78610 42430
rect 78550 42384 78555 42418
rect 78555 42384 78589 42418
rect 78589 42384 78610 42418
rect 78550 42370 78610 42384
rect 78130 42270 78190 42330
rect 78130 42160 78190 42220
rect 77710 42108 77770 42120
rect 77710 42074 77738 42108
rect 77738 42074 77770 42108
rect 77710 42060 77770 42074
rect 78130 41990 78190 42050
rect 78550 42108 78610 42120
rect 78550 42074 78555 42108
rect 78555 42074 78589 42108
rect 78589 42074 78610 42108
rect 78550 42060 78610 42074
rect 77710 40708 77770 40720
rect 78130 40730 78190 40790
rect 77710 40674 77738 40708
rect 77738 40674 77770 40708
rect 77710 40660 77770 40674
rect 78550 40708 78610 40720
rect 78550 40674 78555 40708
rect 78555 40674 78589 40708
rect 78589 40674 78610 40708
rect 78550 40660 78610 40674
rect 78130 40560 78190 40620
rect 78130 40450 78190 40510
rect 77710 40398 77770 40410
rect 77710 40364 77738 40398
rect 77738 40364 77770 40398
rect 77710 40350 77770 40364
rect 78130 40280 78190 40340
rect 78550 40398 78610 40410
rect 78550 40364 78555 40398
rect 78555 40364 78589 40398
rect 78589 40364 78610 40398
rect 78550 40350 78610 40364
rect 77600 39620 77660 39680
rect 78670 39620 78730 39680
rect 78770 66410 78830 66470
rect 78830 65880 78890 65940
rect 78770 64700 78830 64760
rect 78830 64170 78890 64230
rect 78770 62990 78830 63050
rect 78830 62460 78890 62520
rect 78770 61280 78830 61340
rect 78830 60750 78890 60810
rect 78770 59570 78830 59630
rect 78830 59040 78890 59100
rect 78770 57860 78830 57920
rect 78830 57330 78890 57390
rect 78770 56150 78830 56210
rect 78830 55620 78890 55680
rect 78770 54440 78830 54500
rect 78830 53910 78890 53970
rect 78770 52730 78830 52790
rect 78830 52200 78890 52260
rect 78770 51020 78830 51080
rect 78830 50490 78890 50550
rect 78770 49310 78830 49370
rect 78830 48780 78890 48840
rect 78770 47600 78830 47660
rect 78830 47070 78890 47130
rect 78770 45890 78830 45950
rect 78830 45360 78890 45420
rect 78770 44180 78830 44240
rect 78830 43650 78890 43710
rect 78770 42470 78830 42530
rect 78830 41940 78890 42000
rect 78770 40760 78830 40820
rect 74130 39170 74190 39230
rect 77300 39170 77360 39230
rect 78830 40230 78890 40290
rect 78830 39620 78890 39680
rect 78920 66320 78980 66380
rect 78920 64610 78980 64670
rect 78920 62900 78980 62960
rect 78920 61190 78980 61250
rect 78920 59480 78980 59540
rect 78920 57770 78980 57830
rect 78920 56060 78980 56120
rect 78920 54350 78980 54410
rect 78920 52640 78980 52700
rect 78920 50930 78980 50990
rect 78920 49220 78980 49280
rect 78920 47510 78980 47570
rect 78920 45800 78980 45860
rect 78920 44090 78980 44150
rect 78920 42380 78980 42440
rect 78920 40670 78980 40730
rect 79120 39170 79180 39230
rect 3970 38640 4030 38700
rect 8960 38640 9020 38700
rect 13950 38640 14010 38700
rect 18940 38640 19000 38700
rect 23930 38640 23990 38700
rect 28920 38640 28980 38700
rect 33910 38640 33970 38700
rect 38900 38640 38960 38700
rect 43890 38640 43950 38700
rect 48880 38640 48940 38700
rect 53870 38640 53930 38700
rect 58860 38640 58920 38700
rect 63850 38640 63910 38700
rect 68840 38640 68900 38700
rect 73830 38640 73890 38700
rect 78820 38640 78880 38700
rect 40200 38500 40260 38560
rect 40270 38360 40330 38420
rect 45020 38220 45080 38280
rect 45110 38080 45170 38140
rect 40030 37940 40090 38000
rect 45200 37940 45260 38000
rect 40090 37800 40150 37860
rect 45260 37800 45320 37860
rect 34860 37660 34920 37720
rect 49830 37660 49890 37720
rect 34920 37520 34980 37580
rect 49890 37520 49950 37580
rect 35040 37380 35100 37440
rect 39850 37380 39910 37440
rect 44840 37380 44900 37440
rect 50010 37380 50070 37440
rect 35100 37240 35160 37300
rect 39910 37240 39970 37300
rect 44900 37240 44960 37300
rect 50070 37240 50130 37300
rect 24520 37100 24580 37160
rect 29510 37100 29570 37160
rect 34680 37100 34740 37160
rect 39670 37100 39730 37160
rect 44660 37100 44720 37160
rect 49650 37100 49710 37160
rect 54460 37100 54520 37160
rect 59450 37100 59510 37160
rect 24580 36960 24640 37020
rect 29570 36960 29630 37020
rect 34740 36960 34800 37020
rect 39730 36960 39790 37020
rect 44720 36960 44780 37020
rect 49710 36960 49770 37020
rect 54520 36960 54580 37020
rect 59510 36960 59570 37020
rect 24700 36820 24760 36880
rect 29690 36820 29750 36880
rect 34500 36820 34560 36880
rect 39490 36820 39550 36880
rect 44480 36820 44540 36880
rect 49470 36820 49530 36880
rect 54640 36820 54700 36880
rect 59630 36820 59690 36880
rect 24760 36680 24820 36740
rect 29750 36680 29810 36740
rect 34560 36680 34620 36740
rect 39550 36680 39610 36740
rect 44540 36680 44600 36740
rect 49530 36680 49590 36740
rect 54700 36680 54760 36740
rect 59690 36680 59750 36740
rect 14360 36540 14420 36600
rect 19350 36540 19410 36600
rect 24340 36540 24400 36600
rect 29330 36540 29390 36600
rect 34320 36540 34380 36600
rect 39310 36540 39370 36600
rect 44300 36540 44360 36600
rect 49290 36540 49350 36600
rect 54280 36540 54340 36600
rect 59270 36540 59330 36600
rect 64260 36540 64320 36600
rect 69250 36540 69310 36600
rect 14420 36400 14480 36460
rect 19410 36400 19470 36460
rect 24400 36400 24460 36460
rect 29390 36400 29450 36460
rect 34380 36400 34440 36460
rect 39370 36400 39430 36460
rect 44360 36400 44420 36460
rect 49350 36400 49410 36460
rect 54340 36400 54400 36460
rect 59330 36400 59390 36460
rect 64320 36400 64380 36460
rect 69310 36400 69370 36460
rect 4200 36260 4260 36320
rect 9190 36260 9250 36320
rect 14180 36260 14240 36320
rect 19170 36260 19230 36320
rect 24160 36260 24220 36320
rect 29150 36260 29210 36320
rect 34140 36260 34200 36320
rect 39130 36260 39190 36320
rect 44120 36260 44180 36320
rect 49110 36260 49170 36320
rect 54100 36260 54160 36320
rect 59090 36260 59150 36320
rect 64080 36260 64140 36320
rect 69070 36260 69130 36320
rect 74060 36260 74120 36320
rect 79050 36260 79110 36320
rect 4260 36120 4320 36180
rect 9250 36120 9310 36180
rect 14240 36120 14300 36180
rect 19230 36120 19290 36180
rect 24220 36120 24280 36180
rect 29210 36120 29270 36180
rect 34200 36120 34260 36180
rect 39190 36120 39250 36180
rect 44180 36120 44240 36180
rect 49170 36120 49230 36180
rect 54160 36120 54220 36180
rect 59150 36120 59210 36180
rect 64140 36120 64200 36180
rect 69130 36120 69190 36180
rect 74120 36120 74180 36180
rect 79110 36120 79170 36180
rect 4160 30870 4220 30930
rect 9150 30870 9210 30930
rect 14140 30870 14200 30930
rect 19130 30870 19190 30930
rect 24120 30870 24180 30930
rect 29110 30870 29170 30930
rect 34100 30870 34160 30930
rect 39090 30870 39150 30930
rect 44080 30870 44140 30930
rect 49070 30870 49130 30930
rect 54060 30870 54120 30930
rect 59050 30870 59110 30930
rect 64040 30870 64100 30930
rect 69030 30870 69090 30930
rect 74020 30870 74080 30930
rect 79010 30870 79070 30930
rect 4100 30730 4160 30790
rect 9090 30730 9150 30790
rect 14080 30730 14140 30790
rect 19070 30730 19130 30790
rect 24060 30730 24120 30790
rect 29050 30730 29110 30790
rect 34040 30730 34100 30790
rect 39030 30730 39090 30790
rect 44020 30730 44080 30790
rect 49010 30730 49070 30790
rect 54000 30730 54060 30790
rect 58990 30730 59050 30790
rect 63980 30730 64040 30790
rect 68970 30730 69030 30790
rect 73960 30730 74020 30790
rect 78950 30730 79010 30790
rect 14320 30590 14380 30650
rect 19310 30590 19370 30650
rect 24300 30590 24360 30650
rect 29290 30590 29350 30650
rect 34280 30590 34340 30650
rect 39270 30590 39330 30650
rect 44260 30590 44320 30650
rect 49250 30590 49310 30650
rect 54240 30590 54300 30650
rect 59230 30590 59290 30650
rect 64220 30590 64280 30650
rect 69210 30590 69270 30650
rect 14260 30450 14320 30510
rect 19250 30450 19310 30510
rect 24240 30450 24300 30510
rect 29230 30450 29290 30510
rect 34220 30450 34280 30510
rect 39210 30450 39270 30510
rect 44200 30450 44260 30510
rect 49190 30450 49250 30510
rect 54180 30450 54240 30510
rect 59170 30450 59230 30510
rect 64160 30450 64220 30510
rect 69150 30450 69210 30510
rect 24660 30310 24720 30370
rect 29650 30310 29710 30370
rect 34460 30310 34520 30370
rect 39450 30310 39510 30370
rect 44440 30310 44500 30370
rect 49430 30310 49490 30370
rect 54600 30310 54660 30370
rect 59590 30310 59650 30370
rect 24600 30170 24660 30230
rect 29590 30170 29650 30230
rect 34400 30170 34460 30230
rect 39390 30170 39450 30230
rect 44380 30170 44440 30230
rect 49370 30170 49430 30230
rect 54540 30170 54600 30230
rect 59530 30170 59590 30230
rect 24480 30030 24540 30090
rect 29470 30030 29530 30090
rect 34640 30030 34700 30090
rect 39630 30030 39690 30090
rect 44620 30030 44680 30090
rect 49610 30030 49670 30090
rect 54420 30030 54480 30090
rect 59410 30030 59470 30090
rect 24420 29890 24480 29950
rect 29410 29890 29470 29950
rect 34580 29890 34640 29950
rect 39570 29890 39630 29950
rect 44560 29890 44620 29950
rect 49550 29890 49610 29950
rect 54360 29890 54420 29950
rect 59350 29890 59410 29950
rect 35000 29750 35060 29810
rect 39810 29750 39870 29810
rect 44800 29750 44860 29810
rect 49970 29750 50030 29810
rect 34940 29610 35000 29670
rect 39750 29610 39810 29670
rect 44740 29610 44800 29670
rect 49910 29610 49970 29670
rect 34820 29470 34880 29530
rect 49790 29470 49850 29530
rect 34760 29330 34820 29390
rect 49730 29330 49790 29390
rect 39990 29190 40050 29250
rect 45160 29190 45220 29250
rect 39930 29050 39990 29110
rect 45100 29050 45160 29110
rect 45010 28910 45070 28970
rect 44920 28770 44980 28830
rect 40170 28630 40230 28690
rect 40100 28490 40160 28550
rect 3870 28350 3930 28410
rect 8860 28350 8920 28410
rect 13850 28350 13910 28410
rect 18840 28350 18900 28410
rect 23830 28350 23890 28410
rect 28820 28350 28880 28410
rect 33810 28350 33870 28410
rect 38800 28350 38860 28410
rect 43790 28350 43850 28410
rect 48780 28350 48840 28410
rect 53770 28350 53830 28410
rect 58760 28350 58820 28410
rect 63750 28350 63810 28410
rect 68740 28350 68800 28410
rect 73730 28350 73790 28410
rect 78720 28350 78780 28410
rect 2350 27820 2410 27880
rect 2650 27370 2710 27430
rect 3720 27370 3780 27430
rect 4170 27820 4230 27880
rect 7340 27820 7400 27880
rect 3880 27370 3940 27430
rect 7640 27370 7700 27430
rect 8710 27370 8770 27430
rect 9160 27820 9220 27880
rect 8870 27370 8930 27430
rect 12150 27760 12210 27820
rect 12330 27820 12390 27880
rect 12630 27370 12690 27430
rect 13700 27370 13760 27430
rect 14150 27820 14210 27880
rect 13860 27370 13920 27430
rect 14330 27760 14390 27820
rect 17140 27760 17200 27820
rect 17320 27820 17380 27880
rect 17620 27370 17680 27430
rect 18690 27370 18750 27430
rect 19140 27820 19200 27880
rect 18850 27370 18910 27430
rect 19320 27760 19380 27820
rect 21770 27640 21830 27700
rect 21950 27700 22010 27760
rect 22130 27760 22190 27820
rect 22310 27820 22370 27880
rect 22610 27370 22670 27430
rect 23680 27370 23740 27430
rect 24130 27820 24190 27880
rect 23840 27370 23900 27430
rect 24310 27760 24370 27820
rect 24490 27700 24550 27760
rect 24670 27640 24730 27700
rect 26760 27640 26820 27700
rect 26940 27700 27000 27760
rect 27120 27760 27180 27820
rect 27300 27820 27360 27880
rect 27600 27370 27660 27430
rect 28670 27370 28730 27430
rect 29120 27820 29180 27880
rect 28830 27370 28890 27430
rect 29300 27760 29360 27820
rect 29480 27700 29540 27760
rect 29660 27640 29720 27700
rect 31390 27520 31450 27580
rect 31570 27580 31630 27640
rect 31750 27640 31810 27700
rect 31930 27700 31990 27760
rect 32110 27760 32170 27820
rect 32290 27820 32350 27880
rect 32590 27370 32650 27430
rect 33660 27370 33720 27430
rect 34110 27820 34170 27880
rect 33820 27370 33880 27430
rect 34290 27760 34350 27820
rect 34470 27700 34530 27760
rect 34650 27640 34710 27700
rect 34830 27580 34890 27640
rect 35010 27520 35070 27580
rect 36200 27460 36260 27520
rect 36380 27520 36440 27580
rect 36560 27580 36620 27640
rect 36740 27640 36800 27700
rect 36920 27700 36980 27760
rect 37100 27760 37160 27820
rect 37280 27820 37340 27880
rect 37580 27370 37640 27430
rect 38650 27370 38710 27430
rect 39100 27820 39160 27880
rect 38810 27370 38870 27430
rect 39280 27760 39340 27820
rect 39460 27700 39520 27760
rect 39640 27640 39700 27700
rect 39820 27580 39880 27640
rect 40000 27520 40060 27580
rect 40180 27460 40240 27520
rect 41190 27460 41250 27520
rect 41370 27520 41430 27580
rect 41550 27580 41610 27640
rect 41730 27640 41790 27700
rect 41910 27700 41970 27760
rect 42090 27760 42150 27820
rect 42270 27820 42330 27880
rect 42570 27370 42630 27430
rect 43640 27370 43700 27430
rect 44090 27820 44150 27880
rect 43800 27370 43860 27430
rect 44270 27760 44330 27820
rect 44450 27700 44510 27760
rect 44630 27640 44690 27700
rect 44810 27580 44870 27640
rect 44990 27520 45050 27580
rect 45170 27460 45230 27520
rect 46360 27520 46420 27580
rect 46540 27580 46600 27640
rect 46720 27640 46780 27700
rect 46900 27700 46960 27760
rect 47080 27760 47140 27820
rect 47260 27820 47320 27880
rect 47560 27370 47620 27430
rect 48630 27370 48690 27430
rect 49080 27820 49140 27880
rect 48790 27370 48850 27430
rect 49260 27760 49320 27820
rect 49440 27700 49500 27760
rect 49620 27640 49680 27700
rect 49800 27580 49860 27640
rect 51710 27640 51770 27700
rect 51890 27700 51950 27760
rect 52070 27760 52130 27820
rect 52250 27820 52310 27880
rect 49980 27520 50040 27580
rect 52550 27370 52610 27430
rect 53620 27370 53680 27430
rect 54070 27820 54130 27880
rect 53780 27370 53840 27430
rect 54250 27760 54310 27820
rect 54430 27700 54490 27760
rect 54610 27640 54670 27700
rect 56700 27640 56760 27700
rect 56880 27700 56940 27760
rect 57060 27760 57120 27820
rect 57240 27820 57300 27880
rect 57540 27370 57600 27430
rect 58610 27370 58670 27430
rect 59060 27820 59120 27880
rect 58770 27370 58830 27430
rect 59240 27760 59300 27820
rect 59420 27700 59480 27760
rect 62050 27760 62110 27820
rect 62230 27820 62290 27880
rect 59600 27640 59660 27700
rect 62530 27370 62590 27430
rect 63600 27370 63660 27430
rect 64050 27820 64110 27880
rect 63760 27370 63820 27430
rect 64230 27760 64290 27820
rect 67040 27760 67100 27820
rect 67220 27820 67280 27880
rect 67520 27370 67580 27430
rect 68590 27370 68650 27430
rect 69040 27820 69100 27880
rect 68750 27370 68810 27430
rect 69220 27760 69280 27820
rect 72210 27820 72270 27880
rect 72510 27370 72570 27430
rect 73580 27370 73640 27430
rect 74030 27820 74090 27880
rect 77200 27820 77260 27880
rect 73740 27370 73800 27430
rect 77500 27370 77560 27430
rect 78570 27370 78630 27430
rect 79020 27820 79080 27880
rect 78730 27370 78790 27430
<< metal2 >>
rect 2680 66590 2710 67050
rect 2630 66580 2710 66590
rect 2630 66520 2640 66580
rect 2700 66520 2710 66580
rect 2630 66510 2710 66520
rect 4070 66590 4100 67050
rect 7670 66590 7700 67050
rect 4070 66580 4150 66590
rect 4070 66520 4080 66580
rect 4140 66520 4150 66580
rect 4070 66510 4150 66520
rect 7620 66580 7700 66590
rect 7620 66520 7630 66580
rect 7690 66520 7700 66580
rect 7620 66510 7700 66520
rect 9060 66590 9090 67050
rect 9060 66580 9140 66590
rect 9060 66520 9070 66580
rect 9130 66520 9140 66580
rect 9060 66510 9140 66520
rect 3920 66470 3980 66480
rect 3270 66440 3920 66450
rect 2650 66380 2710 66390
rect 3270 66380 3280 66440
rect 3340 66420 3920 66440
rect 3340 66380 3350 66420
rect 8910 66470 8970 66480
rect 3920 66400 3980 66410
rect 8260 66440 8910 66450
rect 4070 66380 4130 66390
rect 2850 66370 2930 66380
rect 3270 66370 3350 66380
rect 3690 66370 3770 66380
rect 2850 66360 2860 66370
rect 2710 66330 2860 66360
rect 2650 66310 2710 66320
rect 2850 66310 2860 66330
rect 2920 66310 2930 66370
rect 2850 66300 2930 66310
rect 3690 66310 3700 66370
rect 3760 66360 3770 66370
rect 3760 66330 4070 66360
rect 3760 66310 3770 66330
rect 4070 66310 4130 66320
rect 7640 66380 7700 66390
rect 8260 66380 8270 66440
rect 8330 66420 8910 66440
rect 8330 66380 8340 66420
rect 8910 66400 8970 66410
rect 9060 66380 9120 66390
rect 7840 66370 7920 66380
rect 8260 66370 8340 66380
rect 8680 66370 8760 66380
rect 7840 66360 7850 66370
rect 7700 66330 7850 66360
rect 7640 66310 7700 66320
rect 7840 66310 7850 66330
rect 7910 66310 7920 66370
rect 3690 66300 3770 66310
rect 7840 66300 7920 66310
rect 8680 66310 8690 66370
rect 8750 66360 8760 66370
rect 8750 66330 9060 66360
rect 8750 66310 8760 66330
rect 9060 66310 9120 66320
rect 8680 66300 8760 66310
rect 3260 66280 3360 66290
rect 3260 66210 3280 66280
rect 3350 66210 3360 66280
rect 3260 66170 3360 66210
rect 3260 66100 3280 66170
rect 3350 66100 3360 66170
rect 3260 66080 3360 66100
rect 8250 66280 8350 66290
rect 8250 66210 8270 66280
rect 8340 66210 8350 66280
rect 8250 66170 8350 66210
rect 8250 66100 8270 66170
rect 8340 66100 8350 66170
rect 8250 66080 8350 66100
rect 2630 66060 2710 66070
rect 2630 66000 2640 66060
rect 2700 66050 2710 66060
rect 2850 66060 2930 66070
rect 2850 66050 2860 66060
rect 2700 66020 2860 66050
rect 2700 66000 2710 66020
rect 2630 65990 2710 66000
rect 2850 66000 2860 66020
rect 2920 66000 2930 66060
rect 3690 66060 3770 66070
rect 3690 66000 3700 66060
rect 3760 66050 3770 66060
rect 4070 66060 4150 66070
rect 4070 66050 4080 66060
rect 3760 66020 4080 66050
rect 3760 66000 3770 66020
rect 2850 65990 2930 66000
rect 3270 65990 3350 66000
rect 3690 65990 3770 66000
rect 4070 66000 4080 66020
rect 4140 66000 4150 66060
rect 4070 65990 4150 66000
rect 7620 66060 7700 66070
rect 7620 66000 7630 66060
rect 7690 66050 7700 66060
rect 7840 66060 7920 66070
rect 7840 66050 7850 66060
rect 7690 66020 7850 66050
rect 7690 66000 7700 66020
rect 7620 65990 7700 66000
rect 7840 66000 7850 66020
rect 7910 66000 7920 66060
rect 8680 66060 8760 66070
rect 8680 66000 8690 66060
rect 8750 66050 8760 66060
rect 9060 66060 9140 66070
rect 9060 66050 9070 66060
rect 8750 66020 9070 66050
rect 8750 66000 8760 66020
rect 7840 65990 7920 66000
rect 8260 65990 8340 66000
rect 8680 65990 8760 66000
rect 9060 66000 9070 66020
rect 9130 66000 9140 66060
rect 9060 65990 9140 66000
rect 3270 65930 3280 65990
rect 3340 65950 3350 65990
rect 3340 65940 4040 65950
rect 3340 65930 3980 65940
rect 3270 65920 3980 65930
rect 8260 65930 8270 65990
rect 8330 65950 8340 65990
rect 8330 65940 9030 65950
rect 8330 65930 8970 65940
rect 8260 65920 8970 65930
rect 3980 65870 4040 65880
rect 8970 65870 9030 65880
rect 3920 64760 3980 64770
rect 3270 64730 3920 64740
rect 2650 64670 2710 64680
rect 3270 64670 3280 64730
rect 3340 64710 3920 64730
rect 3340 64670 3350 64710
rect 8910 64760 8970 64770
rect 3920 64690 3980 64700
rect 8260 64730 8910 64740
rect 4070 64670 4130 64680
rect 2850 64660 2930 64670
rect 3270 64660 3350 64670
rect 3690 64660 3770 64670
rect 2850 64650 2860 64660
rect 2710 64620 2860 64650
rect 2650 64600 2710 64610
rect 2850 64600 2860 64620
rect 2920 64600 2930 64660
rect 2850 64590 2930 64600
rect 3690 64600 3700 64660
rect 3760 64650 3770 64660
rect 3760 64620 4070 64650
rect 3760 64600 3770 64620
rect 4070 64600 4130 64610
rect 7640 64670 7700 64680
rect 8260 64670 8270 64730
rect 8330 64710 8910 64730
rect 8330 64670 8340 64710
rect 8910 64690 8970 64700
rect 9060 64670 9120 64680
rect 7840 64660 7920 64670
rect 8260 64660 8340 64670
rect 8680 64660 8760 64670
rect 7840 64650 7850 64660
rect 7700 64620 7850 64650
rect 7640 64600 7700 64610
rect 7840 64600 7850 64620
rect 7910 64600 7920 64660
rect 3690 64590 3770 64600
rect 7840 64590 7920 64600
rect 8680 64600 8690 64660
rect 8750 64650 8760 64660
rect 8750 64620 9060 64650
rect 8750 64600 8760 64620
rect 9060 64600 9120 64610
rect 8680 64590 8760 64600
rect 3260 64570 3360 64580
rect 3260 64500 3280 64570
rect 3350 64500 3360 64570
rect 3260 64460 3360 64500
rect 3260 64390 3280 64460
rect 3350 64390 3360 64460
rect 3260 64370 3360 64390
rect 8250 64570 8350 64580
rect 8250 64500 8270 64570
rect 8340 64500 8350 64570
rect 8250 64460 8350 64500
rect 8250 64390 8270 64460
rect 8340 64390 8350 64460
rect 8250 64370 8350 64390
rect 2630 64350 2710 64360
rect 2630 64290 2640 64350
rect 2700 64340 2710 64350
rect 2850 64350 2930 64360
rect 2850 64340 2860 64350
rect 2700 64310 2860 64340
rect 2700 64290 2710 64310
rect 2630 64280 2710 64290
rect 2850 64290 2860 64310
rect 2920 64290 2930 64350
rect 3690 64350 3770 64360
rect 3690 64290 3700 64350
rect 3760 64340 3770 64350
rect 4070 64350 4150 64360
rect 4070 64340 4080 64350
rect 3760 64310 4080 64340
rect 3760 64290 3770 64310
rect 2850 64280 2930 64290
rect 3270 64280 3350 64290
rect 3690 64280 3770 64290
rect 4070 64290 4080 64310
rect 4140 64290 4150 64350
rect 4070 64280 4150 64290
rect 7620 64350 7700 64360
rect 7620 64290 7630 64350
rect 7690 64340 7700 64350
rect 7840 64350 7920 64360
rect 7840 64340 7850 64350
rect 7690 64310 7850 64340
rect 7690 64290 7700 64310
rect 7620 64280 7700 64290
rect 7840 64290 7850 64310
rect 7910 64290 7920 64350
rect 8680 64350 8760 64360
rect 8680 64290 8690 64350
rect 8750 64340 8760 64350
rect 9060 64350 9140 64360
rect 9060 64340 9070 64350
rect 8750 64310 9070 64340
rect 8750 64290 8760 64310
rect 7840 64280 7920 64290
rect 8260 64280 8340 64290
rect 8680 64280 8760 64290
rect 9060 64290 9070 64310
rect 9130 64290 9140 64350
rect 9060 64280 9140 64290
rect 3270 64220 3280 64280
rect 3340 64240 3350 64280
rect 3340 64230 4040 64240
rect 3340 64220 3980 64230
rect 3270 64210 3980 64220
rect 8260 64220 8270 64280
rect 8330 64240 8340 64280
rect 8330 64230 9030 64240
rect 8330 64220 8970 64230
rect 8260 64210 8970 64220
rect 3980 64160 4040 64170
rect 8970 64160 9030 64170
rect 3920 63050 3980 63060
rect 3270 63020 3920 63030
rect 2650 62960 2710 62970
rect 3270 62960 3280 63020
rect 3340 63000 3920 63020
rect 3340 62960 3350 63000
rect 8910 63050 8970 63060
rect 3920 62980 3980 62990
rect 8260 63020 8910 63030
rect 4070 62960 4130 62970
rect 2850 62950 2930 62960
rect 3270 62950 3350 62960
rect 3690 62950 3770 62960
rect 2850 62940 2860 62950
rect 2710 62910 2860 62940
rect 2650 62890 2710 62900
rect 2850 62890 2860 62910
rect 2920 62890 2930 62950
rect 2850 62880 2930 62890
rect 3690 62890 3700 62950
rect 3760 62940 3770 62950
rect 3760 62910 4070 62940
rect 3760 62890 3770 62910
rect 4070 62890 4130 62900
rect 7640 62960 7700 62970
rect 8260 62960 8270 63020
rect 8330 63000 8910 63020
rect 8330 62960 8340 63000
rect 8910 62980 8970 62990
rect 9060 62960 9120 62970
rect 7840 62950 7920 62960
rect 8260 62950 8340 62960
rect 8680 62950 8760 62960
rect 7840 62940 7850 62950
rect 7700 62910 7850 62940
rect 7640 62890 7700 62900
rect 7840 62890 7850 62910
rect 7910 62890 7920 62950
rect 3690 62880 3770 62890
rect 7840 62880 7920 62890
rect 8680 62890 8690 62950
rect 8750 62940 8760 62950
rect 8750 62910 9060 62940
rect 8750 62890 8760 62910
rect 9060 62890 9120 62900
rect 8680 62880 8760 62890
rect 3260 62860 3360 62870
rect 3260 62790 3280 62860
rect 3350 62790 3360 62860
rect 3260 62750 3360 62790
rect 3260 62680 3280 62750
rect 3350 62680 3360 62750
rect 3260 62660 3360 62680
rect 8250 62860 8350 62870
rect 8250 62790 8270 62860
rect 8340 62790 8350 62860
rect 8250 62750 8350 62790
rect 8250 62680 8270 62750
rect 8340 62680 8350 62750
rect 8250 62660 8350 62680
rect 2630 62640 2710 62650
rect 2630 62580 2640 62640
rect 2700 62630 2710 62640
rect 2850 62640 2930 62650
rect 2850 62630 2860 62640
rect 2700 62600 2860 62630
rect 2700 62580 2710 62600
rect 2630 62570 2710 62580
rect 2850 62580 2860 62600
rect 2920 62580 2930 62640
rect 3690 62640 3770 62650
rect 3690 62580 3700 62640
rect 3760 62630 3770 62640
rect 4070 62640 4150 62650
rect 4070 62630 4080 62640
rect 3760 62600 4080 62630
rect 3760 62580 3770 62600
rect 2850 62570 2930 62580
rect 3270 62570 3350 62580
rect 3690 62570 3770 62580
rect 4070 62580 4080 62600
rect 4140 62580 4150 62640
rect 4070 62570 4150 62580
rect 7620 62640 7700 62650
rect 7620 62580 7630 62640
rect 7690 62630 7700 62640
rect 7840 62640 7920 62650
rect 7840 62630 7850 62640
rect 7690 62600 7850 62630
rect 7690 62580 7700 62600
rect 7620 62570 7700 62580
rect 7840 62580 7850 62600
rect 7910 62580 7920 62640
rect 8680 62640 8760 62650
rect 8680 62580 8690 62640
rect 8750 62630 8760 62640
rect 9060 62640 9140 62650
rect 9060 62630 9070 62640
rect 8750 62600 9070 62630
rect 8750 62580 8760 62600
rect 7840 62570 7920 62580
rect 8260 62570 8340 62580
rect 8680 62570 8760 62580
rect 9060 62580 9070 62600
rect 9130 62580 9140 62640
rect 9060 62570 9140 62580
rect 3270 62510 3280 62570
rect 3340 62530 3350 62570
rect 3340 62520 4040 62530
rect 3340 62510 3980 62520
rect 3270 62500 3980 62510
rect 8260 62510 8270 62570
rect 8330 62530 8340 62570
rect 8330 62520 9030 62530
rect 8330 62510 8970 62520
rect 8260 62500 8970 62510
rect 3980 62450 4040 62460
rect 8970 62450 9030 62460
rect 3920 61340 3980 61350
rect 3270 61310 3920 61320
rect 2650 61250 2710 61260
rect 3270 61250 3280 61310
rect 3340 61290 3920 61310
rect 3340 61250 3350 61290
rect 8910 61340 8970 61350
rect 3920 61270 3980 61280
rect 8260 61310 8910 61320
rect 4070 61250 4130 61260
rect 2850 61240 2930 61250
rect 3270 61240 3350 61250
rect 3690 61240 3770 61250
rect 2850 61230 2860 61240
rect 2710 61200 2860 61230
rect 2650 61180 2710 61190
rect 2850 61180 2860 61200
rect 2920 61180 2930 61240
rect 2850 61170 2930 61180
rect 3690 61180 3700 61240
rect 3760 61230 3770 61240
rect 3760 61200 4070 61230
rect 3760 61180 3770 61200
rect 4070 61180 4130 61190
rect 7640 61250 7700 61260
rect 8260 61250 8270 61310
rect 8330 61290 8910 61310
rect 8330 61250 8340 61290
rect 8910 61270 8970 61280
rect 9060 61250 9120 61260
rect 7840 61240 7920 61250
rect 8260 61240 8340 61250
rect 8680 61240 8760 61250
rect 7840 61230 7850 61240
rect 7700 61200 7850 61230
rect 7640 61180 7700 61190
rect 7840 61180 7850 61200
rect 7910 61180 7920 61240
rect 3690 61170 3770 61180
rect 7840 61170 7920 61180
rect 8680 61180 8690 61240
rect 8750 61230 8760 61240
rect 8750 61200 9060 61230
rect 8750 61180 8760 61200
rect 9060 61180 9120 61190
rect 8680 61170 8760 61180
rect 3260 61150 3360 61160
rect 3260 61080 3280 61150
rect 3350 61080 3360 61150
rect 3260 61040 3360 61080
rect 3260 60970 3280 61040
rect 3350 60970 3360 61040
rect 3260 60950 3360 60970
rect 8250 61150 8350 61160
rect 8250 61080 8270 61150
rect 8340 61080 8350 61150
rect 8250 61040 8350 61080
rect 8250 60970 8270 61040
rect 8340 60970 8350 61040
rect 8250 60950 8350 60970
rect 2630 60930 2710 60940
rect 2630 60870 2640 60930
rect 2700 60920 2710 60930
rect 2850 60930 2930 60940
rect 2850 60920 2860 60930
rect 2700 60890 2860 60920
rect 2700 60870 2710 60890
rect 2630 60860 2710 60870
rect 2850 60870 2860 60890
rect 2920 60870 2930 60930
rect 3690 60930 3770 60940
rect 3690 60870 3700 60930
rect 3760 60920 3770 60930
rect 4070 60930 4150 60940
rect 4070 60920 4080 60930
rect 3760 60890 4080 60920
rect 3760 60870 3770 60890
rect 2850 60860 2930 60870
rect 3270 60860 3350 60870
rect 3690 60860 3770 60870
rect 4070 60870 4080 60890
rect 4140 60870 4150 60930
rect 4070 60860 4150 60870
rect 7620 60930 7700 60940
rect 7620 60870 7630 60930
rect 7690 60920 7700 60930
rect 7840 60930 7920 60940
rect 7840 60920 7850 60930
rect 7690 60890 7850 60920
rect 7690 60870 7700 60890
rect 7620 60860 7700 60870
rect 7840 60870 7850 60890
rect 7910 60870 7920 60930
rect 8680 60930 8760 60940
rect 8680 60870 8690 60930
rect 8750 60920 8760 60930
rect 9060 60930 9140 60940
rect 9060 60920 9070 60930
rect 8750 60890 9070 60920
rect 8750 60870 8760 60890
rect 7840 60860 7920 60870
rect 8260 60860 8340 60870
rect 8680 60860 8760 60870
rect 9060 60870 9070 60890
rect 9130 60870 9140 60930
rect 9060 60860 9140 60870
rect 3270 60800 3280 60860
rect 3340 60820 3350 60860
rect 3340 60810 4040 60820
rect 3340 60800 3980 60810
rect 3270 60790 3980 60800
rect 8260 60800 8270 60860
rect 8330 60820 8340 60860
rect 8330 60810 9030 60820
rect 8330 60800 8970 60810
rect 8260 60790 8970 60800
rect 3980 60740 4040 60750
rect 8970 60740 9030 60750
rect 12540 59750 12570 67050
rect 12660 66590 12690 67050
rect 12610 66580 12690 66590
rect 12610 66520 12620 66580
rect 12680 66520 12690 66580
rect 12610 66510 12690 66520
rect 14050 66590 14080 67050
rect 14050 66580 14130 66590
rect 14050 66520 14060 66580
rect 14120 66520 14130 66580
rect 14050 66510 14130 66520
rect 13900 66470 13960 66480
rect 13250 66440 13900 66450
rect 12630 66380 12690 66390
rect 13250 66380 13260 66440
rect 13320 66420 13900 66440
rect 13320 66380 13330 66420
rect 13900 66400 13960 66410
rect 14050 66380 14110 66390
rect 12830 66370 12910 66380
rect 13250 66370 13330 66380
rect 13670 66370 13750 66380
rect 12830 66360 12840 66370
rect 12690 66330 12840 66360
rect 12630 66310 12690 66320
rect 12830 66310 12840 66330
rect 12900 66310 12910 66370
rect 12830 66300 12910 66310
rect 13670 66310 13680 66370
rect 13740 66360 13750 66370
rect 13740 66330 14050 66360
rect 13740 66310 13750 66330
rect 14050 66310 14110 66320
rect 13670 66300 13750 66310
rect 13240 66280 13340 66290
rect 13240 66210 13260 66280
rect 13330 66210 13340 66280
rect 13240 66170 13340 66210
rect 13240 66100 13260 66170
rect 13330 66100 13340 66170
rect 13240 66080 13340 66100
rect 12610 66060 12690 66070
rect 12610 66000 12620 66060
rect 12680 66050 12690 66060
rect 12830 66060 12910 66070
rect 12830 66050 12840 66060
rect 12680 66020 12840 66050
rect 12680 66000 12690 66020
rect 12610 65990 12690 66000
rect 12830 66000 12840 66020
rect 12900 66000 12910 66060
rect 13670 66060 13750 66070
rect 13670 66000 13680 66060
rect 13740 66050 13750 66060
rect 14050 66060 14130 66070
rect 14050 66050 14060 66060
rect 13740 66020 14060 66050
rect 13740 66000 13750 66020
rect 12830 65990 12910 66000
rect 13250 65990 13330 66000
rect 13670 65990 13750 66000
rect 14050 66000 14060 66020
rect 14120 66000 14130 66060
rect 14050 65990 14130 66000
rect 13250 65930 13260 65990
rect 13320 65950 13330 65990
rect 13320 65940 14020 65950
rect 13320 65930 13960 65940
rect 13250 65920 13960 65930
rect 13960 65870 14020 65880
rect 13900 64760 13960 64770
rect 13250 64730 13900 64740
rect 12630 64670 12690 64680
rect 13250 64670 13260 64730
rect 13320 64710 13900 64730
rect 13320 64670 13330 64710
rect 13900 64690 13960 64700
rect 14050 64670 14110 64680
rect 12830 64660 12910 64670
rect 13250 64660 13330 64670
rect 13670 64660 13750 64670
rect 12830 64650 12840 64660
rect 12690 64620 12840 64650
rect 12630 64600 12690 64610
rect 12830 64600 12840 64620
rect 12900 64600 12910 64660
rect 12830 64590 12910 64600
rect 13670 64600 13680 64660
rect 13740 64650 13750 64660
rect 13740 64620 14050 64650
rect 13740 64600 13750 64620
rect 14050 64600 14110 64610
rect 13670 64590 13750 64600
rect 13240 64570 13340 64580
rect 13240 64500 13260 64570
rect 13330 64500 13340 64570
rect 13240 64460 13340 64500
rect 13240 64390 13260 64460
rect 13330 64390 13340 64460
rect 13240 64370 13340 64390
rect 12610 64350 12690 64360
rect 12610 64290 12620 64350
rect 12680 64340 12690 64350
rect 12830 64350 12910 64360
rect 12830 64340 12840 64350
rect 12680 64310 12840 64340
rect 12680 64290 12690 64310
rect 12610 64280 12690 64290
rect 12830 64290 12840 64310
rect 12900 64290 12910 64350
rect 13670 64350 13750 64360
rect 13670 64290 13680 64350
rect 13740 64340 13750 64350
rect 14050 64350 14130 64360
rect 14050 64340 14060 64350
rect 13740 64310 14060 64340
rect 13740 64290 13750 64310
rect 12830 64280 12910 64290
rect 13250 64280 13330 64290
rect 13670 64280 13750 64290
rect 14050 64290 14060 64310
rect 14120 64290 14130 64350
rect 14050 64280 14130 64290
rect 13250 64220 13260 64280
rect 13320 64240 13330 64280
rect 13320 64230 14020 64240
rect 13320 64220 13960 64230
rect 13250 64210 13960 64220
rect 13960 64160 14020 64170
rect 13900 63050 13960 63060
rect 13250 63020 13900 63030
rect 12630 62960 12690 62970
rect 13250 62960 13260 63020
rect 13320 63000 13900 63020
rect 13320 62960 13330 63000
rect 13900 62980 13960 62990
rect 14050 62960 14110 62970
rect 12830 62950 12910 62960
rect 13250 62950 13330 62960
rect 13670 62950 13750 62960
rect 12830 62940 12840 62950
rect 12690 62910 12840 62940
rect 12630 62890 12690 62900
rect 12830 62890 12840 62910
rect 12900 62890 12910 62950
rect 12830 62880 12910 62890
rect 13670 62890 13680 62950
rect 13740 62940 13750 62950
rect 13740 62910 14050 62940
rect 13740 62890 13750 62910
rect 14050 62890 14110 62900
rect 13670 62880 13750 62890
rect 13240 62860 13340 62870
rect 13240 62790 13260 62860
rect 13330 62790 13340 62860
rect 13240 62750 13340 62790
rect 13240 62680 13260 62750
rect 13330 62680 13340 62750
rect 13240 62660 13340 62680
rect 12610 62640 12690 62650
rect 12610 62580 12620 62640
rect 12680 62630 12690 62640
rect 12830 62640 12910 62650
rect 12830 62630 12840 62640
rect 12680 62600 12840 62630
rect 12680 62580 12690 62600
rect 12610 62570 12690 62580
rect 12830 62580 12840 62600
rect 12900 62580 12910 62640
rect 13670 62640 13750 62650
rect 13670 62580 13680 62640
rect 13740 62630 13750 62640
rect 14050 62640 14130 62650
rect 14050 62630 14060 62640
rect 13740 62600 14060 62630
rect 13740 62580 13750 62600
rect 12830 62570 12910 62580
rect 13250 62570 13330 62580
rect 13670 62570 13750 62580
rect 14050 62580 14060 62600
rect 14120 62580 14130 62640
rect 14050 62570 14130 62580
rect 13250 62510 13260 62570
rect 13320 62530 13330 62570
rect 13320 62520 14020 62530
rect 13320 62510 13960 62520
rect 13250 62500 13960 62510
rect 13960 62450 14020 62460
rect 13900 61340 13960 61350
rect 13250 61310 13900 61320
rect 12630 61250 12690 61260
rect 13250 61250 13260 61310
rect 13320 61290 13900 61310
rect 13320 61250 13330 61290
rect 13900 61270 13960 61280
rect 14050 61250 14110 61260
rect 12830 61240 12910 61250
rect 13250 61240 13330 61250
rect 13670 61240 13750 61250
rect 12830 61230 12840 61240
rect 12690 61200 12840 61230
rect 12630 61180 12690 61190
rect 12830 61180 12840 61200
rect 12900 61180 12910 61240
rect 12830 61170 12910 61180
rect 13670 61180 13680 61240
rect 13740 61230 13750 61240
rect 13740 61200 14050 61230
rect 13740 61180 13750 61200
rect 14050 61180 14110 61190
rect 13670 61170 13750 61180
rect 13240 61150 13340 61160
rect 13240 61080 13260 61150
rect 13330 61080 13340 61150
rect 13240 61040 13340 61080
rect 13240 60970 13260 61040
rect 13330 60970 13340 61040
rect 13240 60950 13340 60970
rect 12610 60930 12690 60940
rect 12610 60870 12620 60930
rect 12680 60920 12690 60930
rect 12830 60930 12910 60940
rect 12830 60920 12840 60930
rect 12680 60890 12840 60920
rect 12680 60870 12690 60890
rect 12610 60860 12690 60870
rect 12830 60870 12840 60890
rect 12900 60870 12910 60930
rect 13670 60930 13750 60940
rect 13670 60870 13680 60930
rect 13740 60920 13750 60930
rect 14050 60930 14130 60940
rect 14050 60920 14060 60930
rect 13740 60890 14060 60920
rect 13740 60870 13750 60890
rect 12830 60860 12910 60870
rect 13250 60860 13330 60870
rect 13670 60860 13750 60870
rect 14050 60870 14060 60890
rect 14120 60870 14130 60930
rect 14050 60860 14130 60870
rect 13250 60800 13260 60860
rect 13320 60820 13330 60860
rect 13320 60810 14020 60820
rect 13320 60800 13960 60810
rect 13250 60790 13960 60800
rect 13960 60740 14020 60750
rect 12490 59740 12570 59750
rect 12490 59680 12500 59740
rect 12560 59680 12570 59740
rect 12490 59670 12570 59680
rect 14170 59750 14200 67050
rect 17530 59750 17560 67050
rect 17650 66590 17680 67050
rect 17600 66580 17680 66590
rect 17600 66520 17610 66580
rect 17670 66520 17680 66580
rect 17600 66510 17680 66520
rect 19040 66590 19070 67050
rect 19040 66580 19120 66590
rect 19040 66520 19050 66580
rect 19110 66520 19120 66580
rect 19040 66510 19120 66520
rect 18890 66470 18950 66480
rect 18240 66440 18890 66450
rect 17620 66380 17680 66390
rect 18240 66380 18250 66440
rect 18310 66420 18890 66440
rect 18310 66380 18320 66420
rect 18890 66400 18950 66410
rect 19040 66380 19100 66390
rect 17820 66370 17900 66380
rect 18240 66370 18320 66380
rect 18660 66370 18740 66380
rect 17820 66360 17830 66370
rect 17680 66330 17830 66360
rect 17620 66310 17680 66320
rect 17820 66310 17830 66330
rect 17890 66310 17900 66370
rect 17820 66300 17900 66310
rect 18660 66310 18670 66370
rect 18730 66360 18740 66370
rect 18730 66330 19040 66360
rect 18730 66310 18740 66330
rect 19040 66310 19100 66320
rect 18660 66300 18740 66310
rect 18230 66280 18330 66290
rect 18230 66210 18250 66280
rect 18320 66210 18330 66280
rect 18230 66170 18330 66210
rect 18230 66100 18250 66170
rect 18320 66100 18330 66170
rect 18230 66080 18330 66100
rect 17600 66060 17680 66070
rect 17600 66000 17610 66060
rect 17670 66050 17680 66060
rect 17820 66060 17900 66070
rect 17820 66050 17830 66060
rect 17670 66020 17830 66050
rect 17670 66000 17680 66020
rect 17600 65990 17680 66000
rect 17820 66000 17830 66020
rect 17890 66000 17900 66060
rect 18660 66060 18740 66070
rect 18660 66000 18670 66060
rect 18730 66050 18740 66060
rect 19040 66060 19120 66070
rect 19040 66050 19050 66060
rect 18730 66020 19050 66050
rect 18730 66000 18740 66020
rect 17820 65990 17900 66000
rect 18240 65990 18320 66000
rect 18660 65990 18740 66000
rect 19040 66000 19050 66020
rect 19110 66000 19120 66060
rect 19040 65990 19120 66000
rect 18240 65930 18250 65990
rect 18310 65950 18320 65990
rect 18310 65940 19010 65950
rect 18310 65930 18950 65940
rect 18240 65920 18950 65930
rect 18950 65870 19010 65880
rect 18890 64760 18950 64770
rect 18240 64730 18890 64740
rect 17620 64670 17680 64680
rect 18240 64670 18250 64730
rect 18310 64710 18890 64730
rect 18310 64670 18320 64710
rect 18890 64690 18950 64700
rect 19040 64670 19100 64680
rect 17820 64660 17900 64670
rect 18240 64660 18320 64670
rect 18660 64660 18740 64670
rect 17820 64650 17830 64660
rect 17680 64620 17830 64650
rect 17620 64600 17680 64610
rect 17820 64600 17830 64620
rect 17890 64600 17900 64660
rect 17820 64590 17900 64600
rect 18660 64600 18670 64660
rect 18730 64650 18740 64660
rect 18730 64620 19040 64650
rect 18730 64600 18740 64620
rect 19040 64600 19100 64610
rect 18660 64590 18740 64600
rect 18230 64570 18330 64580
rect 18230 64500 18250 64570
rect 18320 64500 18330 64570
rect 18230 64460 18330 64500
rect 18230 64390 18250 64460
rect 18320 64390 18330 64460
rect 18230 64370 18330 64390
rect 17600 64350 17680 64360
rect 17600 64290 17610 64350
rect 17670 64340 17680 64350
rect 17820 64350 17900 64360
rect 17820 64340 17830 64350
rect 17670 64310 17830 64340
rect 17670 64290 17680 64310
rect 17600 64280 17680 64290
rect 17820 64290 17830 64310
rect 17890 64290 17900 64350
rect 18660 64350 18740 64360
rect 18660 64290 18670 64350
rect 18730 64340 18740 64350
rect 19040 64350 19120 64360
rect 19040 64340 19050 64350
rect 18730 64310 19050 64340
rect 18730 64290 18740 64310
rect 17820 64280 17900 64290
rect 18240 64280 18320 64290
rect 18660 64280 18740 64290
rect 19040 64290 19050 64310
rect 19110 64290 19120 64350
rect 19040 64280 19120 64290
rect 18240 64220 18250 64280
rect 18310 64240 18320 64280
rect 18310 64230 19010 64240
rect 18310 64220 18950 64230
rect 18240 64210 18950 64220
rect 18950 64160 19010 64170
rect 18890 63050 18950 63060
rect 18240 63020 18890 63030
rect 17620 62960 17680 62970
rect 18240 62960 18250 63020
rect 18310 63000 18890 63020
rect 18310 62960 18320 63000
rect 18890 62980 18950 62990
rect 19040 62960 19100 62970
rect 17820 62950 17900 62960
rect 18240 62950 18320 62960
rect 18660 62950 18740 62960
rect 17820 62940 17830 62950
rect 17680 62910 17830 62940
rect 17620 62890 17680 62900
rect 17820 62890 17830 62910
rect 17890 62890 17900 62950
rect 17820 62880 17900 62890
rect 18660 62890 18670 62950
rect 18730 62940 18740 62950
rect 18730 62910 19040 62940
rect 18730 62890 18740 62910
rect 19040 62890 19100 62900
rect 18660 62880 18740 62890
rect 18230 62860 18330 62870
rect 18230 62790 18250 62860
rect 18320 62790 18330 62860
rect 18230 62750 18330 62790
rect 18230 62680 18250 62750
rect 18320 62680 18330 62750
rect 18230 62660 18330 62680
rect 17600 62640 17680 62650
rect 17600 62580 17610 62640
rect 17670 62630 17680 62640
rect 17820 62640 17900 62650
rect 17820 62630 17830 62640
rect 17670 62600 17830 62630
rect 17670 62580 17680 62600
rect 17600 62570 17680 62580
rect 17820 62580 17830 62600
rect 17890 62580 17900 62640
rect 18660 62640 18740 62650
rect 18660 62580 18670 62640
rect 18730 62630 18740 62640
rect 19040 62640 19120 62650
rect 19040 62630 19050 62640
rect 18730 62600 19050 62630
rect 18730 62580 18740 62600
rect 17820 62570 17900 62580
rect 18240 62570 18320 62580
rect 18660 62570 18740 62580
rect 19040 62580 19050 62600
rect 19110 62580 19120 62640
rect 19040 62570 19120 62580
rect 18240 62510 18250 62570
rect 18310 62530 18320 62570
rect 18310 62520 19010 62530
rect 18310 62510 18950 62520
rect 18240 62500 18950 62510
rect 18950 62450 19010 62460
rect 18890 61340 18950 61350
rect 18240 61310 18890 61320
rect 17620 61250 17680 61260
rect 18240 61250 18250 61310
rect 18310 61290 18890 61310
rect 18310 61250 18320 61290
rect 18890 61270 18950 61280
rect 19040 61250 19100 61260
rect 17820 61240 17900 61250
rect 18240 61240 18320 61250
rect 18660 61240 18740 61250
rect 17820 61230 17830 61240
rect 17680 61200 17830 61230
rect 17620 61180 17680 61190
rect 17820 61180 17830 61200
rect 17890 61180 17900 61240
rect 17820 61170 17900 61180
rect 18660 61180 18670 61240
rect 18730 61230 18740 61240
rect 18730 61200 19040 61230
rect 18730 61180 18740 61200
rect 19040 61180 19100 61190
rect 18660 61170 18740 61180
rect 18230 61150 18330 61160
rect 18230 61080 18250 61150
rect 18320 61080 18330 61150
rect 18230 61040 18330 61080
rect 18230 60970 18250 61040
rect 18320 60970 18330 61040
rect 18230 60950 18330 60970
rect 17600 60930 17680 60940
rect 17600 60870 17610 60930
rect 17670 60920 17680 60930
rect 17820 60930 17900 60940
rect 17820 60920 17830 60930
rect 17670 60890 17830 60920
rect 17670 60870 17680 60890
rect 17600 60860 17680 60870
rect 17820 60870 17830 60890
rect 17890 60870 17900 60930
rect 18660 60930 18740 60940
rect 18660 60870 18670 60930
rect 18730 60920 18740 60930
rect 19040 60930 19120 60940
rect 19040 60920 19050 60930
rect 18730 60890 19050 60920
rect 18730 60870 18740 60890
rect 17820 60860 17900 60870
rect 18240 60860 18320 60870
rect 18660 60860 18740 60870
rect 19040 60870 19050 60890
rect 19110 60870 19120 60930
rect 19040 60860 19120 60870
rect 18240 60800 18250 60860
rect 18310 60820 18320 60860
rect 18310 60810 19010 60820
rect 18310 60800 18950 60810
rect 18240 60790 18950 60800
rect 18950 60740 19010 60750
rect 14170 59740 14250 59750
rect 14170 59680 14180 59740
rect 14240 59680 14250 59740
rect 14170 59670 14250 59680
rect 17480 59740 17560 59750
rect 17480 59680 17490 59740
rect 17550 59680 17560 59740
rect 17480 59670 17560 59680
rect 19160 59750 19190 67050
rect 19160 59740 19240 59750
rect 19160 59680 19170 59740
rect 19230 59680 19240 59740
rect 19160 59670 19240 59680
rect 3920 59630 3980 59640
rect 3270 59600 3920 59610
rect 2650 59540 2710 59550
rect 3270 59540 3280 59600
rect 3340 59580 3920 59600
rect 3340 59540 3350 59580
rect 8910 59630 8970 59640
rect 3920 59560 3980 59570
rect 8260 59600 8910 59610
rect 4070 59540 4130 59550
rect 2850 59530 2930 59540
rect 3270 59530 3350 59540
rect 3690 59530 3770 59540
rect 2850 59520 2860 59530
rect 2710 59490 2860 59520
rect 2650 59470 2710 59480
rect 2850 59470 2860 59490
rect 2920 59470 2930 59530
rect 2850 59460 2930 59470
rect 3690 59470 3700 59530
rect 3760 59520 3770 59530
rect 3760 59490 4070 59520
rect 3760 59470 3770 59490
rect 4070 59470 4130 59480
rect 7640 59540 7700 59550
rect 8260 59540 8270 59600
rect 8330 59580 8910 59600
rect 8330 59540 8340 59580
rect 13900 59630 13960 59640
rect 8910 59560 8970 59570
rect 13250 59600 13900 59610
rect 9060 59540 9120 59550
rect 7840 59530 7920 59540
rect 8260 59530 8340 59540
rect 8680 59530 8760 59540
rect 7840 59520 7850 59530
rect 7700 59490 7850 59520
rect 7640 59470 7700 59480
rect 7840 59470 7850 59490
rect 7910 59470 7920 59530
rect 3690 59460 3770 59470
rect 7840 59460 7920 59470
rect 8680 59470 8690 59530
rect 8750 59520 8760 59530
rect 8750 59490 9060 59520
rect 8750 59470 8760 59490
rect 9060 59470 9120 59480
rect 12510 59540 12570 59550
rect 13250 59540 13260 59600
rect 13320 59580 13900 59600
rect 13320 59540 13330 59580
rect 18890 59630 18950 59640
rect 13900 59560 13960 59570
rect 18240 59600 18890 59610
rect 14170 59540 14230 59550
rect 12830 59530 12910 59540
rect 13250 59530 13330 59540
rect 13670 59530 13750 59540
rect 12830 59520 12840 59530
rect 12570 59490 12840 59520
rect 12510 59470 12570 59480
rect 12830 59470 12840 59490
rect 12900 59470 12910 59530
rect 8680 59460 8760 59470
rect 12830 59460 12910 59470
rect 13670 59470 13680 59530
rect 13740 59520 13750 59530
rect 13740 59490 14170 59520
rect 13740 59470 13750 59490
rect 14170 59470 14230 59480
rect 17500 59540 17560 59550
rect 18240 59540 18250 59600
rect 18310 59580 18890 59600
rect 18310 59540 18320 59580
rect 18890 59560 18950 59570
rect 19160 59540 19220 59550
rect 17820 59530 17900 59540
rect 18240 59530 18320 59540
rect 18660 59530 18740 59540
rect 17820 59520 17830 59530
rect 17560 59490 17830 59520
rect 17500 59470 17560 59480
rect 17820 59470 17830 59490
rect 17890 59470 17900 59530
rect 13670 59460 13750 59470
rect 17820 59460 17900 59470
rect 18660 59470 18670 59530
rect 18730 59520 18740 59530
rect 18730 59490 19160 59520
rect 18730 59470 18740 59490
rect 19160 59470 19220 59480
rect 18660 59460 18740 59470
rect 3260 59440 3360 59450
rect 3260 59370 3280 59440
rect 3350 59370 3360 59440
rect 3260 59330 3360 59370
rect 3260 59260 3280 59330
rect 3350 59260 3360 59330
rect 3260 59240 3360 59260
rect 8250 59440 8350 59450
rect 8250 59370 8270 59440
rect 8340 59370 8350 59440
rect 8250 59330 8350 59370
rect 8250 59260 8270 59330
rect 8340 59260 8350 59330
rect 8250 59240 8350 59260
rect 13240 59440 13340 59450
rect 13240 59370 13260 59440
rect 13330 59370 13340 59440
rect 13240 59330 13340 59370
rect 13240 59260 13260 59330
rect 13330 59260 13340 59330
rect 13240 59240 13340 59260
rect 18230 59440 18330 59450
rect 18230 59370 18250 59440
rect 18320 59370 18330 59440
rect 18230 59330 18330 59370
rect 18230 59260 18250 59330
rect 18320 59260 18330 59330
rect 18230 59240 18330 59260
rect 2630 59220 2710 59230
rect 2630 59160 2640 59220
rect 2700 59210 2710 59220
rect 2850 59220 2930 59230
rect 2850 59210 2860 59220
rect 2700 59180 2860 59210
rect 2700 59160 2710 59180
rect 2630 59150 2710 59160
rect 2850 59160 2860 59180
rect 2920 59160 2930 59220
rect 3690 59220 3770 59230
rect 3690 59160 3700 59220
rect 3760 59210 3770 59220
rect 4070 59220 4150 59230
rect 4070 59210 4080 59220
rect 3760 59180 4080 59210
rect 3760 59160 3770 59180
rect 2850 59150 2930 59160
rect 3270 59150 3350 59160
rect 3690 59150 3770 59160
rect 4070 59160 4080 59180
rect 4140 59160 4150 59220
rect 4070 59150 4150 59160
rect 7620 59220 7700 59230
rect 7620 59160 7630 59220
rect 7690 59210 7700 59220
rect 7840 59220 7920 59230
rect 7840 59210 7850 59220
rect 7690 59180 7850 59210
rect 7690 59160 7700 59180
rect 7620 59150 7700 59160
rect 7840 59160 7850 59180
rect 7910 59160 7920 59220
rect 8680 59220 8760 59230
rect 8680 59160 8690 59220
rect 8750 59210 8760 59220
rect 9060 59220 9140 59230
rect 9060 59210 9070 59220
rect 8750 59180 9070 59210
rect 8750 59160 8760 59180
rect 7840 59150 7920 59160
rect 8260 59150 8340 59160
rect 8680 59150 8760 59160
rect 9060 59160 9070 59180
rect 9130 59160 9140 59220
rect 9060 59150 9140 59160
rect 12490 59220 12570 59230
rect 12490 59160 12500 59220
rect 12560 59210 12570 59220
rect 12830 59220 12910 59230
rect 12830 59210 12840 59220
rect 12560 59180 12840 59210
rect 12560 59160 12570 59180
rect 12490 59150 12570 59160
rect 12830 59160 12840 59180
rect 12900 59160 12910 59220
rect 13670 59220 13750 59230
rect 13670 59160 13680 59220
rect 13740 59210 13750 59220
rect 14170 59220 14250 59230
rect 14170 59210 14180 59220
rect 13740 59180 14180 59210
rect 13740 59160 13750 59180
rect 12830 59150 12910 59160
rect 13250 59150 13330 59160
rect 13670 59150 13750 59160
rect 14170 59160 14180 59180
rect 14240 59160 14250 59220
rect 14170 59150 14250 59160
rect 17480 59220 17560 59230
rect 17480 59160 17490 59220
rect 17550 59210 17560 59220
rect 17820 59220 17900 59230
rect 17820 59210 17830 59220
rect 17550 59180 17830 59210
rect 17550 59160 17560 59180
rect 17480 59150 17560 59160
rect 17820 59160 17830 59180
rect 17890 59160 17900 59220
rect 18660 59220 18740 59230
rect 18660 59160 18670 59220
rect 18730 59210 18740 59220
rect 19160 59220 19240 59230
rect 19160 59210 19170 59220
rect 18730 59180 19170 59210
rect 18730 59160 18740 59180
rect 17820 59150 17900 59160
rect 18240 59150 18320 59160
rect 18660 59150 18740 59160
rect 19160 59160 19170 59180
rect 19230 59160 19240 59220
rect 19160 59150 19240 59160
rect 3270 59090 3280 59150
rect 3340 59110 3350 59150
rect 3340 59100 4040 59110
rect 3340 59090 3980 59100
rect 3270 59080 3980 59090
rect 8260 59090 8270 59150
rect 8330 59110 8340 59150
rect 8330 59100 9030 59110
rect 8330 59090 8970 59100
rect 8260 59080 8970 59090
rect 3980 59030 4040 59040
rect 13250 59090 13260 59150
rect 13320 59110 13330 59150
rect 13320 59100 14020 59110
rect 13320 59090 13960 59100
rect 13250 59080 13960 59090
rect 8970 59030 9030 59040
rect 18240 59090 18250 59150
rect 18310 59110 18320 59150
rect 18310 59100 19010 59110
rect 18310 59090 18950 59100
rect 18240 59080 18950 59090
rect 13960 59030 14020 59040
rect 18950 59030 19010 59040
rect 22280 58040 22310 67050
rect 22400 59750 22430 67050
rect 22520 63170 22550 67050
rect 22640 66590 22670 67050
rect 22590 66580 22670 66590
rect 22590 66520 22600 66580
rect 22660 66520 22670 66580
rect 22590 66510 22670 66520
rect 24030 66590 24060 67050
rect 24030 66580 24110 66590
rect 24030 66520 24040 66580
rect 24100 66520 24110 66580
rect 24030 66510 24110 66520
rect 23880 66470 23940 66480
rect 23230 66440 23880 66450
rect 22610 66380 22670 66390
rect 23230 66380 23240 66440
rect 23300 66420 23880 66440
rect 23300 66380 23310 66420
rect 23880 66400 23940 66410
rect 24030 66380 24090 66390
rect 22810 66370 22890 66380
rect 23230 66370 23310 66380
rect 23650 66370 23730 66380
rect 22810 66360 22820 66370
rect 22670 66330 22820 66360
rect 22610 66310 22670 66320
rect 22810 66310 22820 66330
rect 22880 66310 22890 66370
rect 22810 66300 22890 66310
rect 23650 66310 23660 66370
rect 23720 66360 23730 66370
rect 23720 66330 24030 66360
rect 23720 66310 23730 66330
rect 24030 66310 24090 66320
rect 23650 66300 23730 66310
rect 23220 66280 23320 66290
rect 23220 66210 23240 66280
rect 23310 66210 23320 66280
rect 23220 66170 23320 66210
rect 23220 66100 23240 66170
rect 23310 66100 23320 66170
rect 23220 66080 23320 66100
rect 22590 66060 22670 66070
rect 22590 66000 22600 66060
rect 22660 66050 22670 66060
rect 22810 66060 22890 66070
rect 22810 66050 22820 66060
rect 22660 66020 22820 66050
rect 22660 66000 22670 66020
rect 22590 65990 22670 66000
rect 22810 66000 22820 66020
rect 22880 66000 22890 66060
rect 23650 66060 23730 66070
rect 23650 66000 23660 66060
rect 23720 66050 23730 66060
rect 24030 66060 24110 66070
rect 24030 66050 24040 66060
rect 23720 66020 24040 66050
rect 23720 66000 23730 66020
rect 22810 65990 22890 66000
rect 23230 65990 23310 66000
rect 23650 65990 23730 66000
rect 24030 66000 24040 66020
rect 24100 66000 24110 66060
rect 24030 65990 24110 66000
rect 23230 65930 23240 65990
rect 23300 65950 23310 65990
rect 23300 65940 24000 65950
rect 23300 65930 23940 65940
rect 23230 65920 23940 65930
rect 23940 65870 24000 65880
rect 23880 64760 23940 64770
rect 23230 64730 23880 64740
rect 22610 64670 22670 64680
rect 23230 64670 23240 64730
rect 23300 64710 23880 64730
rect 23300 64670 23310 64710
rect 23880 64690 23940 64700
rect 24030 64670 24090 64680
rect 22810 64660 22890 64670
rect 23230 64660 23310 64670
rect 23650 64660 23730 64670
rect 22810 64650 22820 64660
rect 22670 64620 22820 64650
rect 22610 64600 22670 64610
rect 22810 64600 22820 64620
rect 22880 64600 22890 64660
rect 22810 64590 22890 64600
rect 23650 64600 23660 64660
rect 23720 64650 23730 64660
rect 23720 64620 24030 64650
rect 23720 64600 23730 64620
rect 24030 64600 24090 64610
rect 23650 64590 23730 64600
rect 23220 64570 23320 64580
rect 23220 64500 23240 64570
rect 23310 64500 23320 64570
rect 23220 64460 23320 64500
rect 23220 64390 23240 64460
rect 23310 64390 23320 64460
rect 23220 64370 23320 64390
rect 22590 64350 22670 64360
rect 22590 64290 22600 64350
rect 22660 64340 22670 64350
rect 22810 64350 22890 64360
rect 22810 64340 22820 64350
rect 22660 64310 22820 64340
rect 22660 64290 22670 64310
rect 22590 64280 22670 64290
rect 22810 64290 22820 64310
rect 22880 64290 22890 64350
rect 23650 64350 23730 64360
rect 23650 64290 23660 64350
rect 23720 64340 23730 64350
rect 24030 64350 24110 64360
rect 24030 64340 24040 64350
rect 23720 64310 24040 64340
rect 23720 64290 23730 64310
rect 22810 64280 22890 64290
rect 23230 64280 23310 64290
rect 23650 64280 23730 64290
rect 24030 64290 24040 64310
rect 24100 64290 24110 64350
rect 24030 64280 24110 64290
rect 23230 64220 23240 64280
rect 23300 64240 23310 64280
rect 23300 64230 24000 64240
rect 23300 64220 23940 64230
rect 23230 64210 23940 64220
rect 23940 64160 24000 64170
rect 22470 63160 22550 63170
rect 22470 63100 22480 63160
rect 22540 63100 22550 63160
rect 22470 63090 22550 63100
rect 24150 63170 24180 67050
rect 24150 63160 24230 63170
rect 24150 63100 24160 63160
rect 24220 63100 24230 63160
rect 24150 63090 24230 63100
rect 23880 63050 23940 63060
rect 23230 63020 23880 63030
rect 22490 62960 22550 62970
rect 23230 62960 23240 63020
rect 23300 63000 23880 63020
rect 23300 62960 23310 63000
rect 23880 62980 23940 62990
rect 24150 62960 24210 62970
rect 22810 62950 22890 62960
rect 23230 62950 23310 62960
rect 23650 62950 23730 62960
rect 22810 62940 22820 62950
rect 22550 62910 22820 62940
rect 22490 62890 22550 62900
rect 22810 62890 22820 62910
rect 22880 62890 22890 62950
rect 22810 62880 22890 62890
rect 23650 62890 23660 62950
rect 23720 62940 23730 62950
rect 23720 62910 24150 62940
rect 23720 62890 23730 62910
rect 24150 62890 24210 62900
rect 23650 62880 23730 62890
rect 23220 62860 23320 62870
rect 23220 62790 23240 62860
rect 23310 62790 23320 62860
rect 23220 62750 23320 62790
rect 23220 62680 23240 62750
rect 23310 62680 23320 62750
rect 23220 62660 23320 62680
rect 22470 62640 22550 62650
rect 22470 62580 22480 62640
rect 22540 62630 22550 62640
rect 22810 62640 22890 62650
rect 22810 62630 22820 62640
rect 22540 62600 22820 62630
rect 22540 62580 22550 62600
rect 22470 62570 22550 62580
rect 22810 62580 22820 62600
rect 22880 62580 22890 62640
rect 23650 62640 23730 62650
rect 23650 62580 23660 62640
rect 23720 62630 23730 62640
rect 24150 62640 24230 62650
rect 24150 62630 24160 62640
rect 23720 62600 24160 62630
rect 23720 62580 23730 62600
rect 22810 62570 22890 62580
rect 23230 62570 23310 62580
rect 23650 62570 23730 62580
rect 24150 62580 24160 62600
rect 24220 62580 24230 62640
rect 24150 62570 24230 62580
rect 23230 62510 23240 62570
rect 23300 62530 23310 62570
rect 23300 62520 24000 62530
rect 23300 62510 23940 62520
rect 23230 62500 23940 62510
rect 23940 62450 24000 62460
rect 23880 61340 23940 61350
rect 23230 61310 23880 61320
rect 23230 61250 23240 61310
rect 23300 61290 23880 61310
rect 23300 61250 23310 61290
rect 23880 61270 23940 61280
rect 22490 61240 22550 61250
rect 22810 61240 22890 61250
rect 23230 61240 23310 61250
rect 23650 61240 23730 61250
rect 22810 61230 22820 61240
rect 22550 61200 22820 61230
rect 22490 61170 22550 61180
rect 22810 61180 22820 61200
rect 22880 61180 22890 61240
rect 22810 61170 22890 61180
rect 23650 61180 23660 61240
rect 23720 61230 23730 61240
rect 24150 61240 24210 61250
rect 23720 61200 24150 61230
rect 23720 61180 23730 61200
rect 23650 61170 23730 61180
rect 24150 61170 24210 61180
rect 23220 61150 23320 61160
rect 23220 61080 23240 61150
rect 23310 61080 23320 61150
rect 23220 61040 23320 61080
rect 23220 60970 23240 61040
rect 23310 60970 23320 61040
rect 23220 60950 23320 60970
rect 22810 60930 22890 60940
rect 22470 60920 22550 60930
rect 22810 60920 22820 60930
rect 22470 60860 22480 60920
rect 22540 60890 22820 60920
rect 22540 60860 22550 60890
rect 22810 60870 22820 60890
rect 22880 60870 22890 60930
rect 23650 60930 23730 60940
rect 23650 60870 23660 60930
rect 23720 60920 23730 60930
rect 24150 60920 24230 60930
rect 23720 60890 24160 60920
rect 23720 60870 23730 60890
rect 22810 60860 22890 60870
rect 23230 60860 23310 60870
rect 23650 60860 23730 60870
rect 24150 60860 24160 60890
rect 24220 60860 24230 60920
rect 22470 60850 22550 60860
rect 23230 60800 23240 60860
rect 23300 60820 23310 60860
rect 24150 60850 24230 60860
rect 23300 60810 24000 60820
rect 23300 60800 23940 60810
rect 23230 60790 23940 60800
rect 23940 60740 24000 60750
rect 22350 59740 22430 59750
rect 22350 59680 22360 59740
rect 22420 59680 22430 59740
rect 22350 59670 22430 59680
rect 24270 59750 24300 67050
rect 24270 59740 24350 59750
rect 24270 59680 24280 59740
rect 24340 59680 24350 59740
rect 24270 59670 24350 59680
rect 23880 59630 23940 59640
rect 23230 59600 23880 59610
rect 22370 59540 22430 59550
rect 23230 59540 23240 59600
rect 23300 59580 23880 59600
rect 23300 59540 23310 59580
rect 23880 59560 23940 59570
rect 24270 59540 24330 59550
rect 22810 59530 22890 59540
rect 23230 59530 23310 59540
rect 23650 59530 23730 59540
rect 22810 59520 22820 59530
rect 22430 59490 22820 59520
rect 22370 59470 22430 59480
rect 22810 59470 22820 59490
rect 22880 59470 22890 59530
rect 22810 59460 22890 59470
rect 23650 59470 23660 59530
rect 23720 59520 23730 59530
rect 23720 59490 24270 59520
rect 23720 59470 23730 59490
rect 24270 59470 24330 59480
rect 23650 59460 23730 59470
rect 23220 59440 23320 59450
rect 23220 59370 23240 59440
rect 23310 59370 23320 59440
rect 23220 59330 23320 59370
rect 23220 59260 23240 59330
rect 23310 59260 23320 59330
rect 23220 59240 23320 59260
rect 22350 59220 22430 59230
rect 22350 59160 22360 59220
rect 22420 59210 22430 59220
rect 22810 59220 22890 59230
rect 22810 59210 22820 59220
rect 22420 59180 22820 59210
rect 22420 59160 22430 59180
rect 22350 59150 22430 59160
rect 22810 59160 22820 59180
rect 22880 59160 22890 59220
rect 23650 59220 23730 59230
rect 23650 59160 23660 59220
rect 23720 59210 23730 59220
rect 24270 59220 24350 59230
rect 24270 59210 24280 59220
rect 23720 59180 24280 59210
rect 23720 59160 23730 59180
rect 22810 59150 22890 59160
rect 23230 59150 23310 59160
rect 23650 59150 23730 59160
rect 24270 59160 24280 59180
rect 24340 59160 24350 59220
rect 24270 59150 24350 59160
rect 23230 59090 23240 59150
rect 23300 59110 23310 59150
rect 23300 59100 24000 59110
rect 23300 59090 23940 59100
rect 23230 59080 23940 59090
rect 23940 59030 24000 59040
rect 22230 58030 22310 58040
rect 22230 57970 22240 58030
rect 22300 57970 22310 58030
rect 22230 57960 22310 57970
rect 24390 58040 24420 67050
rect 27270 58040 27300 67050
rect 27390 59750 27420 67050
rect 27510 63170 27540 67050
rect 27630 66590 27660 67050
rect 27580 66580 27660 66590
rect 27580 66520 27590 66580
rect 27650 66520 27660 66580
rect 27580 66510 27660 66520
rect 29020 66590 29050 67050
rect 29020 66580 29100 66590
rect 29020 66520 29030 66580
rect 29090 66520 29100 66580
rect 29020 66510 29100 66520
rect 28870 66470 28930 66480
rect 28220 66440 28870 66450
rect 27600 66380 27660 66390
rect 28220 66380 28230 66440
rect 28290 66420 28870 66440
rect 28290 66380 28300 66420
rect 28870 66400 28930 66410
rect 29020 66380 29080 66390
rect 27800 66370 27880 66380
rect 28220 66370 28300 66380
rect 28640 66370 28720 66380
rect 27800 66360 27810 66370
rect 27660 66330 27810 66360
rect 27600 66310 27660 66320
rect 27800 66310 27810 66330
rect 27870 66310 27880 66370
rect 27800 66300 27880 66310
rect 28640 66310 28650 66370
rect 28710 66360 28720 66370
rect 28710 66330 29020 66360
rect 28710 66310 28720 66330
rect 29020 66310 29080 66320
rect 28640 66300 28720 66310
rect 28210 66280 28310 66290
rect 28210 66210 28230 66280
rect 28300 66210 28310 66280
rect 28210 66170 28310 66210
rect 28210 66100 28230 66170
rect 28300 66100 28310 66170
rect 28210 66080 28310 66100
rect 27580 66060 27660 66070
rect 27580 66000 27590 66060
rect 27650 66050 27660 66060
rect 27800 66060 27880 66070
rect 27800 66050 27810 66060
rect 27650 66020 27810 66050
rect 27650 66000 27660 66020
rect 27580 65990 27660 66000
rect 27800 66000 27810 66020
rect 27870 66000 27880 66060
rect 28640 66060 28720 66070
rect 28640 66000 28650 66060
rect 28710 66050 28720 66060
rect 29020 66060 29100 66070
rect 29020 66050 29030 66060
rect 28710 66020 29030 66050
rect 28710 66000 28720 66020
rect 27800 65990 27880 66000
rect 28220 65990 28300 66000
rect 28640 65990 28720 66000
rect 29020 66000 29030 66020
rect 29090 66000 29100 66060
rect 29020 65990 29100 66000
rect 28220 65930 28230 65990
rect 28290 65950 28300 65990
rect 28290 65940 28990 65950
rect 28290 65930 28930 65940
rect 28220 65920 28930 65930
rect 28930 65870 28990 65880
rect 28870 64760 28930 64770
rect 28220 64730 28870 64740
rect 27600 64670 27660 64680
rect 28220 64670 28230 64730
rect 28290 64710 28870 64730
rect 28290 64670 28300 64710
rect 28870 64690 28930 64700
rect 29020 64670 29080 64680
rect 27800 64660 27880 64670
rect 28220 64660 28300 64670
rect 28640 64660 28720 64670
rect 27800 64650 27810 64660
rect 27660 64620 27810 64650
rect 27600 64600 27660 64610
rect 27800 64600 27810 64620
rect 27870 64600 27880 64660
rect 27800 64590 27880 64600
rect 28640 64600 28650 64660
rect 28710 64650 28720 64660
rect 28710 64620 29020 64650
rect 28710 64600 28720 64620
rect 29020 64600 29080 64610
rect 28640 64590 28720 64600
rect 28210 64570 28310 64580
rect 28210 64500 28230 64570
rect 28300 64500 28310 64570
rect 28210 64460 28310 64500
rect 28210 64390 28230 64460
rect 28300 64390 28310 64460
rect 28210 64370 28310 64390
rect 27580 64350 27660 64360
rect 27580 64290 27590 64350
rect 27650 64340 27660 64350
rect 27800 64350 27880 64360
rect 27800 64340 27810 64350
rect 27650 64310 27810 64340
rect 27650 64290 27660 64310
rect 27580 64280 27660 64290
rect 27800 64290 27810 64310
rect 27870 64290 27880 64350
rect 28640 64350 28720 64360
rect 28640 64290 28650 64350
rect 28710 64340 28720 64350
rect 29020 64350 29100 64360
rect 29020 64340 29030 64350
rect 28710 64310 29030 64340
rect 28710 64290 28720 64310
rect 27800 64280 27880 64290
rect 28220 64280 28300 64290
rect 28640 64280 28720 64290
rect 29020 64290 29030 64310
rect 29090 64290 29100 64350
rect 29020 64280 29100 64290
rect 28220 64220 28230 64280
rect 28290 64240 28300 64280
rect 28290 64230 28990 64240
rect 28290 64220 28930 64230
rect 28220 64210 28930 64220
rect 28930 64160 28990 64170
rect 27460 63160 27540 63170
rect 27460 63100 27470 63160
rect 27530 63100 27540 63160
rect 27460 63090 27540 63100
rect 29140 63170 29170 67050
rect 29140 63160 29220 63170
rect 29140 63100 29150 63160
rect 29210 63100 29220 63160
rect 29140 63090 29220 63100
rect 28870 63050 28930 63060
rect 28220 63020 28870 63030
rect 27480 62960 27540 62970
rect 28220 62960 28230 63020
rect 28290 63000 28870 63020
rect 28290 62960 28300 63000
rect 28870 62980 28930 62990
rect 29140 62960 29200 62970
rect 27800 62950 27880 62960
rect 28220 62950 28300 62960
rect 28640 62950 28720 62960
rect 27800 62940 27810 62950
rect 27540 62910 27810 62940
rect 27480 62890 27540 62900
rect 27800 62890 27810 62910
rect 27870 62890 27880 62950
rect 27800 62880 27880 62890
rect 28640 62890 28650 62950
rect 28710 62940 28720 62950
rect 28710 62910 29140 62940
rect 28710 62890 28720 62910
rect 29140 62890 29200 62900
rect 28640 62880 28720 62890
rect 28210 62860 28310 62870
rect 28210 62790 28230 62860
rect 28300 62790 28310 62860
rect 28210 62750 28310 62790
rect 28210 62680 28230 62750
rect 28300 62680 28310 62750
rect 28210 62660 28310 62680
rect 27460 62640 27540 62650
rect 27460 62580 27470 62640
rect 27530 62630 27540 62640
rect 27800 62640 27880 62650
rect 27800 62630 27810 62640
rect 27530 62600 27810 62630
rect 27530 62580 27540 62600
rect 27460 62570 27540 62580
rect 27800 62580 27810 62600
rect 27870 62580 27880 62640
rect 28640 62640 28720 62650
rect 28640 62580 28650 62640
rect 28710 62630 28720 62640
rect 29140 62640 29220 62650
rect 29140 62630 29150 62640
rect 28710 62600 29150 62630
rect 28710 62580 28720 62600
rect 27800 62570 27880 62580
rect 28220 62570 28300 62580
rect 28640 62570 28720 62580
rect 29140 62580 29150 62600
rect 29210 62580 29220 62640
rect 29140 62570 29220 62580
rect 28220 62510 28230 62570
rect 28290 62530 28300 62570
rect 28290 62520 28990 62530
rect 28290 62510 28930 62520
rect 28220 62500 28930 62510
rect 28930 62450 28990 62460
rect 28870 61340 28930 61350
rect 28220 61310 28870 61320
rect 28220 61250 28230 61310
rect 28290 61290 28870 61310
rect 28290 61250 28300 61290
rect 28870 61270 28930 61280
rect 27480 61240 27540 61250
rect 27800 61240 27880 61250
rect 28220 61240 28300 61250
rect 28640 61240 28720 61250
rect 27800 61230 27810 61240
rect 27540 61200 27810 61230
rect 27480 61170 27540 61180
rect 27800 61180 27810 61200
rect 27870 61180 27880 61240
rect 27800 61170 27880 61180
rect 28640 61180 28650 61240
rect 28710 61230 28720 61240
rect 29140 61240 29200 61250
rect 28710 61200 29140 61230
rect 28710 61180 28720 61200
rect 28640 61170 28720 61180
rect 29140 61170 29200 61180
rect 28210 61150 28310 61160
rect 28210 61080 28230 61150
rect 28300 61080 28310 61150
rect 28210 61040 28310 61080
rect 28210 60970 28230 61040
rect 28300 60970 28310 61040
rect 28210 60950 28310 60970
rect 27800 60930 27880 60940
rect 27460 60920 27540 60930
rect 27800 60920 27810 60930
rect 27460 60860 27470 60920
rect 27530 60890 27810 60920
rect 27530 60860 27540 60890
rect 27800 60870 27810 60890
rect 27870 60870 27880 60930
rect 28640 60930 28720 60940
rect 28640 60870 28650 60930
rect 28710 60920 28720 60930
rect 29140 60920 29220 60930
rect 28710 60890 29150 60920
rect 28710 60870 28720 60890
rect 27800 60860 27880 60870
rect 28220 60860 28300 60870
rect 28640 60860 28720 60870
rect 29140 60860 29150 60890
rect 29210 60860 29220 60920
rect 27460 60850 27540 60860
rect 28220 60800 28230 60860
rect 28290 60820 28300 60860
rect 29140 60850 29220 60860
rect 28290 60810 28990 60820
rect 28290 60800 28930 60810
rect 28220 60790 28930 60800
rect 28930 60740 28990 60750
rect 27340 59740 27420 59750
rect 27340 59680 27350 59740
rect 27410 59680 27420 59740
rect 27340 59670 27420 59680
rect 29260 59750 29290 67050
rect 29260 59740 29340 59750
rect 29260 59680 29270 59740
rect 29330 59680 29340 59740
rect 29260 59670 29340 59680
rect 28870 59630 28930 59640
rect 28220 59600 28870 59610
rect 27360 59540 27420 59550
rect 28220 59540 28230 59600
rect 28290 59580 28870 59600
rect 28290 59540 28300 59580
rect 28870 59560 28930 59570
rect 29260 59540 29320 59550
rect 27800 59530 27880 59540
rect 28220 59530 28300 59540
rect 28640 59530 28720 59540
rect 27800 59520 27810 59530
rect 27420 59490 27810 59520
rect 27360 59470 27420 59480
rect 27800 59470 27810 59490
rect 27870 59470 27880 59530
rect 27800 59460 27880 59470
rect 28640 59470 28650 59530
rect 28710 59520 28720 59530
rect 28710 59490 29260 59520
rect 28710 59470 28720 59490
rect 29260 59470 29320 59480
rect 28640 59460 28720 59470
rect 28210 59440 28310 59450
rect 28210 59370 28230 59440
rect 28300 59370 28310 59440
rect 28210 59330 28310 59370
rect 28210 59260 28230 59330
rect 28300 59260 28310 59330
rect 28210 59240 28310 59260
rect 27340 59220 27420 59230
rect 27340 59160 27350 59220
rect 27410 59210 27420 59220
rect 27800 59220 27880 59230
rect 27800 59210 27810 59220
rect 27410 59180 27810 59210
rect 27410 59160 27420 59180
rect 27340 59150 27420 59160
rect 27800 59160 27810 59180
rect 27870 59160 27880 59220
rect 28640 59220 28720 59230
rect 28640 59160 28650 59220
rect 28710 59210 28720 59220
rect 29260 59220 29340 59230
rect 29260 59210 29270 59220
rect 28710 59180 29270 59210
rect 28710 59160 28720 59180
rect 27800 59150 27880 59160
rect 28220 59150 28300 59160
rect 28640 59150 28720 59160
rect 29260 59160 29270 59180
rect 29330 59160 29340 59220
rect 29260 59150 29340 59160
rect 28220 59090 28230 59150
rect 28290 59110 28300 59150
rect 28290 59100 28990 59110
rect 28290 59090 28930 59100
rect 28220 59080 28930 59090
rect 28930 59030 28990 59040
rect 24390 58030 24470 58040
rect 24390 57970 24400 58030
rect 24460 57970 24470 58030
rect 24390 57960 24470 57970
rect 27220 58030 27300 58040
rect 27220 57970 27230 58030
rect 27290 57970 27300 58030
rect 27220 57960 27300 57970
rect 29380 58040 29410 67050
rect 29380 58030 29460 58040
rect 29380 57970 29390 58030
rect 29450 57970 29460 58030
rect 29380 57960 29460 57970
rect 3920 57920 3980 57930
rect 3270 57890 3920 57900
rect 2650 57830 2710 57840
rect 3270 57830 3280 57890
rect 3340 57870 3920 57890
rect 3340 57830 3350 57870
rect 8910 57920 8970 57930
rect 3920 57850 3980 57860
rect 8260 57890 8910 57900
rect 4070 57830 4130 57840
rect 2850 57820 2930 57830
rect 3270 57820 3350 57830
rect 3690 57820 3770 57830
rect 2850 57810 2860 57820
rect 2710 57780 2860 57810
rect 2650 57760 2710 57770
rect 2850 57760 2860 57780
rect 2920 57760 2930 57820
rect 2850 57750 2930 57760
rect 3690 57760 3700 57820
rect 3760 57810 3770 57820
rect 3760 57780 4070 57810
rect 3760 57760 3770 57780
rect 4070 57760 4130 57770
rect 7640 57830 7700 57840
rect 8260 57830 8270 57890
rect 8330 57870 8910 57890
rect 8330 57830 8340 57870
rect 13900 57920 13960 57930
rect 8910 57850 8970 57860
rect 13250 57890 13900 57900
rect 9060 57830 9120 57840
rect 7840 57820 7920 57830
rect 8260 57820 8340 57830
rect 8680 57820 8760 57830
rect 7840 57810 7850 57820
rect 7700 57780 7850 57810
rect 7640 57760 7700 57770
rect 7840 57760 7850 57780
rect 7910 57760 7920 57820
rect 3690 57750 3770 57760
rect 7840 57750 7920 57760
rect 8680 57760 8690 57820
rect 8750 57810 8760 57820
rect 8750 57780 9060 57810
rect 8750 57760 8760 57780
rect 9060 57760 9120 57770
rect 12510 57830 12570 57840
rect 13250 57830 13260 57890
rect 13320 57870 13900 57890
rect 13320 57830 13330 57870
rect 18890 57920 18950 57930
rect 13900 57850 13960 57860
rect 18240 57890 18890 57900
rect 14170 57830 14230 57840
rect 12830 57820 12910 57830
rect 13250 57820 13330 57830
rect 13670 57820 13750 57830
rect 12830 57810 12840 57820
rect 12570 57780 12840 57810
rect 12510 57760 12570 57770
rect 12830 57760 12840 57780
rect 12900 57760 12910 57820
rect 8680 57750 8760 57760
rect 12830 57750 12910 57760
rect 13670 57760 13680 57820
rect 13740 57810 13750 57820
rect 13740 57780 14170 57810
rect 13740 57760 13750 57780
rect 14170 57760 14230 57770
rect 17500 57830 17560 57840
rect 18240 57830 18250 57890
rect 18310 57870 18890 57890
rect 18310 57830 18320 57870
rect 23880 57920 23940 57930
rect 18890 57850 18950 57860
rect 23230 57890 23880 57900
rect 19160 57830 19220 57840
rect 17820 57820 17900 57830
rect 18240 57820 18320 57830
rect 18660 57820 18740 57830
rect 17820 57810 17830 57820
rect 17560 57780 17830 57810
rect 17500 57760 17560 57770
rect 17820 57760 17830 57780
rect 17890 57760 17900 57820
rect 13670 57750 13750 57760
rect 17820 57750 17900 57760
rect 18660 57760 18670 57820
rect 18730 57810 18740 57820
rect 18730 57780 19160 57810
rect 18730 57760 18740 57780
rect 19160 57760 19220 57770
rect 22250 57830 22310 57840
rect 23230 57830 23240 57890
rect 23300 57870 23880 57890
rect 23300 57830 23310 57870
rect 28870 57920 28930 57930
rect 23880 57850 23940 57860
rect 28220 57890 28870 57900
rect 24390 57830 24450 57840
rect 22810 57820 22890 57830
rect 23230 57820 23310 57830
rect 23650 57820 23730 57830
rect 22810 57810 22820 57820
rect 22310 57780 22820 57810
rect 22250 57760 22310 57770
rect 22810 57760 22820 57780
rect 22880 57760 22890 57820
rect 18660 57750 18740 57760
rect 22810 57750 22890 57760
rect 23650 57760 23660 57820
rect 23720 57810 23730 57820
rect 23720 57780 24390 57810
rect 23720 57760 23730 57780
rect 24390 57760 24450 57770
rect 27240 57830 27300 57840
rect 28220 57830 28230 57890
rect 28290 57870 28870 57890
rect 28290 57830 28300 57870
rect 28870 57850 28930 57860
rect 29380 57830 29440 57840
rect 27800 57820 27880 57830
rect 28220 57820 28300 57830
rect 28640 57820 28720 57830
rect 27800 57810 27810 57820
rect 27300 57780 27810 57810
rect 27240 57760 27300 57770
rect 27800 57760 27810 57780
rect 27870 57760 27880 57820
rect 23650 57750 23730 57760
rect 27800 57750 27880 57760
rect 28640 57760 28650 57820
rect 28710 57810 28720 57820
rect 28710 57780 29380 57810
rect 28710 57760 28720 57780
rect 29380 57760 29440 57770
rect 28640 57750 28720 57760
rect 3260 57730 3360 57740
rect 3260 57660 3280 57730
rect 3350 57660 3360 57730
rect 3260 57620 3360 57660
rect 3260 57550 3280 57620
rect 3350 57550 3360 57620
rect 3260 57530 3360 57550
rect 8250 57730 8350 57740
rect 8250 57660 8270 57730
rect 8340 57660 8350 57730
rect 8250 57620 8350 57660
rect 8250 57550 8270 57620
rect 8340 57550 8350 57620
rect 8250 57530 8350 57550
rect 13240 57730 13340 57740
rect 13240 57660 13260 57730
rect 13330 57660 13340 57730
rect 13240 57620 13340 57660
rect 13240 57550 13260 57620
rect 13330 57550 13340 57620
rect 13240 57530 13340 57550
rect 18230 57730 18330 57740
rect 18230 57660 18250 57730
rect 18320 57660 18330 57730
rect 18230 57620 18330 57660
rect 18230 57550 18250 57620
rect 18320 57550 18330 57620
rect 18230 57530 18330 57550
rect 23220 57730 23320 57740
rect 23220 57660 23240 57730
rect 23310 57660 23320 57730
rect 23220 57620 23320 57660
rect 23220 57550 23240 57620
rect 23310 57550 23320 57620
rect 23220 57530 23320 57550
rect 28210 57730 28310 57740
rect 28210 57660 28230 57730
rect 28300 57660 28310 57730
rect 28210 57620 28310 57660
rect 28210 57550 28230 57620
rect 28300 57550 28310 57620
rect 28210 57530 28310 57550
rect 2630 57510 2710 57520
rect 2630 57450 2640 57510
rect 2700 57500 2710 57510
rect 2850 57510 2930 57520
rect 2850 57500 2860 57510
rect 2700 57470 2860 57500
rect 2700 57450 2710 57470
rect 2630 57440 2710 57450
rect 2850 57450 2860 57470
rect 2920 57450 2930 57510
rect 3690 57510 3770 57520
rect 3690 57450 3700 57510
rect 3760 57500 3770 57510
rect 4070 57510 4150 57520
rect 4070 57500 4080 57510
rect 3760 57470 4080 57500
rect 3760 57450 3770 57470
rect 2850 57440 2930 57450
rect 3270 57440 3350 57450
rect 3690 57440 3770 57450
rect 4070 57450 4080 57470
rect 4140 57450 4150 57510
rect 4070 57440 4150 57450
rect 7620 57510 7700 57520
rect 7620 57450 7630 57510
rect 7690 57500 7700 57510
rect 7840 57510 7920 57520
rect 7840 57500 7850 57510
rect 7690 57470 7850 57500
rect 7690 57450 7700 57470
rect 7620 57440 7700 57450
rect 7840 57450 7850 57470
rect 7910 57450 7920 57510
rect 8680 57510 8760 57520
rect 8680 57450 8690 57510
rect 8750 57500 8760 57510
rect 9060 57510 9140 57520
rect 9060 57500 9070 57510
rect 8750 57470 9070 57500
rect 8750 57450 8760 57470
rect 7840 57440 7920 57450
rect 8260 57440 8340 57450
rect 8680 57440 8760 57450
rect 9060 57450 9070 57470
rect 9130 57450 9140 57510
rect 9060 57440 9140 57450
rect 12490 57510 12570 57520
rect 12490 57450 12500 57510
rect 12560 57500 12570 57510
rect 12830 57510 12910 57520
rect 12830 57500 12840 57510
rect 12560 57470 12840 57500
rect 12560 57450 12570 57470
rect 12490 57440 12570 57450
rect 12830 57450 12840 57470
rect 12900 57450 12910 57510
rect 13670 57510 13750 57520
rect 13670 57450 13680 57510
rect 13740 57500 13750 57510
rect 14170 57510 14250 57520
rect 14170 57500 14180 57510
rect 13740 57470 14180 57500
rect 13740 57450 13750 57470
rect 12830 57440 12910 57450
rect 13250 57440 13330 57450
rect 13670 57440 13750 57450
rect 14170 57450 14180 57470
rect 14240 57450 14250 57510
rect 14170 57440 14250 57450
rect 17480 57510 17560 57520
rect 17480 57450 17490 57510
rect 17550 57500 17560 57510
rect 17820 57510 17900 57520
rect 17820 57500 17830 57510
rect 17550 57470 17830 57500
rect 17550 57450 17560 57470
rect 17480 57440 17560 57450
rect 17820 57450 17830 57470
rect 17890 57450 17900 57510
rect 18660 57510 18740 57520
rect 18660 57450 18670 57510
rect 18730 57500 18740 57510
rect 19160 57510 19240 57520
rect 19160 57500 19170 57510
rect 18730 57470 19170 57500
rect 18730 57450 18740 57470
rect 17820 57440 17900 57450
rect 18240 57440 18320 57450
rect 18660 57440 18740 57450
rect 19160 57450 19170 57470
rect 19230 57450 19240 57510
rect 19160 57440 19240 57450
rect 22230 57510 22310 57520
rect 22230 57450 22240 57510
rect 22300 57500 22310 57510
rect 22810 57510 22890 57520
rect 22810 57500 22820 57510
rect 22300 57470 22820 57500
rect 22300 57450 22310 57470
rect 22230 57440 22310 57450
rect 22810 57450 22820 57470
rect 22880 57450 22890 57510
rect 23650 57510 23730 57520
rect 23650 57450 23660 57510
rect 23720 57500 23730 57510
rect 24390 57510 24470 57520
rect 24390 57500 24400 57510
rect 23720 57470 24400 57500
rect 23720 57450 23730 57470
rect 22810 57440 22890 57450
rect 23230 57440 23310 57450
rect 23650 57440 23730 57450
rect 24390 57450 24400 57470
rect 24460 57450 24470 57510
rect 24390 57440 24470 57450
rect 27220 57510 27300 57520
rect 27220 57450 27230 57510
rect 27290 57500 27300 57510
rect 27800 57510 27880 57520
rect 27800 57500 27810 57510
rect 27290 57470 27810 57500
rect 27290 57450 27300 57470
rect 27220 57440 27300 57450
rect 27800 57450 27810 57470
rect 27870 57450 27880 57510
rect 28640 57510 28720 57520
rect 28640 57450 28650 57510
rect 28710 57500 28720 57510
rect 29380 57510 29460 57520
rect 29380 57500 29390 57510
rect 28710 57470 29390 57500
rect 28710 57450 28720 57470
rect 27800 57440 27880 57450
rect 28220 57440 28300 57450
rect 28640 57440 28720 57450
rect 29380 57450 29390 57470
rect 29450 57450 29460 57510
rect 29380 57440 29460 57450
rect 3270 57380 3280 57440
rect 3340 57400 3350 57440
rect 3340 57390 4040 57400
rect 3340 57380 3980 57390
rect 3270 57370 3980 57380
rect 8260 57380 8270 57440
rect 8330 57400 8340 57440
rect 8330 57390 9030 57400
rect 8330 57380 8970 57390
rect 8260 57370 8970 57380
rect 3980 57320 4040 57330
rect 13250 57380 13260 57440
rect 13320 57400 13330 57440
rect 13320 57390 14020 57400
rect 13320 57380 13960 57390
rect 13250 57370 13960 57380
rect 8970 57320 9030 57330
rect 18240 57380 18250 57440
rect 18310 57400 18320 57440
rect 18310 57390 19010 57400
rect 18310 57380 18950 57390
rect 18240 57370 18950 57380
rect 13960 57320 14020 57330
rect 23230 57380 23240 57440
rect 23300 57400 23310 57440
rect 23300 57390 24000 57400
rect 23300 57380 23940 57390
rect 23230 57370 23940 57380
rect 18950 57320 19010 57330
rect 28220 57380 28230 57440
rect 28290 57400 28300 57440
rect 28290 57390 28990 57400
rect 28290 57380 28930 57390
rect 28220 57370 28930 57380
rect 23940 57320 24000 57330
rect 28930 57320 28990 57330
rect 3920 56210 3980 56220
rect 3270 56180 3920 56190
rect 2650 56120 2710 56130
rect 3270 56120 3280 56180
rect 3340 56160 3920 56180
rect 3340 56120 3350 56160
rect 8910 56210 8970 56220
rect 3920 56140 3980 56150
rect 8260 56180 8910 56190
rect 4070 56120 4130 56130
rect 2850 56110 2930 56120
rect 3270 56110 3350 56120
rect 3690 56110 3770 56120
rect 2850 56100 2860 56110
rect 2710 56070 2860 56100
rect 2650 56050 2710 56060
rect 2850 56050 2860 56070
rect 2920 56050 2930 56110
rect 2850 56040 2930 56050
rect 3690 56050 3700 56110
rect 3760 56100 3770 56110
rect 3760 56070 4070 56100
rect 3760 56050 3770 56070
rect 4070 56050 4130 56060
rect 7640 56120 7700 56130
rect 8260 56120 8270 56180
rect 8330 56160 8910 56180
rect 8330 56120 8340 56160
rect 13900 56210 13960 56220
rect 8910 56140 8970 56150
rect 13250 56180 13900 56190
rect 9060 56120 9120 56130
rect 7840 56110 7920 56120
rect 8260 56110 8340 56120
rect 8680 56110 8760 56120
rect 7840 56100 7850 56110
rect 7700 56070 7850 56100
rect 7640 56050 7700 56060
rect 7840 56050 7850 56070
rect 7910 56050 7920 56110
rect 3690 56040 3770 56050
rect 7840 56040 7920 56050
rect 8680 56050 8690 56110
rect 8750 56100 8760 56110
rect 8750 56070 9060 56100
rect 8750 56050 8760 56070
rect 9060 56050 9120 56060
rect 12510 56120 12570 56130
rect 13250 56120 13260 56180
rect 13320 56160 13900 56180
rect 13320 56120 13330 56160
rect 18890 56210 18950 56220
rect 13900 56140 13960 56150
rect 18240 56180 18890 56190
rect 14170 56120 14230 56130
rect 12830 56110 12910 56120
rect 13250 56110 13330 56120
rect 13670 56110 13750 56120
rect 12830 56100 12840 56110
rect 12570 56070 12840 56100
rect 12510 56050 12570 56060
rect 12830 56050 12840 56070
rect 12900 56050 12910 56110
rect 8680 56040 8760 56050
rect 12830 56040 12910 56050
rect 13670 56050 13680 56110
rect 13740 56100 13750 56110
rect 13740 56070 14170 56100
rect 13740 56050 13750 56070
rect 14170 56050 14230 56060
rect 17500 56120 17560 56130
rect 18240 56120 18250 56180
rect 18310 56160 18890 56180
rect 18310 56120 18320 56160
rect 23880 56210 23940 56220
rect 18890 56140 18950 56150
rect 23230 56180 23880 56190
rect 19160 56120 19220 56130
rect 17820 56110 17900 56120
rect 18240 56110 18320 56120
rect 18660 56110 18740 56120
rect 17820 56100 17830 56110
rect 17560 56070 17830 56100
rect 17500 56050 17560 56060
rect 17820 56050 17830 56070
rect 17890 56050 17900 56110
rect 13670 56040 13750 56050
rect 17820 56040 17900 56050
rect 18660 56050 18670 56110
rect 18730 56100 18740 56110
rect 18730 56070 19160 56100
rect 18730 56050 18740 56070
rect 19160 56050 19220 56060
rect 22250 56120 22310 56130
rect 23230 56120 23240 56180
rect 23300 56160 23880 56180
rect 23300 56120 23310 56160
rect 28870 56210 28930 56220
rect 23880 56140 23940 56150
rect 28220 56180 28870 56190
rect 24390 56120 24450 56130
rect 22810 56110 22890 56120
rect 23230 56110 23310 56120
rect 23650 56110 23730 56120
rect 22810 56100 22820 56110
rect 22310 56070 22820 56100
rect 22250 56050 22310 56060
rect 22810 56050 22820 56070
rect 22880 56050 22890 56110
rect 18660 56040 18740 56050
rect 22810 56040 22890 56050
rect 23650 56050 23660 56110
rect 23720 56100 23730 56110
rect 23720 56070 24390 56100
rect 23720 56050 23730 56070
rect 24390 56050 24450 56060
rect 27240 56120 27300 56130
rect 28220 56120 28230 56180
rect 28290 56160 28870 56180
rect 28290 56120 28300 56160
rect 28870 56140 28930 56150
rect 29380 56120 29440 56130
rect 27800 56110 27880 56120
rect 28220 56110 28300 56120
rect 28640 56110 28720 56120
rect 27800 56100 27810 56110
rect 27300 56070 27810 56100
rect 27240 56050 27300 56060
rect 27800 56050 27810 56070
rect 27870 56050 27880 56110
rect 23650 56040 23730 56050
rect 27800 56040 27880 56050
rect 28640 56050 28650 56110
rect 28710 56100 28720 56110
rect 28710 56070 29380 56100
rect 28710 56050 28720 56070
rect 29380 56050 29440 56060
rect 28640 56040 28720 56050
rect 3260 56020 3360 56030
rect 3260 55950 3280 56020
rect 3350 55950 3360 56020
rect 3260 55910 3360 55950
rect 3260 55840 3280 55910
rect 3350 55840 3360 55910
rect 3260 55820 3360 55840
rect 8250 56020 8350 56030
rect 8250 55950 8270 56020
rect 8340 55950 8350 56020
rect 8250 55910 8350 55950
rect 8250 55840 8270 55910
rect 8340 55840 8350 55910
rect 8250 55820 8350 55840
rect 13240 56020 13340 56030
rect 13240 55950 13260 56020
rect 13330 55950 13340 56020
rect 13240 55910 13340 55950
rect 13240 55840 13260 55910
rect 13330 55840 13340 55910
rect 13240 55820 13340 55840
rect 18230 56020 18330 56030
rect 18230 55950 18250 56020
rect 18320 55950 18330 56020
rect 18230 55910 18330 55950
rect 18230 55840 18250 55910
rect 18320 55840 18330 55910
rect 18230 55820 18330 55840
rect 23220 56020 23320 56030
rect 23220 55950 23240 56020
rect 23310 55950 23320 56020
rect 23220 55910 23320 55950
rect 23220 55840 23240 55910
rect 23310 55840 23320 55910
rect 23220 55820 23320 55840
rect 28210 56020 28310 56030
rect 28210 55950 28230 56020
rect 28300 55950 28310 56020
rect 28210 55910 28310 55950
rect 28210 55840 28230 55910
rect 28300 55840 28310 55910
rect 28210 55820 28310 55840
rect 2630 55800 2710 55810
rect 2630 55740 2640 55800
rect 2700 55790 2710 55800
rect 2850 55800 2930 55810
rect 2850 55790 2860 55800
rect 2700 55760 2860 55790
rect 2700 55740 2710 55760
rect 2630 55730 2710 55740
rect 2850 55740 2860 55760
rect 2920 55740 2930 55800
rect 3690 55800 3770 55810
rect 3690 55740 3700 55800
rect 3760 55790 3770 55800
rect 4070 55800 4150 55810
rect 4070 55790 4080 55800
rect 3760 55760 4080 55790
rect 3760 55740 3770 55760
rect 2850 55730 2930 55740
rect 3270 55730 3350 55740
rect 3690 55730 3770 55740
rect 4070 55740 4080 55760
rect 4140 55740 4150 55800
rect 4070 55730 4150 55740
rect 7620 55800 7700 55810
rect 7620 55740 7630 55800
rect 7690 55790 7700 55800
rect 7840 55800 7920 55810
rect 7840 55790 7850 55800
rect 7690 55760 7850 55790
rect 7690 55740 7700 55760
rect 7620 55730 7700 55740
rect 7840 55740 7850 55760
rect 7910 55740 7920 55800
rect 8680 55800 8760 55810
rect 8680 55740 8690 55800
rect 8750 55790 8760 55800
rect 9060 55800 9140 55810
rect 9060 55790 9070 55800
rect 8750 55760 9070 55790
rect 8750 55740 8760 55760
rect 7840 55730 7920 55740
rect 8260 55730 8340 55740
rect 8680 55730 8760 55740
rect 9060 55740 9070 55760
rect 9130 55740 9140 55800
rect 9060 55730 9140 55740
rect 12490 55800 12570 55810
rect 12490 55740 12500 55800
rect 12560 55790 12570 55800
rect 12830 55800 12910 55810
rect 12830 55790 12840 55800
rect 12560 55760 12840 55790
rect 12560 55740 12570 55760
rect 12490 55730 12570 55740
rect 12830 55740 12840 55760
rect 12900 55740 12910 55800
rect 13670 55800 13750 55810
rect 13670 55740 13680 55800
rect 13740 55790 13750 55800
rect 14170 55800 14250 55810
rect 14170 55790 14180 55800
rect 13740 55760 14180 55790
rect 13740 55740 13750 55760
rect 12830 55730 12910 55740
rect 13250 55730 13330 55740
rect 13670 55730 13750 55740
rect 14170 55740 14180 55760
rect 14240 55740 14250 55800
rect 14170 55730 14250 55740
rect 17480 55800 17560 55810
rect 17480 55740 17490 55800
rect 17550 55790 17560 55800
rect 17820 55800 17900 55810
rect 17820 55790 17830 55800
rect 17550 55760 17830 55790
rect 17550 55740 17560 55760
rect 17480 55730 17560 55740
rect 17820 55740 17830 55760
rect 17890 55740 17900 55800
rect 18660 55800 18740 55810
rect 18660 55740 18670 55800
rect 18730 55790 18740 55800
rect 19160 55800 19240 55810
rect 19160 55790 19170 55800
rect 18730 55760 19170 55790
rect 18730 55740 18740 55760
rect 17820 55730 17900 55740
rect 18240 55730 18320 55740
rect 18660 55730 18740 55740
rect 19160 55740 19170 55760
rect 19230 55740 19240 55800
rect 19160 55730 19240 55740
rect 22230 55800 22310 55810
rect 22230 55740 22240 55800
rect 22300 55790 22310 55800
rect 22810 55800 22890 55810
rect 22810 55790 22820 55800
rect 22300 55760 22820 55790
rect 22300 55740 22310 55760
rect 22230 55730 22310 55740
rect 22810 55740 22820 55760
rect 22880 55740 22890 55800
rect 23650 55800 23730 55810
rect 23650 55740 23660 55800
rect 23720 55790 23730 55800
rect 24390 55800 24470 55810
rect 24390 55790 24400 55800
rect 23720 55760 24400 55790
rect 23720 55740 23730 55760
rect 22810 55730 22890 55740
rect 23230 55730 23310 55740
rect 23650 55730 23730 55740
rect 24390 55740 24400 55760
rect 24460 55740 24470 55800
rect 24390 55730 24470 55740
rect 27220 55800 27300 55810
rect 27220 55740 27230 55800
rect 27290 55790 27300 55800
rect 27800 55800 27880 55810
rect 27800 55790 27810 55800
rect 27290 55760 27810 55790
rect 27290 55740 27300 55760
rect 27220 55730 27300 55740
rect 27800 55740 27810 55760
rect 27870 55740 27880 55800
rect 28640 55800 28720 55810
rect 28640 55740 28650 55800
rect 28710 55790 28720 55800
rect 29380 55800 29460 55810
rect 29380 55790 29390 55800
rect 28710 55760 29390 55790
rect 28710 55740 28720 55760
rect 27800 55730 27880 55740
rect 28220 55730 28300 55740
rect 28640 55730 28720 55740
rect 29380 55740 29390 55760
rect 29450 55740 29460 55800
rect 29380 55730 29460 55740
rect 3270 55670 3280 55730
rect 3340 55690 3350 55730
rect 3340 55680 4040 55690
rect 3340 55670 3980 55680
rect 3270 55660 3980 55670
rect 8260 55670 8270 55730
rect 8330 55690 8340 55730
rect 8330 55680 9030 55690
rect 8330 55670 8970 55680
rect 8260 55660 8970 55670
rect 3980 55610 4040 55620
rect 13250 55670 13260 55730
rect 13320 55690 13330 55730
rect 13320 55680 14020 55690
rect 13320 55670 13960 55680
rect 13250 55660 13960 55670
rect 8970 55610 9030 55620
rect 18240 55670 18250 55730
rect 18310 55690 18320 55730
rect 18310 55680 19010 55690
rect 18310 55670 18950 55680
rect 18240 55660 18950 55670
rect 13960 55610 14020 55620
rect 23230 55670 23240 55730
rect 23300 55690 23310 55730
rect 23300 55680 24000 55690
rect 23300 55670 23940 55680
rect 23230 55660 23940 55670
rect 18950 55610 19010 55620
rect 28220 55670 28230 55730
rect 28290 55690 28300 55730
rect 28290 55680 28990 55690
rect 28290 55670 28930 55680
rect 28220 55660 28930 55670
rect 23940 55610 24000 55620
rect 28930 55610 28990 55620
rect 32020 54620 32050 67050
rect 32140 56330 32170 67050
rect 32260 58040 32290 67050
rect 32380 59750 32410 67050
rect 32500 63170 32530 67050
rect 32620 66590 32650 67050
rect 32570 66580 32650 66590
rect 32570 66520 32580 66580
rect 32640 66520 32650 66580
rect 32570 66510 32650 66520
rect 34010 66590 34040 67050
rect 34010 66580 34090 66590
rect 34010 66520 34020 66580
rect 34080 66520 34090 66580
rect 34010 66510 34090 66520
rect 33860 66470 33920 66480
rect 33210 66440 33860 66450
rect 32590 66380 32650 66390
rect 33210 66380 33220 66440
rect 33280 66420 33860 66440
rect 33280 66380 33290 66420
rect 33860 66400 33920 66410
rect 34010 66380 34070 66390
rect 32790 66370 32870 66380
rect 33210 66370 33290 66380
rect 33630 66370 33710 66380
rect 32790 66360 32800 66370
rect 32650 66330 32800 66360
rect 32590 66310 32650 66320
rect 32790 66310 32800 66330
rect 32860 66310 32870 66370
rect 32790 66300 32870 66310
rect 33630 66310 33640 66370
rect 33700 66360 33710 66370
rect 33700 66330 34010 66360
rect 33700 66310 33710 66330
rect 34010 66310 34070 66320
rect 33630 66300 33710 66310
rect 33200 66280 33300 66290
rect 33200 66210 33220 66280
rect 33290 66210 33300 66280
rect 33200 66170 33300 66210
rect 33200 66100 33220 66170
rect 33290 66100 33300 66170
rect 33200 66080 33300 66100
rect 32570 66060 32650 66070
rect 32570 66000 32580 66060
rect 32640 66050 32650 66060
rect 32790 66060 32870 66070
rect 32790 66050 32800 66060
rect 32640 66020 32800 66050
rect 32640 66000 32650 66020
rect 32570 65990 32650 66000
rect 32790 66000 32800 66020
rect 32860 66000 32870 66060
rect 33630 66060 33710 66070
rect 33630 66000 33640 66060
rect 33700 66050 33710 66060
rect 34010 66060 34090 66070
rect 34010 66050 34020 66060
rect 33700 66020 34020 66050
rect 33700 66000 33710 66020
rect 32790 65990 32870 66000
rect 33210 65990 33290 66000
rect 33630 65990 33710 66000
rect 34010 66000 34020 66020
rect 34080 66000 34090 66060
rect 34010 65990 34090 66000
rect 33210 65930 33220 65990
rect 33280 65950 33290 65990
rect 33280 65940 33980 65950
rect 33280 65930 33920 65940
rect 33210 65920 33920 65930
rect 33920 65870 33980 65880
rect 33860 64760 33920 64770
rect 33210 64730 33860 64740
rect 32590 64670 32650 64680
rect 33210 64670 33220 64730
rect 33280 64710 33860 64730
rect 33280 64670 33290 64710
rect 33860 64690 33920 64700
rect 34010 64670 34070 64680
rect 32790 64660 32870 64670
rect 33210 64660 33290 64670
rect 33630 64660 33710 64670
rect 32790 64650 32800 64660
rect 32650 64620 32800 64650
rect 32590 64600 32650 64610
rect 32790 64600 32800 64620
rect 32860 64600 32870 64660
rect 32790 64590 32870 64600
rect 33630 64600 33640 64660
rect 33700 64650 33710 64660
rect 33700 64620 34010 64650
rect 33700 64600 33710 64620
rect 34010 64600 34070 64610
rect 33630 64590 33710 64600
rect 33200 64570 33300 64580
rect 33200 64500 33220 64570
rect 33290 64500 33300 64570
rect 33200 64460 33300 64500
rect 33200 64390 33220 64460
rect 33290 64390 33300 64460
rect 33200 64370 33300 64390
rect 32570 64350 32650 64360
rect 32570 64290 32580 64350
rect 32640 64340 32650 64350
rect 32790 64350 32870 64360
rect 32790 64340 32800 64350
rect 32640 64310 32800 64340
rect 32640 64290 32650 64310
rect 32570 64280 32650 64290
rect 32790 64290 32800 64310
rect 32860 64290 32870 64350
rect 33630 64350 33710 64360
rect 33630 64290 33640 64350
rect 33700 64340 33710 64350
rect 34010 64350 34090 64360
rect 34010 64340 34020 64350
rect 33700 64310 34020 64340
rect 33700 64290 33710 64310
rect 32790 64280 32870 64290
rect 33210 64280 33290 64290
rect 33630 64280 33710 64290
rect 34010 64290 34020 64310
rect 34080 64290 34090 64350
rect 34010 64280 34090 64290
rect 33210 64220 33220 64280
rect 33280 64240 33290 64280
rect 33280 64230 33980 64240
rect 33280 64220 33920 64230
rect 33210 64210 33920 64220
rect 33920 64160 33980 64170
rect 32450 63160 32530 63170
rect 32450 63100 32460 63160
rect 32520 63100 32530 63160
rect 32450 63090 32530 63100
rect 34130 63170 34160 67050
rect 34130 63160 34210 63170
rect 34130 63100 34140 63160
rect 34200 63100 34210 63160
rect 34130 63090 34210 63100
rect 33860 63050 33920 63060
rect 33210 63020 33860 63030
rect 32470 62960 32530 62970
rect 33210 62960 33220 63020
rect 33280 63000 33860 63020
rect 33280 62960 33290 63000
rect 33860 62980 33920 62990
rect 34130 62960 34190 62970
rect 32790 62950 32870 62960
rect 33210 62950 33290 62960
rect 33630 62950 33710 62960
rect 32790 62940 32800 62950
rect 32530 62910 32800 62940
rect 32470 62890 32530 62900
rect 32790 62890 32800 62910
rect 32860 62890 32870 62950
rect 32790 62880 32870 62890
rect 33630 62890 33640 62950
rect 33700 62940 33710 62950
rect 33700 62910 34130 62940
rect 33700 62890 33710 62910
rect 34130 62890 34190 62900
rect 33630 62880 33710 62890
rect 33200 62860 33300 62870
rect 33200 62790 33220 62860
rect 33290 62790 33300 62860
rect 33200 62750 33300 62790
rect 33200 62680 33220 62750
rect 33290 62680 33300 62750
rect 33200 62660 33300 62680
rect 32450 62640 32530 62650
rect 32450 62580 32460 62640
rect 32520 62630 32530 62640
rect 32790 62640 32870 62650
rect 32790 62630 32800 62640
rect 32520 62600 32800 62630
rect 32520 62580 32530 62600
rect 32450 62570 32530 62580
rect 32790 62580 32800 62600
rect 32860 62580 32870 62640
rect 33630 62640 33710 62650
rect 33630 62580 33640 62640
rect 33700 62630 33710 62640
rect 34130 62640 34210 62650
rect 34130 62630 34140 62640
rect 33700 62600 34140 62630
rect 33700 62580 33710 62600
rect 32790 62570 32870 62580
rect 33210 62570 33290 62580
rect 33630 62570 33710 62580
rect 34130 62580 34140 62600
rect 34200 62580 34210 62640
rect 34130 62570 34210 62580
rect 33210 62510 33220 62570
rect 33280 62530 33290 62570
rect 33280 62520 33980 62530
rect 33280 62510 33920 62520
rect 33210 62500 33920 62510
rect 33920 62450 33980 62460
rect 33860 61340 33920 61350
rect 33210 61310 33860 61320
rect 32470 61250 32530 61260
rect 33210 61250 33220 61310
rect 33280 61290 33860 61310
rect 33280 61250 33290 61290
rect 33860 61270 33920 61280
rect 34130 61250 34190 61260
rect 32790 61240 32870 61250
rect 33210 61240 33290 61250
rect 33630 61240 33710 61250
rect 32790 61230 32800 61240
rect 32530 61200 32800 61230
rect 32470 61180 32530 61190
rect 32790 61180 32800 61200
rect 32860 61180 32870 61240
rect 32790 61170 32870 61180
rect 33630 61180 33640 61240
rect 33700 61230 33710 61240
rect 33700 61200 34130 61230
rect 33700 61180 33710 61200
rect 34130 61180 34190 61190
rect 33630 61170 33710 61180
rect 33200 61150 33300 61160
rect 33200 61080 33220 61150
rect 33290 61080 33300 61150
rect 33200 61040 33300 61080
rect 33200 60970 33220 61040
rect 33290 60970 33300 61040
rect 33200 60950 33300 60970
rect 32450 60930 32530 60940
rect 32450 60870 32460 60930
rect 32520 60920 32530 60930
rect 32790 60930 32870 60940
rect 32790 60920 32800 60930
rect 32520 60890 32800 60920
rect 32520 60870 32530 60890
rect 32450 60860 32530 60870
rect 32790 60870 32800 60890
rect 32860 60870 32870 60930
rect 33630 60930 33710 60940
rect 33630 60870 33640 60930
rect 33700 60920 33710 60930
rect 34130 60930 34210 60940
rect 34130 60920 34140 60930
rect 33700 60890 34140 60920
rect 33700 60870 33710 60890
rect 32790 60860 32870 60870
rect 33210 60860 33290 60870
rect 33630 60860 33710 60870
rect 34130 60870 34140 60890
rect 34200 60870 34210 60930
rect 34130 60860 34210 60870
rect 33210 60800 33220 60860
rect 33280 60820 33290 60860
rect 33280 60810 33980 60820
rect 33280 60800 33920 60810
rect 33210 60790 33920 60800
rect 33920 60740 33980 60750
rect 32330 59740 32410 59750
rect 32330 59680 32340 59740
rect 32400 59680 32410 59740
rect 32330 59670 32410 59680
rect 34250 59750 34280 67050
rect 34250 59740 34330 59750
rect 34250 59680 34260 59740
rect 34320 59680 34330 59740
rect 34250 59670 34330 59680
rect 33860 59630 33920 59640
rect 33210 59600 33860 59610
rect 32350 59540 32410 59550
rect 33210 59540 33220 59600
rect 33280 59580 33860 59600
rect 33280 59540 33290 59580
rect 33860 59560 33920 59570
rect 34250 59540 34310 59550
rect 32790 59530 32870 59540
rect 33210 59530 33290 59540
rect 33630 59530 33710 59540
rect 32790 59520 32800 59530
rect 32410 59490 32800 59520
rect 32350 59470 32410 59480
rect 32790 59470 32800 59490
rect 32860 59470 32870 59530
rect 32790 59460 32870 59470
rect 33630 59470 33640 59530
rect 33700 59520 33710 59530
rect 33700 59490 34250 59520
rect 33700 59470 33710 59490
rect 34250 59470 34310 59480
rect 33630 59460 33710 59470
rect 33200 59440 33300 59450
rect 33200 59370 33220 59440
rect 33290 59370 33300 59440
rect 33200 59330 33300 59370
rect 33200 59260 33220 59330
rect 33290 59260 33300 59330
rect 33200 59240 33300 59260
rect 32330 59220 32410 59230
rect 32330 59160 32340 59220
rect 32400 59210 32410 59220
rect 32790 59220 32870 59230
rect 32790 59210 32800 59220
rect 32400 59180 32800 59210
rect 32400 59160 32410 59180
rect 32330 59150 32410 59160
rect 32790 59160 32800 59180
rect 32860 59160 32870 59220
rect 33630 59220 33710 59230
rect 33630 59160 33640 59220
rect 33700 59210 33710 59220
rect 34250 59220 34330 59230
rect 34250 59210 34260 59220
rect 33700 59180 34260 59210
rect 33700 59160 33710 59180
rect 32790 59150 32870 59160
rect 33210 59150 33290 59160
rect 33630 59150 33710 59160
rect 34250 59160 34260 59180
rect 34320 59160 34330 59220
rect 34250 59150 34330 59160
rect 33210 59090 33220 59150
rect 33280 59110 33290 59150
rect 33280 59100 33980 59110
rect 33280 59090 33920 59100
rect 33210 59080 33920 59090
rect 33920 59030 33980 59040
rect 32210 58030 32290 58040
rect 32210 57970 32220 58030
rect 32280 57970 32290 58030
rect 32210 57960 32290 57970
rect 34370 58040 34400 67050
rect 34370 58030 34450 58040
rect 34370 57970 34380 58030
rect 34440 57970 34450 58030
rect 34370 57960 34450 57970
rect 33860 57920 33920 57930
rect 33210 57890 33860 57900
rect 32230 57830 32290 57840
rect 33210 57830 33220 57890
rect 33280 57870 33860 57890
rect 33280 57830 33290 57870
rect 33860 57850 33920 57860
rect 34370 57830 34430 57840
rect 32790 57820 32870 57830
rect 33210 57820 33290 57830
rect 33630 57820 33710 57830
rect 32790 57810 32800 57820
rect 32290 57780 32800 57810
rect 32230 57760 32290 57770
rect 32790 57760 32800 57780
rect 32860 57760 32870 57820
rect 32790 57750 32870 57760
rect 33630 57760 33640 57820
rect 33700 57810 33710 57820
rect 33700 57780 34370 57810
rect 33700 57760 33710 57780
rect 34370 57760 34430 57770
rect 33630 57750 33710 57760
rect 33200 57730 33300 57740
rect 33200 57660 33220 57730
rect 33290 57660 33300 57730
rect 33200 57620 33300 57660
rect 33200 57550 33220 57620
rect 33290 57550 33300 57620
rect 33200 57530 33300 57550
rect 32210 57510 32290 57520
rect 32210 57450 32220 57510
rect 32280 57500 32290 57510
rect 32790 57510 32870 57520
rect 32790 57500 32800 57510
rect 32280 57470 32800 57500
rect 32280 57450 32290 57470
rect 32210 57440 32290 57450
rect 32790 57450 32800 57470
rect 32860 57450 32870 57510
rect 33630 57510 33710 57520
rect 33630 57450 33640 57510
rect 33700 57500 33710 57510
rect 34370 57510 34450 57520
rect 34370 57500 34380 57510
rect 33700 57470 34380 57500
rect 33700 57450 33710 57470
rect 32790 57440 32870 57450
rect 33210 57440 33290 57450
rect 33630 57440 33710 57450
rect 34370 57450 34380 57470
rect 34440 57450 34450 57510
rect 34370 57440 34450 57450
rect 33210 57380 33220 57440
rect 33280 57400 33290 57440
rect 33280 57390 33980 57400
rect 33280 57380 33920 57390
rect 33210 57370 33920 57380
rect 33920 57320 33980 57330
rect 32090 56320 32170 56330
rect 32090 56260 32100 56320
rect 32160 56260 32170 56320
rect 32090 56250 32170 56260
rect 34490 56330 34520 67050
rect 34490 56320 34570 56330
rect 34490 56260 34500 56320
rect 34560 56260 34570 56320
rect 34490 56250 34570 56260
rect 33860 56210 33920 56220
rect 33210 56180 33860 56190
rect 32110 56120 32170 56130
rect 33210 56120 33220 56180
rect 33280 56160 33860 56180
rect 33280 56120 33290 56160
rect 33860 56140 33920 56150
rect 34490 56120 34550 56130
rect 32790 56110 32870 56120
rect 33210 56110 33290 56120
rect 33630 56110 33710 56120
rect 32790 56100 32800 56110
rect 32170 56070 32800 56100
rect 32110 56050 32170 56060
rect 32790 56050 32800 56070
rect 32860 56050 32870 56110
rect 32790 56040 32870 56050
rect 33630 56050 33640 56110
rect 33700 56100 33710 56110
rect 33700 56070 34490 56100
rect 33700 56050 33710 56070
rect 34490 56050 34550 56060
rect 33630 56040 33710 56050
rect 33200 56020 33300 56030
rect 33200 55950 33220 56020
rect 33290 55950 33300 56020
rect 33200 55910 33300 55950
rect 33200 55840 33220 55910
rect 33290 55840 33300 55910
rect 33200 55820 33300 55840
rect 32090 55800 32170 55810
rect 32090 55740 32100 55800
rect 32160 55790 32170 55800
rect 32790 55800 32870 55810
rect 32790 55790 32800 55800
rect 32160 55760 32800 55790
rect 32160 55740 32170 55760
rect 32090 55730 32170 55740
rect 32790 55740 32800 55760
rect 32860 55740 32870 55800
rect 33630 55800 33710 55810
rect 33630 55740 33640 55800
rect 33700 55790 33710 55800
rect 34490 55800 34570 55810
rect 34490 55790 34500 55800
rect 33700 55760 34500 55790
rect 33700 55740 33710 55760
rect 32790 55730 32870 55740
rect 33210 55730 33290 55740
rect 33630 55730 33710 55740
rect 34490 55740 34500 55760
rect 34560 55740 34570 55800
rect 34490 55730 34570 55740
rect 33210 55670 33220 55730
rect 33280 55690 33290 55730
rect 33280 55680 33980 55690
rect 33280 55670 33920 55680
rect 33210 55660 33920 55670
rect 33920 55610 33980 55620
rect 31970 54610 32050 54620
rect 31970 54550 31980 54610
rect 32040 54550 32050 54610
rect 31970 54540 32050 54550
rect 34610 54620 34640 67050
rect 34610 54610 34690 54620
rect 34610 54550 34620 54610
rect 34680 54550 34690 54610
rect 34610 54540 34690 54550
rect 3920 54500 3980 54510
rect 3270 54470 3920 54480
rect 2650 54410 2710 54420
rect 3270 54410 3280 54470
rect 3340 54450 3920 54470
rect 3340 54410 3350 54450
rect 8910 54500 8970 54510
rect 3920 54430 3980 54440
rect 8260 54470 8910 54480
rect 4070 54410 4130 54420
rect 2850 54400 2930 54410
rect 3270 54400 3350 54410
rect 3690 54400 3770 54410
rect 2850 54390 2860 54400
rect 2710 54360 2860 54390
rect 2650 54340 2710 54350
rect 2850 54340 2860 54360
rect 2920 54340 2930 54400
rect 2850 54330 2930 54340
rect 3690 54340 3700 54400
rect 3760 54390 3770 54400
rect 3760 54360 4070 54390
rect 3760 54340 3770 54360
rect 4070 54340 4130 54350
rect 7640 54410 7700 54420
rect 8260 54410 8270 54470
rect 8330 54450 8910 54470
rect 8330 54410 8340 54450
rect 13900 54500 13960 54510
rect 8910 54430 8970 54440
rect 13250 54470 13900 54480
rect 9060 54410 9120 54420
rect 7840 54400 7920 54410
rect 8260 54400 8340 54410
rect 8680 54400 8760 54410
rect 7840 54390 7850 54400
rect 7700 54360 7850 54390
rect 7640 54340 7700 54350
rect 7840 54340 7850 54360
rect 7910 54340 7920 54400
rect 3690 54330 3770 54340
rect 7840 54330 7920 54340
rect 8680 54340 8690 54400
rect 8750 54390 8760 54400
rect 8750 54360 9060 54390
rect 8750 54340 8760 54360
rect 9060 54340 9120 54350
rect 12510 54410 12570 54420
rect 13250 54410 13260 54470
rect 13320 54450 13900 54470
rect 13320 54410 13330 54450
rect 18890 54500 18950 54510
rect 13900 54430 13960 54440
rect 18240 54470 18890 54480
rect 14170 54410 14230 54420
rect 12830 54400 12910 54410
rect 13250 54400 13330 54410
rect 13670 54400 13750 54410
rect 12830 54390 12840 54400
rect 12570 54360 12840 54390
rect 12510 54340 12570 54350
rect 12830 54340 12840 54360
rect 12900 54340 12910 54400
rect 8680 54330 8760 54340
rect 12830 54330 12910 54340
rect 13670 54340 13680 54400
rect 13740 54390 13750 54400
rect 13740 54360 14170 54390
rect 13740 54340 13750 54360
rect 14170 54340 14230 54350
rect 17500 54410 17560 54420
rect 18240 54410 18250 54470
rect 18310 54450 18890 54470
rect 18310 54410 18320 54450
rect 23880 54500 23940 54510
rect 18890 54430 18950 54440
rect 23230 54470 23880 54480
rect 19160 54410 19220 54420
rect 17820 54400 17900 54410
rect 18240 54400 18320 54410
rect 18660 54400 18740 54410
rect 17820 54390 17830 54400
rect 17560 54360 17830 54390
rect 17500 54340 17560 54350
rect 17820 54340 17830 54360
rect 17890 54340 17900 54400
rect 13670 54330 13750 54340
rect 17820 54330 17900 54340
rect 18660 54340 18670 54400
rect 18730 54390 18740 54400
rect 18730 54360 19160 54390
rect 18730 54340 18740 54360
rect 19160 54340 19220 54350
rect 22250 54410 22310 54420
rect 23230 54410 23240 54470
rect 23300 54450 23880 54470
rect 23300 54410 23310 54450
rect 28870 54500 28930 54510
rect 23880 54430 23940 54440
rect 28220 54470 28870 54480
rect 24390 54410 24450 54420
rect 22810 54400 22890 54410
rect 23230 54400 23310 54410
rect 23650 54400 23730 54410
rect 22810 54390 22820 54400
rect 22310 54360 22820 54390
rect 22250 54340 22310 54350
rect 22810 54340 22820 54360
rect 22880 54340 22890 54400
rect 18660 54330 18740 54340
rect 22810 54330 22890 54340
rect 23650 54340 23660 54400
rect 23720 54390 23730 54400
rect 23720 54360 24390 54390
rect 23720 54340 23730 54360
rect 24390 54340 24450 54350
rect 27240 54410 27300 54420
rect 28220 54410 28230 54470
rect 28290 54450 28870 54470
rect 28290 54410 28300 54450
rect 33860 54500 33920 54510
rect 28870 54430 28930 54440
rect 33210 54470 33860 54480
rect 29380 54410 29440 54420
rect 27800 54400 27880 54410
rect 28220 54400 28300 54410
rect 28640 54400 28720 54410
rect 27800 54390 27810 54400
rect 27300 54360 27810 54390
rect 27240 54340 27300 54350
rect 27800 54340 27810 54360
rect 27870 54340 27880 54400
rect 23650 54330 23730 54340
rect 27800 54330 27880 54340
rect 28640 54340 28650 54400
rect 28710 54390 28720 54400
rect 28710 54360 29380 54390
rect 28710 54340 28720 54360
rect 29380 54340 29440 54350
rect 31990 54410 32050 54420
rect 33210 54410 33220 54470
rect 33280 54450 33860 54470
rect 33280 54410 33290 54450
rect 36890 54470 36920 67050
rect 37010 54620 37040 67050
rect 37130 56340 37160 67050
rect 37250 58050 37280 67050
rect 37370 59760 37400 67050
rect 37490 63180 37520 67050
rect 37610 66600 37640 67050
rect 37560 66590 37640 66600
rect 37560 66530 37570 66590
rect 37630 66530 37640 66590
rect 37560 66520 37640 66530
rect 39000 66600 39030 67050
rect 39000 66590 39080 66600
rect 39000 66530 39010 66590
rect 39070 66530 39080 66590
rect 39000 66520 39080 66530
rect 38850 66470 38910 66480
rect 38200 66440 38850 66450
rect 37580 66380 37640 66390
rect 38200 66380 38210 66440
rect 38270 66420 38850 66440
rect 38270 66380 38280 66420
rect 38850 66400 38910 66410
rect 39000 66380 39060 66390
rect 37780 66370 37860 66380
rect 38200 66370 38280 66380
rect 38620 66370 38700 66380
rect 37780 66360 37790 66370
rect 37640 66330 37790 66360
rect 37580 66310 37640 66320
rect 37780 66310 37790 66330
rect 37850 66310 37860 66370
rect 37780 66300 37860 66310
rect 38620 66310 38630 66370
rect 38690 66360 38700 66370
rect 38690 66330 39000 66360
rect 38690 66310 38700 66330
rect 39000 66310 39060 66320
rect 38620 66300 38700 66310
rect 38190 66280 38290 66290
rect 38190 66210 38210 66280
rect 38280 66210 38290 66280
rect 38190 66170 38290 66210
rect 38190 66100 38210 66170
rect 38280 66100 38290 66170
rect 38190 66080 38290 66100
rect 37560 66070 37640 66080
rect 39000 66070 39080 66080
rect 37560 66010 37570 66070
rect 37630 66050 37640 66070
rect 37780 66060 37860 66070
rect 37780 66050 37790 66060
rect 37630 66020 37790 66050
rect 37630 66010 37640 66020
rect 37560 66000 37640 66010
rect 37780 66000 37790 66020
rect 37850 66000 37860 66060
rect 38620 66060 38700 66070
rect 38620 66000 38630 66060
rect 38690 66050 38700 66060
rect 39000 66050 39010 66070
rect 38690 66020 39010 66050
rect 38690 66000 38700 66020
rect 39000 66010 39010 66020
rect 39070 66010 39080 66070
rect 39000 66000 39080 66010
rect 37780 65990 37860 66000
rect 38200 65990 38280 66000
rect 38620 65990 38700 66000
rect 38200 65930 38210 65990
rect 38270 65950 38280 65990
rect 38270 65940 38970 65950
rect 38270 65930 38910 65940
rect 38200 65920 38910 65930
rect 38910 65870 38970 65880
rect 38850 64760 38910 64770
rect 38200 64730 38850 64740
rect 37580 64670 37640 64680
rect 38200 64670 38210 64730
rect 38270 64710 38850 64730
rect 38270 64670 38280 64710
rect 38850 64690 38910 64700
rect 39000 64670 39060 64680
rect 37780 64660 37860 64670
rect 38200 64660 38280 64670
rect 38620 64660 38700 64670
rect 37780 64650 37790 64660
rect 37640 64620 37790 64650
rect 37580 64600 37640 64610
rect 37780 64600 37790 64620
rect 37850 64600 37860 64660
rect 37780 64590 37860 64600
rect 38620 64600 38630 64660
rect 38690 64650 38700 64660
rect 38690 64620 39000 64650
rect 38690 64600 38700 64620
rect 39000 64600 39060 64610
rect 38620 64590 38700 64600
rect 38190 64570 38290 64580
rect 38190 64500 38210 64570
rect 38280 64500 38290 64570
rect 38190 64460 38290 64500
rect 38190 64390 38210 64460
rect 38280 64390 38290 64460
rect 38190 64370 38290 64390
rect 37560 64360 37640 64370
rect 39000 64360 39080 64370
rect 37560 64300 37570 64360
rect 37630 64340 37640 64360
rect 37780 64350 37860 64360
rect 37780 64340 37790 64350
rect 37630 64310 37790 64340
rect 37630 64300 37640 64310
rect 37560 64290 37640 64300
rect 37780 64290 37790 64310
rect 37850 64290 37860 64350
rect 38620 64350 38700 64360
rect 38620 64290 38630 64350
rect 38690 64340 38700 64350
rect 39000 64340 39010 64360
rect 38690 64310 39010 64340
rect 38690 64290 38700 64310
rect 39000 64300 39010 64310
rect 39070 64300 39080 64360
rect 39000 64290 39080 64300
rect 37780 64280 37860 64290
rect 38200 64280 38280 64290
rect 38620 64280 38700 64290
rect 38200 64220 38210 64280
rect 38270 64240 38280 64280
rect 38270 64230 38970 64240
rect 38270 64220 38910 64230
rect 38200 64210 38910 64220
rect 38910 64160 38970 64170
rect 37440 63170 37520 63180
rect 37440 63110 37450 63170
rect 37510 63110 37520 63170
rect 37440 63100 37520 63110
rect 39120 63180 39150 67050
rect 39120 63170 39200 63180
rect 39120 63110 39130 63170
rect 39190 63110 39200 63170
rect 39120 63100 39200 63110
rect 38850 63050 38910 63060
rect 38200 63020 38850 63030
rect 37460 62960 37520 62970
rect 38200 62960 38210 63020
rect 38270 63000 38850 63020
rect 38270 62960 38280 63000
rect 38850 62980 38910 62990
rect 39120 62960 39180 62970
rect 37780 62950 37860 62960
rect 38200 62950 38280 62960
rect 38620 62950 38700 62960
rect 37780 62940 37790 62950
rect 37520 62910 37790 62940
rect 37460 62890 37520 62900
rect 37780 62890 37790 62910
rect 37850 62890 37860 62950
rect 37780 62880 37860 62890
rect 38620 62890 38630 62950
rect 38690 62940 38700 62950
rect 38690 62910 39120 62940
rect 38690 62890 38700 62910
rect 39120 62890 39180 62900
rect 38620 62880 38700 62890
rect 38190 62860 38290 62870
rect 38190 62790 38210 62860
rect 38280 62790 38290 62860
rect 38190 62750 38290 62790
rect 38190 62680 38210 62750
rect 38280 62680 38290 62750
rect 38190 62660 38290 62680
rect 37440 62650 37520 62660
rect 39120 62650 39200 62660
rect 37440 62590 37450 62650
rect 37510 62630 37520 62650
rect 37780 62640 37860 62650
rect 37780 62630 37790 62640
rect 37510 62600 37790 62630
rect 37510 62590 37520 62600
rect 37440 62580 37520 62590
rect 37780 62580 37790 62600
rect 37850 62580 37860 62640
rect 38620 62640 38700 62650
rect 38620 62580 38630 62640
rect 38690 62630 38700 62640
rect 39120 62630 39130 62650
rect 38690 62600 39130 62630
rect 38690 62580 38700 62600
rect 39120 62590 39130 62600
rect 39190 62590 39200 62650
rect 39120 62580 39200 62590
rect 37780 62570 37860 62580
rect 38200 62570 38280 62580
rect 38620 62570 38700 62580
rect 38200 62510 38210 62570
rect 38270 62530 38280 62570
rect 38270 62520 38970 62530
rect 38270 62510 38910 62520
rect 38200 62500 38910 62510
rect 38910 62450 38970 62460
rect 38850 61340 38910 61350
rect 38200 61310 38850 61320
rect 37460 61250 37520 61260
rect 38200 61250 38210 61310
rect 38270 61290 38850 61310
rect 38270 61250 38280 61290
rect 38850 61270 38910 61280
rect 39120 61250 39180 61260
rect 37780 61240 37860 61250
rect 38200 61240 38280 61250
rect 38620 61240 38700 61250
rect 37780 61230 37790 61240
rect 37520 61200 37790 61230
rect 37460 61180 37520 61190
rect 37780 61180 37790 61200
rect 37850 61180 37860 61240
rect 37780 61170 37860 61180
rect 38620 61180 38630 61240
rect 38690 61230 38700 61240
rect 38690 61200 39120 61230
rect 38690 61180 38700 61200
rect 39120 61180 39180 61190
rect 38620 61170 38700 61180
rect 38190 61150 38290 61160
rect 38190 61080 38210 61150
rect 38280 61080 38290 61150
rect 38190 61040 38290 61080
rect 38190 60970 38210 61040
rect 38280 60970 38290 61040
rect 38190 60950 38290 60970
rect 37440 60940 37520 60950
rect 39120 60940 39200 60950
rect 37440 60880 37450 60940
rect 37510 60920 37520 60940
rect 37780 60930 37860 60940
rect 37780 60920 37790 60930
rect 37510 60890 37790 60920
rect 37510 60880 37520 60890
rect 37440 60870 37520 60880
rect 37780 60870 37790 60890
rect 37850 60870 37860 60930
rect 38620 60930 38700 60940
rect 38620 60870 38630 60930
rect 38690 60920 38700 60930
rect 39120 60920 39130 60940
rect 38690 60890 39130 60920
rect 38690 60870 38700 60890
rect 39120 60880 39130 60890
rect 39190 60880 39200 60940
rect 39120 60870 39200 60880
rect 37780 60860 37860 60870
rect 38200 60860 38280 60870
rect 38620 60860 38700 60870
rect 38200 60800 38210 60860
rect 38270 60820 38280 60860
rect 38270 60810 38970 60820
rect 38270 60800 38910 60810
rect 38200 60790 38910 60800
rect 38910 60740 38970 60750
rect 37320 59750 37400 59760
rect 37320 59690 37330 59750
rect 37390 59690 37400 59750
rect 37320 59680 37400 59690
rect 39240 59760 39270 67050
rect 39240 59750 39320 59760
rect 39240 59690 39250 59750
rect 39310 59690 39320 59750
rect 39240 59680 39320 59690
rect 38850 59630 38910 59640
rect 38200 59600 38850 59610
rect 37340 59540 37400 59550
rect 38200 59540 38210 59600
rect 38270 59580 38850 59600
rect 38270 59540 38280 59580
rect 38850 59560 38910 59570
rect 39240 59540 39300 59550
rect 37780 59530 37860 59540
rect 38200 59530 38280 59540
rect 38620 59530 38700 59540
rect 37780 59520 37790 59530
rect 37400 59490 37790 59520
rect 37340 59470 37400 59480
rect 37780 59470 37790 59490
rect 37850 59470 37860 59530
rect 37780 59460 37860 59470
rect 38620 59470 38630 59530
rect 38690 59520 38700 59530
rect 38690 59490 39240 59520
rect 38690 59470 38700 59490
rect 39240 59470 39300 59480
rect 38620 59460 38700 59470
rect 38190 59440 38290 59450
rect 38190 59370 38210 59440
rect 38280 59370 38290 59440
rect 38190 59330 38290 59370
rect 38190 59260 38210 59330
rect 38280 59260 38290 59330
rect 38190 59240 38290 59260
rect 37320 59230 37400 59240
rect 39240 59230 39320 59240
rect 37320 59170 37330 59230
rect 37390 59210 37400 59230
rect 37780 59220 37860 59230
rect 37780 59210 37790 59220
rect 37390 59180 37790 59210
rect 37390 59170 37400 59180
rect 37320 59160 37400 59170
rect 37780 59160 37790 59180
rect 37850 59160 37860 59220
rect 38620 59220 38700 59230
rect 38620 59160 38630 59220
rect 38690 59210 38700 59220
rect 39240 59210 39250 59230
rect 38690 59180 39250 59210
rect 38690 59160 38700 59180
rect 39240 59170 39250 59180
rect 39310 59170 39320 59230
rect 39240 59160 39320 59170
rect 37780 59150 37860 59160
rect 38200 59150 38280 59160
rect 38620 59150 38700 59160
rect 38200 59090 38210 59150
rect 38270 59110 38280 59150
rect 38270 59100 38970 59110
rect 38270 59090 38910 59100
rect 38200 59080 38910 59090
rect 38910 59030 38970 59040
rect 37200 58040 37280 58050
rect 37200 57980 37210 58040
rect 37270 57980 37280 58040
rect 37200 57970 37280 57980
rect 39360 58050 39390 67050
rect 39360 58040 39440 58050
rect 39360 57980 39370 58040
rect 39430 57980 39440 58040
rect 39360 57970 39440 57980
rect 38850 57920 38910 57930
rect 38200 57890 38850 57900
rect 37220 57830 37280 57840
rect 38200 57830 38210 57890
rect 38270 57870 38850 57890
rect 38270 57830 38280 57870
rect 38850 57850 38910 57860
rect 39360 57830 39420 57840
rect 37780 57820 37860 57830
rect 38200 57820 38280 57830
rect 38620 57820 38700 57830
rect 37780 57810 37790 57820
rect 37280 57780 37790 57810
rect 37220 57760 37280 57770
rect 37780 57760 37790 57780
rect 37850 57760 37860 57820
rect 37780 57750 37860 57760
rect 38620 57760 38630 57820
rect 38690 57810 38700 57820
rect 38690 57780 39360 57810
rect 38690 57760 38700 57780
rect 39360 57760 39420 57770
rect 38620 57750 38700 57760
rect 38190 57730 38290 57740
rect 38190 57660 38210 57730
rect 38280 57660 38290 57730
rect 38190 57620 38290 57660
rect 38190 57550 38210 57620
rect 38280 57550 38290 57620
rect 38190 57530 38290 57550
rect 37200 57520 37280 57530
rect 39360 57520 39440 57530
rect 37200 57460 37210 57520
rect 37270 57500 37280 57520
rect 37780 57510 37860 57520
rect 37780 57500 37790 57510
rect 37270 57470 37790 57500
rect 37270 57460 37280 57470
rect 37200 57450 37280 57460
rect 37780 57450 37790 57470
rect 37850 57450 37860 57510
rect 38620 57510 38700 57520
rect 38620 57450 38630 57510
rect 38690 57500 38700 57510
rect 39360 57500 39370 57520
rect 38690 57470 39370 57500
rect 38690 57450 38700 57470
rect 39360 57460 39370 57470
rect 39430 57460 39440 57520
rect 39360 57450 39440 57460
rect 37780 57440 37860 57450
rect 38200 57440 38280 57450
rect 38620 57440 38700 57450
rect 38200 57380 38210 57440
rect 38270 57400 38280 57440
rect 38270 57390 38970 57400
rect 38270 57380 38910 57390
rect 38200 57370 38910 57380
rect 38910 57320 38970 57330
rect 37080 56330 37160 56340
rect 37080 56270 37090 56330
rect 37150 56270 37160 56330
rect 37080 56260 37160 56270
rect 39480 56340 39510 67050
rect 39480 56330 39560 56340
rect 39480 56270 39490 56330
rect 39550 56270 39560 56330
rect 39480 56260 39560 56270
rect 38850 56210 38910 56220
rect 38200 56180 38850 56190
rect 37100 56120 37160 56130
rect 38200 56120 38210 56180
rect 38270 56160 38850 56180
rect 38270 56120 38280 56160
rect 38850 56140 38910 56150
rect 39480 56120 39540 56130
rect 37780 56110 37860 56120
rect 38200 56110 38280 56120
rect 38620 56110 38700 56120
rect 37780 56100 37790 56110
rect 37160 56070 37790 56100
rect 37100 56050 37160 56060
rect 37780 56050 37790 56070
rect 37850 56050 37860 56110
rect 37780 56040 37860 56050
rect 38620 56050 38630 56110
rect 38690 56100 38700 56110
rect 38690 56070 39480 56100
rect 38690 56050 38700 56070
rect 39480 56050 39540 56060
rect 38620 56040 38700 56050
rect 38190 56020 38290 56030
rect 38190 55950 38210 56020
rect 38280 55950 38290 56020
rect 38190 55910 38290 55950
rect 38190 55840 38210 55910
rect 38280 55840 38290 55910
rect 38190 55820 38290 55840
rect 37080 55810 37160 55820
rect 39480 55810 39560 55820
rect 37080 55750 37090 55810
rect 37150 55790 37160 55810
rect 37780 55800 37860 55810
rect 37780 55790 37790 55800
rect 37150 55760 37790 55790
rect 37150 55750 37160 55760
rect 37080 55740 37160 55750
rect 37780 55740 37790 55760
rect 37850 55740 37860 55800
rect 38620 55800 38700 55810
rect 38620 55740 38630 55800
rect 38690 55790 38700 55800
rect 39480 55790 39490 55810
rect 38690 55760 39490 55790
rect 38690 55740 38700 55760
rect 39480 55750 39490 55760
rect 39550 55750 39560 55810
rect 39480 55740 39560 55750
rect 37780 55730 37860 55740
rect 38200 55730 38280 55740
rect 38620 55730 38700 55740
rect 38200 55670 38210 55730
rect 38270 55690 38280 55730
rect 38270 55680 38970 55690
rect 38270 55670 38910 55680
rect 38200 55660 38910 55670
rect 38910 55610 38970 55620
rect 36960 54610 37040 54620
rect 36960 54550 36970 54610
rect 37030 54550 37040 54610
rect 39600 54670 39630 67050
rect 39600 54660 39680 54670
rect 39600 54600 39610 54660
rect 39670 54600 39680 54660
rect 39600 54590 39680 54600
rect 36960 54540 37040 54550
rect 38850 54500 38910 54510
rect 33860 54430 33920 54440
rect 36800 54440 36920 54470
rect 38200 54470 38850 54480
rect 34610 54410 34670 54420
rect 32790 54400 32870 54410
rect 33210 54400 33290 54410
rect 33630 54400 33710 54410
rect 32790 54390 32800 54400
rect 32050 54360 32800 54390
rect 31990 54340 32050 54350
rect 32790 54340 32800 54360
rect 32860 54340 32870 54400
rect 28640 54330 28720 54340
rect 32790 54330 32870 54340
rect 33630 54340 33640 54400
rect 33700 54390 33710 54400
rect 33700 54360 34610 54390
rect 33700 54340 33710 54360
rect 34610 54340 34670 54350
rect 33630 54330 33710 54340
rect 3260 54310 3360 54320
rect 3260 54240 3280 54310
rect 3350 54240 3360 54310
rect 3260 54200 3360 54240
rect 3260 54130 3280 54200
rect 3350 54130 3360 54200
rect 3260 54110 3360 54130
rect 8250 54310 8350 54320
rect 8250 54240 8270 54310
rect 8340 54240 8350 54310
rect 8250 54200 8350 54240
rect 8250 54130 8270 54200
rect 8340 54130 8350 54200
rect 8250 54110 8350 54130
rect 13240 54310 13340 54320
rect 13240 54240 13260 54310
rect 13330 54240 13340 54310
rect 13240 54200 13340 54240
rect 13240 54130 13260 54200
rect 13330 54130 13340 54200
rect 13240 54110 13340 54130
rect 18230 54310 18330 54320
rect 18230 54240 18250 54310
rect 18320 54240 18330 54310
rect 18230 54200 18330 54240
rect 18230 54130 18250 54200
rect 18320 54130 18330 54200
rect 18230 54110 18330 54130
rect 23220 54310 23320 54320
rect 23220 54240 23240 54310
rect 23310 54240 23320 54310
rect 23220 54200 23320 54240
rect 23220 54130 23240 54200
rect 23310 54130 23320 54200
rect 23220 54110 23320 54130
rect 28210 54310 28310 54320
rect 28210 54240 28230 54310
rect 28300 54240 28310 54310
rect 28210 54200 28310 54240
rect 28210 54130 28230 54200
rect 28300 54130 28310 54200
rect 28210 54110 28310 54130
rect 33200 54310 33300 54320
rect 33200 54240 33220 54310
rect 33290 54240 33300 54310
rect 36800 54300 36830 54440
rect 38200 54410 38210 54470
rect 38270 54450 38850 54470
rect 38270 54410 38280 54450
rect 39720 54470 39750 67050
rect 41880 54470 41910 67050
rect 42000 54620 42030 67050
rect 42120 56340 42150 67050
rect 42240 58050 42270 67050
rect 42360 59760 42390 67050
rect 42480 63180 42510 67050
rect 42600 66600 42630 67050
rect 42550 66590 42630 66600
rect 42550 66530 42560 66590
rect 42620 66530 42630 66590
rect 42550 66520 42630 66530
rect 43990 66600 44020 67050
rect 43990 66590 44070 66600
rect 43990 66530 44000 66590
rect 44060 66530 44070 66590
rect 43990 66520 44070 66530
rect 43840 66470 43900 66480
rect 43190 66440 43840 66450
rect 42570 66380 42630 66390
rect 43190 66380 43200 66440
rect 43260 66420 43840 66440
rect 43260 66380 43270 66420
rect 43840 66400 43900 66410
rect 43990 66380 44050 66390
rect 42770 66370 42850 66380
rect 43190 66370 43270 66380
rect 43610 66370 43690 66380
rect 42770 66360 42780 66370
rect 42630 66330 42780 66360
rect 42570 66310 42630 66320
rect 42770 66310 42780 66330
rect 42840 66310 42850 66370
rect 42770 66300 42850 66310
rect 43610 66310 43620 66370
rect 43680 66360 43690 66370
rect 43680 66330 43990 66360
rect 43680 66310 43690 66330
rect 43990 66310 44050 66320
rect 43610 66300 43690 66310
rect 43180 66280 43280 66290
rect 43180 66210 43200 66280
rect 43270 66210 43280 66280
rect 43180 66170 43280 66210
rect 43180 66100 43200 66170
rect 43270 66100 43280 66170
rect 43180 66080 43280 66100
rect 42550 66070 42630 66080
rect 43990 66070 44070 66080
rect 42550 66010 42560 66070
rect 42620 66050 42630 66070
rect 42770 66060 42850 66070
rect 42770 66050 42780 66060
rect 42620 66020 42780 66050
rect 42620 66010 42630 66020
rect 42550 66000 42630 66010
rect 42770 66000 42780 66020
rect 42840 66000 42850 66060
rect 43610 66060 43690 66070
rect 43610 66000 43620 66060
rect 43680 66050 43690 66060
rect 43990 66050 44000 66070
rect 43680 66020 44000 66050
rect 43680 66000 43690 66020
rect 43990 66010 44000 66020
rect 44060 66010 44070 66070
rect 43990 66000 44070 66010
rect 42770 65990 42850 66000
rect 43190 65990 43270 66000
rect 43610 65990 43690 66000
rect 43190 65930 43200 65990
rect 43260 65950 43270 65990
rect 43260 65940 43960 65950
rect 43260 65930 43900 65940
rect 43190 65920 43900 65930
rect 43900 65870 43960 65880
rect 43840 64760 43900 64770
rect 43190 64730 43840 64740
rect 42570 64670 42630 64680
rect 43190 64670 43200 64730
rect 43260 64710 43840 64730
rect 43260 64670 43270 64710
rect 43840 64690 43900 64700
rect 43990 64670 44050 64680
rect 42770 64660 42850 64670
rect 43190 64660 43270 64670
rect 43610 64660 43690 64670
rect 42770 64650 42780 64660
rect 42630 64620 42780 64650
rect 42570 64600 42630 64610
rect 42770 64600 42780 64620
rect 42840 64600 42850 64660
rect 42770 64590 42850 64600
rect 43610 64600 43620 64660
rect 43680 64650 43690 64660
rect 43680 64620 43990 64650
rect 43680 64600 43690 64620
rect 43990 64600 44050 64610
rect 43610 64590 43690 64600
rect 43180 64570 43280 64580
rect 43180 64500 43200 64570
rect 43270 64500 43280 64570
rect 43180 64460 43280 64500
rect 43180 64390 43200 64460
rect 43270 64390 43280 64460
rect 43180 64370 43280 64390
rect 42550 64360 42630 64370
rect 43990 64360 44070 64370
rect 42550 64300 42560 64360
rect 42620 64340 42630 64360
rect 42770 64350 42850 64360
rect 42770 64340 42780 64350
rect 42620 64310 42780 64340
rect 42620 64300 42630 64310
rect 42550 64290 42630 64300
rect 42770 64290 42780 64310
rect 42840 64290 42850 64350
rect 43610 64350 43690 64360
rect 43610 64290 43620 64350
rect 43680 64340 43690 64350
rect 43990 64340 44000 64360
rect 43680 64310 44000 64340
rect 43680 64290 43690 64310
rect 43990 64300 44000 64310
rect 44060 64300 44070 64360
rect 43990 64290 44070 64300
rect 42770 64280 42850 64290
rect 43190 64280 43270 64290
rect 43610 64280 43690 64290
rect 43190 64220 43200 64280
rect 43260 64240 43270 64280
rect 43260 64230 43960 64240
rect 43260 64220 43900 64230
rect 43190 64210 43900 64220
rect 43900 64160 43960 64170
rect 42430 63170 42510 63180
rect 42430 63110 42440 63170
rect 42500 63110 42510 63170
rect 42430 63100 42510 63110
rect 44110 63180 44140 67050
rect 44110 63170 44190 63180
rect 44110 63110 44120 63170
rect 44180 63110 44190 63170
rect 44110 63100 44190 63110
rect 43840 63050 43900 63060
rect 43190 63020 43840 63030
rect 42450 62960 42510 62970
rect 43190 62960 43200 63020
rect 43260 63000 43840 63020
rect 43260 62960 43270 63000
rect 43840 62980 43900 62990
rect 44110 62960 44170 62970
rect 42770 62950 42850 62960
rect 43190 62950 43270 62960
rect 43610 62950 43690 62960
rect 42770 62940 42780 62950
rect 42510 62910 42780 62940
rect 42450 62890 42510 62900
rect 42770 62890 42780 62910
rect 42840 62890 42850 62950
rect 42770 62880 42850 62890
rect 43610 62890 43620 62950
rect 43680 62940 43690 62950
rect 43680 62910 44110 62940
rect 43680 62890 43690 62910
rect 44110 62890 44170 62900
rect 43610 62880 43690 62890
rect 43180 62860 43280 62870
rect 43180 62790 43200 62860
rect 43270 62790 43280 62860
rect 43180 62750 43280 62790
rect 43180 62680 43200 62750
rect 43270 62680 43280 62750
rect 43180 62660 43280 62680
rect 42430 62650 42510 62660
rect 44110 62650 44190 62660
rect 42430 62590 42440 62650
rect 42500 62630 42510 62650
rect 42770 62640 42850 62650
rect 42770 62630 42780 62640
rect 42500 62600 42780 62630
rect 42500 62590 42510 62600
rect 42430 62580 42510 62590
rect 42770 62580 42780 62600
rect 42840 62580 42850 62640
rect 43610 62640 43690 62650
rect 43610 62580 43620 62640
rect 43680 62630 43690 62640
rect 44110 62630 44120 62650
rect 43680 62600 44120 62630
rect 43680 62580 43690 62600
rect 44110 62590 44120 62600
rect 44180 62590 44190 62650
rect 44110 62580 44190 62590
rect 42770 62570 42850 62580
rect 43190 62570 43270 62580
rect 43610 62570 43690 62580
rect 43190 62510 43200 62570
rect 43260 62530 43270 62570
rect 43260 62520 43960 62530
rect 43260 62510 43900 62520
rect 43190 62500 43900 62510
rect 43900 62450 43960 62460
rect 43840 61340 43900 61350
rect 43190 61310 43840 61320
rect 42450 61250 42510 61260
rect 43190 61250 43200 61310
rect 43260 61290 43840 61310
rect 43260 61250 43270 61290
rect 43840 61270 43900 61280
rect 44110 61250 44170 61260
rect 42770 61240 42850 61250
rect 43190 61240 43270 61250
rect 43610 61240 43690 61250
rect 42770 61230 42780 61240
rect 42510 61200 42780 61230
rect 42450 61180 42510 61190
rect 42770 61180 42780 61200
rect 42840 61180 42850 61240
rect 42770 61170 42850 61180
rect 43610 61180 43620 61240
rect 43680 61230 43690 61240
rect 43680 61200 44110 61230
rect 43680 61180 43690 61200
rect 44110 61180 44170 61190
rect 43610 61170 43690 61180
rect 43180 61150 43280 61160
rect 43180 61080 43200 61150
rect 43270 61080 43280 61150
rect 43180 61040 43280 61080
rect 43180 60970 43200 61040
rect 43270 60970 43280 61040
rect 43180 60950 43280 60970
rect 42430 60940 42510 60950
rect 44110 60940 44190 60950
rect 42430 60880 42440 60940
rect 42500 60920 42510 60940
rect 42770 60930 42850 60940
rect 42770 60920 42780 60930
rect 42500 60890 42780 60920
rect 42500 60880 42510 60890
rect 42430 60870 42510 60880
rect 42770 60870 42780 60890
rect 42840 60870 42850 60930
rect 43610 60930 43690 60940
rect 43610 60870 43620 60930
rect 43680 60920 43690 60930
rect 44110 60920 44120 60940
rect 43680 60890 44120 60920
rect 43680 60870 43690 60890
rect 44110 60880 44120 60890
rect 44180 60880 44190 60940
rect 44110 60870 44190 60880
rect 42770 60860 42850 60870
rect 43190 60860 43270 60870
rect 43610 60860 43690 60870
rect 43190 60800 43200 60860
rect 43260 60820 43270 60860
rect 43260 60810 43960 60820
rect 43260 60800 43900 60810
rect 43190 60790 43900 60800
rect 43900 60740 43960 60750
rect 42310 59750 42390 59760
rect 42310 59690 42320 59750
rect 42380 59690 42390 59750
rect 42310 59680 42390 59690
rect 44230 59760 44260 67050
rect 44230 59750 44310 59760
rect 44230 59690 44240 59750
rect 44300 59690 44310 59750
rect 44230 59680 44310 59690
rect 43840 59630 43900 59640
rect 43190 59600 43840 59610
rect 42330 59540 42390 59550
rect 43190 59540 43200 59600
rect 43260 59580 43840 59600
rect 43260 59540 43270 59580
rect 43840 59560 43900 59570
rect 44230 59540 44290 59550
rect 42770 59530 42850 59540
rect 43190 59530 43270 59540
rect 43610 59530 43690 59540
rect 42770 59520 42780 59530
rect 42390 59490 42780 59520
rect 42330 59470 42390 59480
rect 42770 59470 42780 59490
rect 42840 59470 42850 59530
rect 42770 59460 42850 59470
rect 43610 59470 43620 59530
rect 43680 59520 43690 59530
rect 43680 59490 44230 59520
rect 43680 59470 43690 59490
rect 44230 59470 44290 59480
rect 43610 59460 43690 59470
rect 43180 59440 43280 59450
rect 43180 59370 43200 59440
rect 43270 59370 43280 59440
rect 43180 59330 43280 59370
rect 43180 59260 43200 59330
rect 43270 59260 43280 59330
rect 43180 59240 43280 59260
rect 42310 59230 42390 59240
rect 44230 59230 44310 59240
rect 42310 59170 42320 59230
rect 42380 59210 42390 59230
rect 42770 59220 42850 59230
rect 42770 59210 42780 59220
rect 42380 59180 42780 59210
rect 42380 59170 42390 59180
rect 42310 59160 42390 59170
rect 42770 59160 42780 59180
rect 42840 59160 42850 59220
rect 43610 59220 43690 59230
rect 43610 59160 43620 59220
rect 43680 59210 43690 59220
rect 44230 59210 44240 59230
rect 43680 59180 44240 59210
rect 43680 59160 43690 59180
rect 44230 59170 44240 59180
rect 44300 59170 44310 59230
rect 44230 59160 44310 59170
rect 42770 59150 42850 59160
rect 43190 59150 43270 59160
rect 43610 59150 43690 59160
rect 43190 59090 43200 59150
rect 43260 59110 43270 59150
rect 43260 59100 43960 59110
rect 43260 59090 43900 59100
rect 43190 59080 43900 59090
rect 43900 59030 43960 59040
rect 42190 58040 42270 58050
rect 42190 57980 42200 58040
rect 42260 57980 42270 58040
rect 42190 57970 42270 57980
rect 44350 58050 44380 67050
rect 44350 58040 44430 58050
rect 44350 57980 44360 58040
rect 44420 57980 44430 58040
rect 44350 57970 44430 57980
rect 43840 57920 43900 57930
rect 43190 57890 43840 57900
rect 42210 57830 42270 57840
rect 43190 57830 43200 57890
rect 43260 57870 43840 57890
rect 43260 57830 43270 57870
rect 43840 57850 43900 57860
rect 44350 57830 44410 57840
rect 42770 57820 42850 57830
rect 43190 57820 43270 57830
rect 43610 57820 43690 57830
rect 42770 57810 42780 57820
rect 42270 57780 42780 57810
rect 42210 57760 42270 57770
rect 42770 57760 42780 57780
rect 42840 57760 42850 57820
rect 42770 57750 42850 57760
rect 43610 57760 43620 57820
rect 43680 57810 43690 57820
rect 43680 57780 44350 57810
rect 43680 57760 43690 57780
rect 44350 57760 44410 57770
rect 43610 57750 43690 57760
rect 43180 57730 43280 57740
rect 43180 57660 43200 57730
rect 43270 57660 43280 57730
rect 43180 57620 43280 57660
rect 43180 57550 43200 57620
rect 43270 57550 43280 57620
rect 43180 57530 43280 57550
rect 42190 57520 42270 57530
rect 44350 57520 44430 57530
rect 42190 57460 42200 57520
rect 42260 57500 42270 57520
rect 42770 57510 42850 57520
rect 42770 57500 42780 57510
rect 42260 57470 42780 57500
rect 42260 57460 42270 57470
rect 42190 57450 42270 57460
rect 42770 57450 42780 57470
rect 42840 57450 42850 57510
rect 43610 57510 43690 57520
rect 43610 57450 43620 57510
rect 43680 57500 43690 57510
rect 44350 57500 44360 57520
rect 43680 57470 44360 57500
rect 43680 57450 43690 57470
rect 44350 57460 44360 57470
rect 44420 57460 44430 57520
rect 44350 57450 44430 57460
rect 42770 57440 42850 57450
rect 43190 57440 43270 57450
rect 43610 57440 43690 57450
rect 43190 57380 43200 57440
rect 43260 57400 43270 57440
rect 43260 57390 43960 57400
rect 43260 57380 43900 57390
rect 43190 57370 43900 57380
rect 43900 57320 43960 57330
rect 42070 56330 42150 56340
rect 42070 56270 42080 56330
rect 42140 56270 42150 56330
rect 42070 56260 42150 56270
rect 44470 56340 44500 67050
rect 44470 56330 44550 56340
rect 44470 56270 44480 56330
rect 44540 56270 44550 56330
rect 44470 56260 44550 56270
rect 43840 56210 43900 56220
rect 43190 56180 43840 56190
rect 42090 56120 42150 56130
rect 43190 56120 43200 56180
rect 43260 56160 43840 56180
rect 43260 56120 43270 56160
rect 43840 56140 43900 56150
rect 44470 56120 44530 56130
rect 42770 56110 42850 56120
rect 43190 56110 43270 56120
rect 43610 56110 43690 56120
rect 42770 56100 42780 56110
rect 42150 56070 42780 56100
rect 42090 56050 42150 56060
rect 42770 56050 42780 56070
rect 42840 56050 42850 56110
rect 42770 56040 42850 56050
rect 43610 56050 43620 56110
rect 43680 56100 43690 56110
rect 43680 56070 44470 56100
rect 43680 56050 43690 56070
rect 44470 56050 44530 56060
rect 43610 56040 43690 56050
rect 43180 56020 43280 56030
rect 43180 55950 43200 56020
rect 43270 55950 43280 56020
rect 43180 55910 43280 55950
rect 43180 55840 43200 55910
rect 43270 55840 43280 55910
rect 43180 55820 43280 55840
rect 42070 55810 42150 55820
rect 44470 55810 44550 55820
rect 42070 55750 42080 55810
rect 42140 55790 42150 55810
rect 42770 55800 42850 55810
rect 42770 55790 42780 55800
rect 42140 55760 42780 55790
rect 42140 55750 42150 55760
rect 42070 55740 42150 55750
rect 42770 55740 42780 55760
rect 42840 55740 42850 55800
rect 43610 55800 43690 55810
rect 43610 55740 43620 55800
rect 43680 55790 43690 55800
rect 44470 55790 44480 55810
rect 43680 55760 44480 55790
rect 43680 55740 43690 55760
rect 44470 55750 44480 55760
rect 44540 55750 44550 55810
rect 44470 55740 44550 55750
rect 42770 55730 42850 55740
rect 43190 55730 43270 55740
rect 43610 55730 43690 55740
rect 43190 55670 43200 55730
rect 43260 55690 43270 55730
rect 43260 55680 43960 55690
rect 43260 55670 43900 55680
rect 43190 55660 43900 55670
rect 43900 55610 43960 55620
rect 41950 54610 42030 54620
rect 41950 54550 41960 54610
rect 42020 54550 42030 54610
rect 44590 54670 44620 67050
rect 44590 54660 44670 54670
rect 44590 54600 44600 54660
rect 44660 54600 44670 54660
rect 44590 54590 44670 54600
rect 41950 54540 42030 54550
rect 43840 54500 43900 54510
rect 39720 54440 39840 54470
rect 38850 54430 38910 54440
rect 36860 54400 36920 54410
rect 37780 54400 37860 54410
rect 38200 54400 38280 54410
rect 38620 54400 38700 54410
rect 37780 54390 37790 54400
rect 36920 54360 37790 54390
rect 36860 54330 36920 54340
rect 37780 54340 37790 54360
rect 37850 54340 37860 54400
rect 37780 54330 37860 54340
rect 38620 54340 38630 54400
rect 38690 54390 38700 54400
rect 39720 54400 39780 54410
rect 38690 54360 39720 54390
rect 38690 54340 38700 54360
rect 38620 54330 38700 54340
rect 39720 54330 39780 54340
rect 38190 54310 38290 54320
rect 36800 54270 36920 54300
rect 33200 54200 33300 54240
rect 33200 54130 33220 54200
rect 33290 54130 33300 54200
rect 33200 54110 33300 54130
rect 2630 54090 2710 54100
rect 2630 54030 2640 54090
rect 2700 54080 2710 54090
rect 2850 54090 2930 54100
rect 2850 54080 2860 54090
rect 2700 54050 2860 54080
rect 2700 54030 2710 54050
rect 2630 54020 2710 54030
rect 2850 54030 2860 54050
rect 2920 54030 2930 54090
rect 3690 54090 3770 54100
rect 3690 54030 3700 54090
rect 3760 54080 3770 54090
rect 4070 54090 4150 54100
rect 4070 54080 4080 54090
rect 3760 54050 4080 54080
rect 3760 54030 3770 54050
rect 2850 54020 2930 54030
rect 3270 54020 3350 54030
rect 3690 54020 3770 54030
rect 4070 54030 4080 54050
rect 4140 54030 4150 54090
rect 4070 54020 4150 54030
rect 7620 54090 7700 54100
rect 7620 54030 7630 54090
rect 7690 54080 7700 54090
rect 7840 54090 7920 54100
rect 7840 54080 7850 54090
rect 7690 54050 7850 54080
rect 7690 54030 7700 54050
rect 7620 54020 7700 54030
rect 7840 54030 7850 54050
rect 7910 54030 7920 54090
rect 8680 54090 8760 54100
rect 8680 54030 8690 54090
rect 8750 54080 8760 54090
rect 9060 54090 9140 54100
rect 9060 54080 9070 54090
rect 8750 54050 9070 54080
rect 8750 54030 8760 54050
rect 7840 54020 7920 54030
rect 8260 54020 8340 54030
rect 8680 54020 8760 54030
rect 9060 54030 9070 54050
rect 9130 54030 9140 54090
rect 9060 54020 9140 54030
rect 12490 54090 12570 54100
rect 12490 54030 12500 54090
rect 12560 54080 12570 54090
rect 12830 54090 12910 54100
rect 12830 54080 12840 54090
rect 12560 54050 12840 54080
rect 12560 54030 12570 54050
rect 12490 54020 12570 54030
rect 12830 54030 12840 54050
rect 12900 54030 12910 54090
rect 13670 54090 13750 54100
rect 13670 54030 13680 54090
rect 13740 54080 13750 54090
rect 14170 54090 14250 54100
rect 14170 54080 14180 54090
rect 13740 54050 14180 54080
rect 13740 54030 13750 54050
rect 12830 54020 12910 54030
rect 13250 54020 13330 54030
rect 13670 54020 13750 54030
rect 14170 54030 14180 54050
rect 14240 54030 14250 54090
rect 14170 54020 14250 54030
rect 17480 54090 17560 54100
rect 17480 54030 17490 54090
rect 17550 54080 17560 54090
rect 17820 54090 17900 54100
rect 17820 54080 17830 54090
rect 17550 54050 17830 54080
rect 17550 54030 17560 54050
rect 17480 54020 17560 54030
rect 17820 54030 17830 54050
rect 17890 54030 17900 54090
rect 18660 54090 18740 54100
rect 18660 54030 18670 54090
rect 18730 54080 18740 54090
rect 19160 54090 19240 54100
rect 19160 54080 19170 54090
rect 18730 54050 19170 54080
rect 18730 54030 18740 54050
rect 17820 54020 17900 54030
rect 18240 54020 18320 54030
rect 18660 54020 18740 54030
rect 19160 54030 19170 54050
rect 19230 54030 19240 54090
rect 19160 54020 19240 54030
rect 22230 54090 22310 54100
rect 22230 54030 22240 54090
rect 22300 54080 22310 54090
rect 22810 54090 22890 54100
rect 22810 54080 22820 54090
rect 22300 54050 22820 54080
rect 22300 54030 22310 54050
rect 22230 54020 22310 54030
rect 22810 54030 22820 54050
rect 22880 54030 22890 54090
rect 23650 54090 23730 54100
rect 23650 54030 23660 54090
rect 23720 54080 23730 54090
rect 24390 54090 24470 54100
rect 24390 54080 24400 54090
rect 23720 54050 24400 54080
rect 23720 54030 23730 54050
rect 22810 54020 22890 54030
rect 23230 54020 23310 54030
rect 23650 54020 23730 54030
rect 24390 54030 24400 54050
rect 24460 54030 24470 54090
rect 24390 54020 24470 54030
rect 27220 54090 27300 54100
rect 27220 54030 27230 54090
rect 27290 54080 27300 54090
rect 27800 54090 27880 54100
rect 27800 54080 27810 54090
rect 27290 54050 27810 54080
rect 27290 54030 27300 54050
rect 27220 54020 27300 54030
rect 27800 54030 27810 54050
rect 27870 54030 27880 54090
rect 28640 54090 28720 54100
rect 28640 54030 28650 54090
rect 28710 54080 28720 54090
rect 29380 54090 29460 54100
rect 29380 54080 29390 54090
rect 28710 54050 29390 54080
rect 28710 54030 28720 54050
rect 27800 54020 27880 54030
rect 28220 54020 28300 54030
rect 28640 54020 28720 54030
rect 29380 54030 29390 54050
rect 29450 54030 29460 54090
rect 29380 54020 29460 54030
rect 31970 54090 32050 54100
rect 31970 54030 31980 54090
rect 32040 54080 32050 54090
rect 32790 54090 32870 54100
rect 32790 54080 32800 54090
rect 32040 54050 32800 54080
rect 32040 54030 32050 54050
rect 31970 54020 32050 54030
rect 32790 54030 32800 54050
rect 32860 54030 32870 54090
rect 33630 54090 33710 54100
rect 33630 54030 33640 54090
rect 33700 54080 33710 54090
rect 34610 54090 34690 54100
rect 34610 54080 34620 54090
rect 33700 54050 34620 54080
rect 33700 54030 33710 54050
rect 32790 54020 32870 54030
rect 33210 54020 33290 54030
rect 33630 54020 33710 54030
rect 34610 54030 34620 54050
rect 34680 54030 34690 54090
rect 34610 54020 34690 54030
rect 36890 54080 36920 54270
rect 38190 54240 38210 54310
rect 38280 54240 38290 54310
rect 39810 54300 39840 54440
rect 38190 54200 38290 54240
rect 38190 54130 38210 54200
rect 38280 54130 38290 54200
rect 38190 54110 38290 54130
rect 39720 54270 39840 54300
rect 41790 54440 41910 54470
rect 43190 54470 43840 54480
rect 41790 54300 41820 54440
rect 43190 54410 43200 54470
rect 43260 54450 43840 54470
rect 43260 54410 43270 54450
rect 44710 54470 44740 67050
rect 46990 54620 47020 67050
rect 47110 56330 47140 67050
rect 47230 58040 47260 67050
rect 47350 59750 47380 67050
rect 47470 63170 47500 67050
rect 47590 66590 47620 67050
rect 47540 66580 47620 66590
rect 47540 66520 47550 66580
rect 47610 66520 47620 66580
rect 47540 66510 47620 66520
rect 48980 66590 49010 67050
rect 48980 66580 49060 66590
rect 48980 66520 48990 66580
rect 49050 66520 49060 66580
rect 48980 66510 49060 66520
rect 48830 66470 48890 66480
rect 48180 66440 48830 66450
rect 47560 66380 47620 66390
rect 48180 66380 48190 66440
rect 48250 66420 48830 66440
rect 48250 66380 48260 66420
rect 48830 66400 48890 66410
rect 48980 66380 49040 66390
rect 47760 66370 47840 66380
rect 48180 66370 48260 66380
rect 48600 66370 48680 66380
rect 47760 66360 47770 66370
rect 47620 66330 47770 66360
rect 47560 66310 47620 66320
rect 47760 66310 47770 66330
rect 47830 66310 47840 66370
rect 47760 66300 47840 66310
rect 48600 66310 48610 66370
rect 48670 66360 48680 66370
rect 48670 66330 48980 66360
rect 48670 66310 48680 66330
rect 48980 66310 49040 66320
rect 48600 66300 48680 66310
rect 48170 66280 48270 66290
rect 48170 66210 48190 66280
rect 48260 66210 48270 66280
rect 48170 66170 48270 66210
rect 48170 66100 48190 66170
rect 48260 66100 48270 66170
rect 48170 66080 48270 66100
rect 47540 66060 47620 66070
rect 47540 66000 47550 66060
rect 47610 66050 47620 66060
rect 47760 66060 47840 66070
rect 47760 66050 47770 66060
rect 47610 66020 47770 66050
rect 47610 66000 47620 66020
rect 47540 65990 47620 66000
rect 47760 66000 47770 66020
rect 47830 66000 47840 66060
rect 48600 66060 48680 66070
rect 48600 66000 48610 66060
rect 48670 66050 48680 66060
rect 48980 66060 49060 66070
rect 48980 66050 48990 66060
rect 48670 66020 48990 66050
rect 48670 66000 48680 66020
rect 47760 65990 47840 66000
rect 48180 65990 48260 66000
rect 48600 65990 48680 66000
rect 48980 66000 48990 66020
rect 49050 66000 49060 66060
rect 48980 65990 49060 66000
rect 48180 65930 48190 65990
rect 48250 65950 48260 65990
rect 48250 65940 48950 65950
rect 48250 65930 48890 65940
rect 48180 65920 48890 65930
rect 48890 65870 48950 65880
rect 48830 64760 48890 64770
rect 48180 64730 48830 64740
rect 47560 64670 47620 64680
rect 48180 64670 48190 64730
rect 48250 64710 48830 64730
rect 48250 64670 48260 64710
rect 48830 64690 48890 64700
rect 48980 64670 49040 64680
rect 47760 64660 47840 64670
rect 48180 64660 48260 64670
rect 48600 64660 48680 64670
rect 47760 64650 47770 64660
rect 47620 64620 47770 64650
rect 47560 64600 47620 64610
rect 47760 64600 47770 64620
rect 47830 64600 47840 64660
rect 47760 64590 47840 64600
rect 48600 64600 48610 64660
rect 48670 64650 48680 64660
rect 48670 64620 48980 64650
rect 48670 64600 48680 64620
rect 48980 64600 49040 64610
rect 48600 64590 48680 64600
rect 48170 64570 48270 64580
rect 48170 64500 48190 64570
rect 48260 64500 48270 64570
rect 48170 64460 48270 64500
rect 48170 64390 48190 64460
rect 48260 64390 48270 64460
rect 48170 64370 48270 64390
rect 47540 64350 47620 64360
rect 47540 64290 47550 64350
rect 47610 64340 47620 64350
rect 47760 64350 47840 64360
rect 47760 64340 47770 64350
rect 47610 64310 47770 64340
rect 47610 64290 47620 64310
rect 47540 64280 47620 64290
rect 47760 64290 47770 64310
rect 47830 64290 47840 64350
rect 48600 64350 48680 64360
rect 48600 64290 48610 64350
rect 48670 64340 48680 64350
rect 48980 64350 49060 64360
rect 48980 64340 48990 64350
rect 48670 64310 48990 64340
rect 48670 64290 48680 64310
rect 47760 64280 47840 64290
rect 48180 64280 48260 64290
rect 48600 64280 48680 64290
rect 48980 64290 48990 64310
rect 49050 64290 49060 64350
rect 48980 64280 49060 64290
rect 48180 64220 48190 64280
rect 48250 64240 48260 64280
rect 48250 64230 48950 64240
rect 48250 64220 48890 64230
rect 48180 64210 48890 64220
rect 48890 64160 48950 64170
rect 47420 63160 47500 63170
rect 47420 63100 47430 63160
rect 47490 63100 47500 63160
rect 47420 63090 47500 63100
rect 49100 63170 49130 67050
rect 49100 63160 49180 63170
rect 49100 63100 49110 63160
rect 49170 63100 49180 63160
rect 49100 63090 49180 63100
rect 48830 63050 48890 63060
rect 48180 63020 48830 63030
rect 47440 62960 47500 62970
rect 48180 62960 48190 63020
rect 48250 63000 48830 63020
rect 48250 62960 48260 63000
rect 48830 62980 48890 62990
rect 49100 62960 49160 62970
rect 47760 62950 47840 62960
rect 48180 62950 48260 62960
rect 48600 62950 48680 62960
rect 47760 62940 47770 62950
rect 47500 62910 47770 62940
rect 47440 62890 47500 62900
rect 47760 62890 47770 62910
rect 47830 62890 47840 62950
rect 47760 62880 47840 62890
rect 48600 62890 48610 62950
rect 48670 62940 48680 62950
rect 48670 62910 49100 62940
rect 48670 62890 48680 62910
rect 49100 62890 49160 62900
rect 48600 62880 48680 62890
rect 48170 62860 48270 62870
rect 48170 62790 48190 62860
rect 48260 62790 48270 62860
rect 48170 62750 48270 62790
rect 48170 62680 48190 62750
rect 48260 62680 48270 62750
rect 48170 62660 48270 62680
rect 47420 62640 47500 62650
rect 47420 62580 47430 62640
rect 47490 62630 47500 62640
rect 47760 62640 47840 62650
rect 47760 62630 47770 62640
rect 47490 62600 47770 62630
rect 47490 62580 47500 62600
rect 47420 62570 47500 62580
rect 47760 62580 47770 62600
rect 47830 62580 47840 62640
rect 48600 62640 48680 62650
rect 48600 62580 48610 62640
rect 48670 62630 48680 62640
rect 49100 62640 49180 62650
rect 49100 62630 49110 62640
rect 48670 62600 49110 62630
rect 48670 62580 48680 62600
rect 47760 62570 47840 62580
rect 48180 62570 48260 62580
rect 48600 62570 48680 62580
rect 49100 62580 49110 62600
rect 49170 62580 49180 62640
rect 49100 62570 49180 62580
rect 48180 62510 48190 62570
rect 48250 62530 48260 62570
rect 48250 62520 48950 62530
rect 48250 62510 48890 62520
rect 48180 62500 48890 62510
rect 48890 62450 48950 62460
rect 48830 61340 48890 61350
rect 48180 61310 48830 61320
rect 47440 61250 47500 61260
rect 48180 61250 48190 61310
rect 48250 61290 48830 61310
rect 48250 61250 48260 61290
rect 48830 61270 48890 61280
rect 49100 61250 49160 61260
rect 47760 61240 47840 61250
rect 48180 61240 48260 61250
rect 48600 61240 48680 61250
rect 47760 61230 47770 61240
rect 47500 61200 47770 61230
rect 47440 61180 47500 61190
rect 47760 61180 47770 61200
rect 47830 61180 47840 61240
rect 47760 61170 47840 61180
rect 48600 61180 48610 61240
rect 48670 61230 48680 61240
rect 48670 61200 49100 61230
rect 48670 61180 48680 61200
rect 49100 61180 49160 61190
rect 48600 61170 48680 61180
rect 48170 61150 48270 61160
rect 48170 61080 48190 61150
rect 48260 61080 48270 61150
rect 48170 61040 48270 61080
rect 48170 60970 48190 61040
rect 48260 60970 48270 61040
rect 48170 60950 48270 60970
rect 47420 60930 47500 60940
rect 47420 60870 47430 60930
rect 47490 60920 47500 60930
rect 47760 60930 47840 60940
rect 47760 60920 47770 60930
rect 47490 60890 47770 60920
rect 47490 60870 47500 60890
rect 47420 60860 47500 60870
rect 47760 60870 47770 60890
rect 47830 60870 47840 60930
rect 48600 60930 48680 60940
rect 48600 60870 48610 60930
rect 48670 60920 48680 60930
rect 49100 60930 49180 60940
rect 49100 60920 49110 60930
rect 48670 60890 49110 60920
rect 48670 60870 48680 60890
rect 47760 60860 47840 60870
rect 48180 60860 48260 60870
rect 48600 60860 48680 60870
rect 49100 60870 49110 60890
rect 49170 60870 49180 60930
rect 49100 60860 49180 60870
rect 48180 60800 48190 60860
rect 48250 60820 48260 60860
rect 48250 60810 48950 60820
rect 48250 60800 48890 60810
rect 48180 60790 48890 60800
rect 48890 60740 48950 60750
rect 47300 59740 47380 59750
rect 47300 59680 47310 59740
rect 47370 59680 47380 59740
rect 47300 59670 47380 59680
rect 49220 59750 49250 67050
rect 49220 59740 49300 59750
rect 49220 59680 49230 59740
rect 49290 59680 49300 59740
rect 49220 59670 49300 59680
rect 48830 59630 48890 59640
rect 48180 59600 48830 59610
rect 47320 59540 47380 59550
rect 48180 59540 48190 59600
rect 48250 59580 48830 59600
rect 48250 59540 48260 59580
rect 48830 59560 48890 59570
rect 49220 59540 49280 59550
rect 47760 59530 47840 59540
rect 48180 59530 48260 59540
rect 48600 59530 48680 59540
rect 47760 59520 47770 59530
rect 47380 59490 47770 59520
rect 47320 59470 47380 59480
rect 47760 59470 47770 59490
rect 47830 59470 47840 59530
rect 47760 59460 47840 59470
rect 48600 59470 48610 59530
rect 48670 59520 48680 59530
rect 48670 59490 49220 59520
rect 48670 59470 48680 59490
rect 49220 59470 49280 59480
rect 48600 59460 48680 59470
rect 48170 59440 48270 59450
rect 48170 59370 48190 59440
rect 48260 59370 48270 59440
rect 48170 59330 48270 59370
rect 48170 59260 48190 59330
rect 48260 59260 48270 59330
rect 48170 59240 48270 59260
rect 47300 59220 47380 59230
rect 47300 59160 47310 59220
rect 47370 59210 47380 59220
rect 47760 59220 47840 59230
rect 47760 59210 47770 59220
rect 47370 59180 47770 59210
rect 47370 59160 47380 59180
rect 47300 59150 47380 59160
rect 47760 59160 47770 59180
rect 47830 59160 47840 59220
rect 48600 59220 48680 59230
rect 48600 59160 48610 59220
rect 48670 59210 48680 59220
rect 49220 59220 49300 59230
rect 49220 59210 49230 59220
rect 48670 59180 49230 59210
rect 48670 59160 48680 59180
rect 47760 59150 47840 59160
rect 48180 59150 48260 59160
rect 48600 59150 48680 59160
rect 49220 59160 49230 59180
rect 49290 59160 49300 59220
rect 49220 59150 49300 59160
rect 48180 59090 48190 59150
rect 48250 59110 48260 59150
rect 48250 59100 48950 59110
rect 48250 59090 48890 59100
rect 48180 59080 48890 59090
rect 48890 59030 48950 59040
rect 47180 58030 47260 58040
rect 47180 57970 47190 58030
rect 47250 57970 47260 58030
rect 47180 57960 47260 57970
rect 49340 58040 49370 67050
rect 49340 58030 49420 58040
rect 49340 57970 49350 58030
rect 49410 57970 49420 58030
rect 49340 57960 49420 57970
rect 48830 57920 48890 57930
rect 48180 57890 48830 57900
rect 47200 57830 47260 57840
rect 48180 57830 48190 57890
rect 48250 57870 48830 57890
rect 48250 57830 48260 57870
rect 48830 57850 48890 57860
rect 49340 57830 49400 57840
rect 47760 57820 47840 57830
rect 48180 57820 48260 57830
rect 48600 57820 48680 57830
rect 47760 57810 47770 57820
rect 47260 57780 47770 57810
rect 47200 57760 47260 57770
rect 47760 57760 47770 57780
rect 47830 57760 47840 57820
rect 47760 57750 47840 57760
rect 48600 57760 48610 57820
rect 48670 57810 48680 57820
rect 48670 57780 49340 57810
rect 48670 57760 48680 57780
rect 49340 57760 49400 57770
rect 48600 57750 48680 57760
rect 48170 57730 48270 57740
rect 48170 57660 48190 57730
rect 48260 57660 48270 57730
rect 48170 57620 48270 57660
rect 48170 57550 48190 57620
rect 48260 57550 48270 57620
rect 48170 57530 48270 57550
rect 47180 57510 47260 57520
rect 47180 57450 47190 57510
rect 47250 57500 47260 57510
rect 47760 57510 47840 57520
rect 47760 57500 47770 57510
rect 47250 57470 47770 57500
rect 47250 57450 47260 57470
rect 47180 57440 47260 57450
rect 47760 57450 47770 57470
rect 47830 57450 47840 57510
rect 48600 57510 48680 57520
rect 48600 57450 48610 57510
rect 48670 57500 48680 57510
rect 49340 57510 49420 57520
rect 49340 57500 49350 57510
rect 48670 57470 49350 57500
rect 48670 57450 48680 57470
rect 47760 57440 47840 57450
rect 48180 57440 48260 57450
rect 48600 57440 48680 57450
rect 49340 57450 49350 57470
rect 49410 57450 49420 57510
rect 49340 57440 49420 57450
rect 48180 57380 48190 57440
rect 48250 57400 48260 57440
rect 48250 57390 48950 57400
rect 48250 57380 48890 57390
rect 48180 57370 48890 57380
rect 48890 57320 48950 57330
rect 47060 56320 47140 56330
rect 47060 56260 47070 56320
rect 47130 56260 47140 56320
rect 47060 56250 47140 56260
rect 49460 56330 49490 67050
rect 49460 56320 49540 56330
rect 49460 56260 49470 56320
rect 49530 56260 49540 56320
rect 49460 56250 49540 56260
rect 48830 56210 48890 56220
rect 48180 56180 48830 56190
rect 47080 56120 47140 56130
rect 48180 56120 48190 56180
rect 48250 56160 48830 56180
rect 48250 56120 48260 56160
rect 48830 56140 48890 56150
rect 49460 56120 49520 56130
rect 47760 56110 47840 56120
rect 48180 56110 48260 56120
rect 48600 56110 48680 56120
rect 47760 56100 47770 56110
rect 47140 56070 47770 56100
rect 47080 56050 47140 56060
rect 47760 56050 47770 56070
rect 47830 56050 47840 56110
rect 47760 56040 47840 56050
rect 48600 56050 48610 56110
rect 48670 56100 48680 56110
rect 48670 56070 49460 56100
rect 48670 56050 48680 56070
rect 49460 56050 49520 56060
rect 48600 56040 48680 56050
rect 48170 56020 48270 56030
rect 48170 55950 48190 56020
rect 48260 55950 48270 56020
rect 48170 55910 48270 55950
rect 48170 55840 48190 55910
rect 48260 55840 48270 55910
rect 48170 55820 48270 55840
rect 47060 55800 47140 55810
rect 47060 55740 47070 55800
rect 47130 55790 47140 55800
rect 47760 55800 47840 55810
rect 47760 55790 47770 55800
rect 47130 55760 47770 55790
rect 47130 55740 47140 55760
rect 47060 55730 47140 55740
rect 47760 55740 47770 55760
rect 47830 55740 47840 55800
rect 48600 55800 48680 55810
rect 48600 55740 48610 55800
rect 48670 55790 48680 55800
rect 49460 55800 49540 55810
rect 49460 55790 49470 55800
rect 48670 55760 49470 55790
rect 48670 55740 48680 55760
rect 47760 55730 47840 55740
rect 48180 55730 48260 55740
rect 48600 55730 48680 55740
rect 49460 55740 49470 55760
rect 49530 55740 49540 55800
rect 49460 55730 49540 55740
rect 48180 55670 48190 55730
rect 48250 55690 48260 55730
rect 48250 55680 48950 55690
rect 48250 55670 48890 55680
rect 48180 55660 48890 55670
rect 48890 55610 48950 55620
rect 46940 54610 47020 54620
rect 46940 54550 46950 54610
rect 47010 54550 47020 54610
rect 46940 54540 47020 54550
rect 49580 54620 49610 67050
rect 52220 58040 52250 67050
rect 52340 59750 52370 67050
rect 52460 63170 52490 67050
rect 52580 66590 52610 67050
rect 52530 66580 52610 66590
rect 52530 66520 52540 66580
rect 52600 66520 52610 66580
rect 52530 66510 52610 66520
rect 53970 66590 54000 67050
rect 53970 66580 54050 66590
rect 53970 66520 53980 66580
rect 54040 66520 54050 66580
rect 53970 66510 54050 66520
rect 53820 66470 53880 66480
rect 53170 66440 53820 66450
rect 52550 66380 52610 66390
rect 53170 66380 53180 66440
rect 53240 66420 53820 66440
rect 53240 66380 53250 66420
rect 53820 66400 53880 66410
rect 53970 66380 54030 66390
rect 52750 66370 52830 66380
rect 53170 66370 53250 66380
rect 53590 66370 53670 66380
rect 52750 66360 52760 66370
rect 52610 66330 52760 66360
rect 52550 66310 52610 66320
rect 52750 66310 52760 66330
rect 52820 66310 52830 66370
rect 52750 66300 52830 66310
rect 53590 66310 53600 66370
rect 53660 66360 53670 66370
rect 53660 66330 53970 66360
rect 53660 66310 53670 66330
rect 53970 66310 54030 66320
rect 53590 66300 53670 66310
rect 53160 66280 53260 66290
rect 53160 66210 53180 66280
rect 53250 66210 53260 66280
rect 53160 66170 53260 66210
rect 53160 66100 53180 66170
rect 53250 66100 53260 66170
rect 53160 66080 53260 66100
rect 52530 66060 52610 66070
rect 52530 66000 52540 66060
rect 52600 66050 52610 66060
rect 52750 66060 52830 66070
rect 52750 66050 52760 66060
rect 52600 66020 52760 66050
rect 52600 66000 52610 66020
rect 52530 65990 52610 66000
rect 52750 66000 52760 66020
rect 52820 66000 52830 66060
rect 53590 66060 53670 66070
rect 53590 66000 53600 66060
rect 53660 66050 53670 66060
rect 53970 66060 54050 66070
rect 53970 66050 53980 66060
rect 53660 66020 53980 66050
rect 53660 66000 53670 66020
rect 52750 65990 52830 66000
rect 53170 65990 53250 66000
rect 53590 65990 53670 66000
rect 53970 66000 53980 66020
rect 54040 66000 54050 66060
rect 53970 65990 54050 66000
rect 53170 65930 53180 65990
rect 53240 65950 53250 65990
rect 53240 65940 53940 65950
rect 53240 65930 53880 65940
rect 53170 65920 53880 65930
rect 53880 65870 53940 65880
rect 53820 64760 53880 64770
rect 53170 64730 53820 64740
rect 52550 64670 52610 64680
rect 53170 64670 53180 64730
rect 53240 64710 53820 64730
rect 53240 64670 53250 64710
rect 53820 64690 53880 64700
rect 53970 64670 54030 64680
rect 52750 64660 52830 64670
rect 53170 64660 53250 64670
rect 53590 64660 53670 64670
rect 52750 64650 52760 64660
rect 52610 64620 52760 64650
rect 52550 64600 52610 64610
rect 52750 64600 52760 64620
rect 52820 64600 52830 64660
rect 52750 64590 52830 64600
rect 53590 64600 53600 64660
rect 53660 64650 53670 64660
rect 53660 64620 53970 64650
rect 53660 64600 53670 64620
rect 53970 64600 54030 64610
rect 53590 64590 53670 64600
rect 53160 64570 53260 64580
rect 53160 64500 53180 64570
rect 53250 64500 53260 64570
rect 53160 64460 53260 64500
rect 53160 64390 53180 64460
rect 53250 64390 53260 64460
rect 53160 64370 53260 64390
rect 52530 64350 52610 64360
rect 52530 64290 52540 64350
rect 52600 64340 52610 64350
rect 52750 64350 52830 64360
rect 52750 64340 52760 64350
rect 52600 64310 52760 64340
rect 52600 64290 52610 64310
rect 52530 64280 52610 64290
rect 52750 64290 52760 64310
rect 52820 64290 52830 64350
rect 53590 64350 53670 64360
rect 53590 64290 53600 64350
rect 53660 64340 53670 64350
rect 53970 64350 54050 64360
rect 53970 64340 53980 64350
rect 53660 64310 53980 64340
rect 53660 64290 53670 64310
rect 52750 64280 52830 64290
rect 53170 64280 53250 64290
rect 53590 64280 53670 64290
rect 53970 64290 53980 64310
rect 54040 64290 54050 64350
rect 53970 64280 54050 64290
rect 53170 64220 53180 64280
rect 53240 64240 53250 64280
rect 53240 64230 53940 64240
rect 53240 64220 53880 64230
rect 53170 64210 53880 64220
rect 53880 64160 53940 64170
rect 52410 63160 52490 63170
rect 52410 63100 52420 63160
rect 52480 63100 52490 63160
rect 52410 63090 52490 63100
rect 54090 63170 54120 67050
rect 54090 63160 54170 63170
rect 54090 63100 54100 63160
rect 54160 63100 54170 63160
rect 54090 63090 54170 63100
rect 53820 63050 53880 63060
rect 53170 63020 53820 63030
rect 52430 62960 52490 62970
rect 53170 62960 53180 63020
rect 53240 63000 53820 63020
rect 53240 62960 53250 63000
rect 53820 62980 53880 62990
rect 54090 62960 54150 62970
rect 52750 62950 52830 62960
rect 53170 62950 53250 62960
rect 53590 62950 53670 62960
rect 52750 62940 52760 62950
rect 52490 62910 52760 62940
rect 52430 62890 52490 62900
rect 52750 62890 52760 62910
rect 52820 62890 52830 62950
rect 52750 62880 52830 62890
rect 53590 62890 53600 62950
rect 53660 62940 53670 62950
rect 53660 62910 54090 62940
rect 53660 62890 53670 62910
rect 54090 62890 54150 62900
rect 53590 62880 53670 62890
rect 53160 62860 53260 62870
rect 53160 62790 53180 62860
rect 53250 62790 53260 62860
rect 53160 62750 53260 62790
rect 53160 62680 53180 62750
rect 53250 62680 53260 62750
rect 53160 62660 53260 62680
rect 52410 62640 52490 62650
rect 52410 62580 52420 62640
rect 52480 62630 52490 62640
rect 52750 62640 52830 62650
rect 52750 62630 52760 62640
rect 52480 62600 52760 62630
rect 52480 62580 52490 62600
rect 52410 62570 52490 62580
rect 52750 62580 52760 62600
rect 52820 62580 52830 62640
rect 53590 62640 53670 62650
rect 53590 62580 53600 62640
rect 53660 62630 53670 62640
rect 54090 62640 54170 62650
rect 54090 62630 54100 62640
rect 53660 62600 54100 62630
rect 53660 62580 53670 62600
rect 52750 62570 52830 62580
rect 53170 62570 53250 62580
rect 53590 62570 53670 62580
rect 54090 62580 54100 62600
rect 54160 62580 54170 62640
rect 54090 62570 54170 62580
rect 53170 62510 53180 62570
rect 53240 62530 53250 62570
rect 53240 62520 53940 62530
rect 53240 62510 53880 62520
rect 53170 62500 53880 62510
rect 53880 62450 53940 62460
rect 53820 61340 53880 61350
rect 53170 61310 53820 61320
rect 53170 61250 53180 61310
rect 53240 61290 53820 61310
rect 53240 61250 53250 61290
rect 53820 61270 53880 61280
rect 52430 61240 52490 61250
rect 52750 61240 52830 61250
rect 53170 61240 53250 61250
rect 53590 61240 53670 61250
rect 52750 61230 52760 61240
rect 52490 61200 52760 61230
rect 52430 61170 52490 61180
rect 52750 61180 52760 61200
rect 52820 61180 52830 61240
rect 52750 61170 52830 61180
rect 53590 61180 53600 61240
rect 53660 61230 53670 61240
rect 54090 61240 54150 61250
rect 53660 61200 54090 61230
rect 53660 61180 53670 61200
rect 53590 61170 53670 61180
rect 54090 61170 54150 61180
rect 53160 61150 53260 61160
rect 53160 61080 53180 61150
rect 53250 61080 53260 61150
rect 53160 61040 53260 61080
rect 53160 60970 53180 61040
rect 53250 60970 53260 61040
rect 53160 60950 53260 60970
rect 52750 60930 52830 60940
rect 52410 60920 52490 60930
rect 52750 60920 52760 60930
rect 52410 60860 52420 60920
rect 52480 60890 52760 60920
rect 52480 60860 52490 60890
rect 52750 60870 52760 60890
rect 52820 60870 52830 60930
rect 53590 60930 53670 60940
rect 53590 60870 53600 60930
rect 53660 60920 53670 60930
rect 54090 60920 54170 60930
rect 53660 60890 54100 60920
rect 53660 60870 53670 60890
rect 52750 60860 52830 60870
rect 53170 60860 53250 60870
rect 53590 60860 53670 60870
rect 54090 60860 54100 60890
rect 54160 60860 54170 60920
rect 52410 60850 52490 60860
rect 53170 60800 53180 60860
rect 53240 60820 53250 60860
rect 54090 60850 54170 60860
rect 53240 60810 53940 60820
rect 53240 60800 53880 60810
rect 53170 60790 53880 60800
rect 53880 60740 53940 60750
rect 52290 59740 52370 59750
rect 52290 59680 52300 59740
rect 52360 59680 52370 59740
rect 52290 59670 52370 59680
rect 54210 59750 54240 67050
rect 54210 59740 54290 59750
rect 54210 59680 54220 59740
rect 54280 59680 54290 59740
rect 54210 59670 54290 59680
rect 53820 59630 53880 59640
rect 53170 59600 53820 59610
rect 52310 59540 52370 59550
rect 53170 59540 53180 59600
rect 53240 59580 53820 59600
rect 53240 59540 53250 59580
rect 53820 59560 53880 59570
rect 54210 59540 54270 59550
rect 52750 59530 52830 59540
rect 53170 59530 53250 59540
rect 53590 59530 53670 59540
rect 52750 59520 52760 59530
rect 52370 59490 52760 59520
rect 52310 59470 52370 59480
rect 52750 59470 52760 59490
rect 52820 59470 52830 59530
rect 52750 59460 52830 59470
rect 53590 59470 53600 59530
rect 53660 59520 53670 59530
rect 53660 59490 54210 59520
rect 53660 59470 53670 59490
rect 54210 59470 54270 59480
rect 53590 59460 53670 59470
rect 53160 59440 53260 59450
rect 53160 59370 53180 59440
rect 53250 59370 53260 59440
rect 53160 59330 53260 59370
rect 53160 59260 53180 59330
rect 53250 59260 53260 59330
rect 53160 59240 53260 59260
rect 52290 59220 52370 59230
rect 52290 59160 52300 59220
rect 52360 59210 52370 59220
rect 52750 59220 52830 59230
rect 52750 59210 52760 59220
rect 52360 59180 52760 59210
rect 52360 59160 52370 59180
rect 52290 59150 52370 59160
rect 52750 59160 52760 59180
rect 52820 59160 52830 59220
rect 53590 59220 53670 59230
rect 53590 59160 53600 59220
rect 53660 59210 53670 59220
rect 54210 59220 54290 59230
rect 54210 59210 54220 59220
rect 53660 59180 54220 59210
rect 53660 59160 53670 59180
rect 52750 59150 52830 59160
rect 53170 59150 53250 59160
rect 53590 59150 53670 59160
rect 54210 59160 54220 59180
rect 54280 59160 54290 59220
rect 54210 59150 54290 59160
rect 53170 59090 53180 59150
rect 53240 59110 53250 59150
rect 53240 59100 53940 59110
rect 53240 59090 53880 59100
rect 53170 59080 53880 59090
rect 53880 59030 53940 59040
rect 52170 58030 52250 58040
rect 52170 57970 52180 58030
rect 52240 57970 52250 58030
rect 52170 57960 52250 57970
rect 54330 58040 54360 67050
rect 57210 58040 57240 67050
rect 57330 59750 57360 67050
rect 57450 63170 57480 67050
rect 57570 66590 57600 67050
rect 57520 66580 57600 66590
rect 57520 66520 57530 66580
rect 57590 66520 57600 66580
rect 57520 66510 57600 66520
rect 58960 66590 58990 67050
rect 58960 66580 59040 66590
rect 58960 66520 58970 66580
rect 59030 66520 59040 66580
rect 58960 66510 59040 66520
rect 58810 66470 58870 66480
rect 58160 66440 58810 66450
rect 57540 66380 57600 66390
rect 58160 66380 58170 66440
rect 58230 66420 58810 66440
rect 58230 66380 58240 66420
rect 58810 66400 58870 66410
rect 58960 66380 59020 66390
rect 57740 66370 57820 66380
rect 58160 66370 58240 66380
rect 58580 66370 58660 66380
rect 57740 66360 57750 66370
rect 57600 66330 57750 66360
rect 57540 66310 57600 66320
rect 57740 66310 57750 66330
rect 57810 66310 57820 66370
rect 57740 66300 57820 66310
rect 58580 66310 58590 66370
rect 58650 66360 58660 66370
rect 58650 66330 58960 66360
rect 58650 66310 58660 66330
rect 58960 66310 59020 66320
rect 58580 66300 58660 66310
rect 58150 66280 58250 66290
rect 58150 66210 58170 66280
rect 58240 66210 58250 66280
rect 58150 66170 58250 66210
rect 58150 66100 58170 66170
rect 58240 66100 58250 66170
rect 58150 66080 58250 66100
rect 57520 66060 57600 66070
rect 57520 66000 57530 66060
rect 57590 66050 57600 66060
rect 57740 66060 57820 66070
rect 57740 66050 57750 66060
rect 57590 66020 57750 66050
rect 57590 66000 57600 66020
rect 57520 65990 57600 66000
rect 57740 66000 57750 66020
rect 57810 66000 57820 66060
rect 58580 66060 58660 66070
rect 58580 66000 58590 66060
rect 58650 66050 58660 66060
rect 58960 66060 59040 66070
rect 58960 66050 58970 66060
rect 58650 66020 58970 66050
rect 58650 66000 58660 66020
rect 57740 65990 57820 66000
rect 58160 65990 58240 66000
rect 58580 65990 58660 66000
rect 58960 66000 58970 66020
rect 59030 66000 59040 66060
rect 58960 65990 59040 66000
rect 58160 65930 58170 65990
rect 58230 65950 58240 65990
rect 58230 65940 58930 65950
rect 58230 65930 58870 65940
rect 58160 65920 58870 65930
rect 58870 65870 58930 65880
rect 58810 64760 58870 64770
rect 58160 64730 58810 64740
rect 57540 64670 57600 64680
rect 58160 64670 58170 64730
rect 58230 64710 58810 64730
rect 58230 64670 58240 64710
rect 58810 64690 58870 64700
rect 58960 64670 59020 64680
rect 57740 64660 57820 64670
rect 58160 64660 58240 64670
rect 58580 64660 58660 64670
rect 57740 64650 57750 64660
rect 57600 64620 57750 64650
rect 57540 64600 57600 64610
rect 57740 64600 57750 64620
rect 57810 64600 57820 64660
rect 57740 64590 57820 64600
rect 58580 64600 58590 64660
rect 58650 64650 58660 64660
rect 58650 64620 58960 64650
rect 58650 64600 58660 64620
rect 58960 64600 59020 64610
rect 58580 64590 58660 64600
rect 58150 64570 58250 64580
rect 58150 64500 58170 64570
rect 58240 64500 58250 64570
rect 58150 64460 58250 64500
rect 58150 64390 58170 64460
rect 58240 64390 58250 64460
rect 58150 64370 58250 64390
rect 57520 64350 57600 64360
rect 57520 64290 57530 64350
rect 57590 64340 57600 64350
rect 57740 64350 57820 64360
rect 57740 64340 57750 64350
rect 57590 64310 57750 64340
rect 57590 64290 57600 64310
rect 57520 64280 57600 64290
rect 57740 64290 57750 64310
rect 57810 64290 57820 64350
rect 58580 64350 58660 64360
rect 58580 64290 58590 64350
rect 58650 64340 58660 64350
rect 58960 64350 59040 64360
rect 58960 64340 58970 64350
rect 58650 64310 58970 64340
rect 58650 64290 58660 64310
rect 57740 64280 57820 64290
rect 58160 64280 58240 64290
rect 58580 64280 58660 64290
rect 58960 64290 58970 64310
rect 59030 64290 59040 64350
rect 58960 64280 59040 64290
rect 58160 64220 58170 64280
rect 58230 64240 58240 64280
rect 58230 64230 58930 64240
rect 58230 64220 58870 64230
rect 58160 64210 58870 64220
rect 58870 64160 58930 64170
rect 57400 63160 57480 63170
rect 57400 63100 57410 63160
rect 57470 63100 57480 63160
rect 57400 63090 57480 63100
rect 59080 63170 59110 67050
rect 59080 63160 59160 63170
rect 59080 63100 59090 63160
rect 59150 63100 59160 63160
rect 59080 63090 59160 63100
rect 58810 63050 58870 63060
rect 58160 63020 58810 63030
rect 57420 62960 57480 62970
rect 58160 62960 58170 63020
rect 58230 63000 58810 63020
rect 58230 62960 58240 63000
rect 58810 62980 58870 62990
rect 59080 62960 59140 62970
rect 57740 62950 57820 62960
rect 58160 62950 58240 62960
rect 58580 62950 58660 62960
rect 57740 62940 57750 62950
rect 57480 62910 57750 62940
rect 57420 62890 57480 62900
rect 57740 62890 57750 62910
rect 57810 62890 57820 62950
rect 57740 62880 57820 62890
rect 58580 62890 58590 62950
rect 58650 62940 58660 62950
rect 58650 62910 59080 62940
rect 58650 62890 58660 62910
rect 59080 62890 59140 62900
rect 58580 62880 58660 62890
rect 58150 62860 58250 62870
rect 58150 62790 58170 62860
rect 58240 62790 58250 62860
rect 58150 62750 58250 62790
rect 58150 62680 58170 62750
rect 58240 62680 58250 62750
rect 58150 62660 58250 62680
rect 57400 62640 57480 62650
rect 57400 62580 57410 62640
rect 57470 62630 57480 62640
rect 57740 62640 57820 62650
rect 57740 62630 57750 62640
rect 57470 62600 57750 62630
rect 57470 62580 57480 62600
rect 57400 62570 57480 62580
rect 57740 62580 57750 62600
rect 57810 62580 57820 62640
rect 58580 62640 58660 62650
rect 58580 62580 58590 62640
rect 58650 62630 58660 62640
rect 59080 62640 59160 62650
rect 59080 62630 59090 62640
rect 58650 62600 59090 62630
rect 58650 62580 58660 62600
rect 57740 62570 57820 62580
rect 58160 62570 58240 62580
rect 58580 62570 58660 62580
rect 59080 62580 59090 62600
rect 59150 62580 59160 62640
rect 59080 62570 59160 62580
rect 58160 62510 58170 62570
rect 58230 62530 58240 62570
rect 58230 62520 58930 62530
rect 58230 62510 58870 62520
rect 58160 62500 58870 62510
rect 58870 62450 58930 62460
rect 58810 61340 58870 61350
rect 58160 61310 58810 61320
rect 58160 61250 58170 61310
rect 58230 61290 58810 61310
rect 58230 61250 58240 61290
rect 58810 61270 58870 61280
rect 57420 61240 57480 61250
rect 57740 61240 57820 61250
rect 58160 61240 58240 61250
rect 58580 61240 58660 61250
rect 57740 61230 57750 61240
rect 57480 61200 57750 61230
rect 57420 61170 57480 61180
rect 57740 61180 57750 61200
rect 57810 61180 57820 61240
rect 57740 61170 57820 61180
rect 58580 61180 58590 61240
rect 58650 61230 58660 61240
rect 59080 61240 59140 61250
rect 58650 61200 59080 61230
rect 58650 61180 58660 61200
rect 58580 61170 58660 61180
rect 59080 61170 59140 61180
rect 58150 61150 58250 61160
rect 58150 61080 58170 61150
rect 58240 61080 58250 61150
rect 58150 61040 58250 61080
rect 58150 60970 58170 61040
rect 58240 60970 58250 61040
rect 58150 60950 58250 60970
rect 57740 60930 57820 60940
rect 57400 60920 57480 60930
rect 57740 60920 57750 60930
rect 57400 60860 57410 60920
rect 57470 60890 57750 60920
rect 57470 60860 57480 60890
rect 57740 60870 57750 60890
rect 57810 60870 57820 60930
rect 58580 60930 58660 60940
rect 58580 60870 58590 60930
rect 58650 60920 58660 60930
rect 59080 60920 59160 60930
rect 58650 60890 59090 60920
rect 58650 60870 58660 60890
rect 57740 60860 57820 60870
rect 58160 60860 58240 60870
rect 58580 60860 58660 60870
rect 59080 60860 59090 60890
rect 59150 60860 59160 60920
rect 57400 60850 57480 60860
rect 58160 60800 58170 60860
rect 58230 60820 58240 60860
rect 59080 60850 59160 60860
rect 58230 60810 58930 60820
rect 58230 60800 58870 60810
rect 58160 60790 58870 60800
rect 58870 60740 58930 60750
rect 57280 59740 57360 59750
rect 57280 59680 57290 59740
rect 57350 59680 57360 59740
rect 57280 59670 57360 59680
rect 59200 59750 59230 67050
rect 59200 59740 59280 59750
rect 59200 59680 59210 59740
rect 59270 59680 59280 59740
rect 59200 59670 59280 59680
rect 58810 59630 58870 59640
rect 58160 59600 58810 59610
rect 57300 59540 57360 59550
rect 58160 59540 58170 59600
rect 58230 59580 58810 59600
rect 58230 59540 58240 59580
rect 58810 59560 58870 59570
rect 59200 59540 59260 59550
rect 57740 59530 57820 59540
rect 58160 59530 58240 59540
rect 58580 59530 58660 59540
rect 57740 59520 57750 59530
rect 57360 59490 57750 59520
rect 57300 59470 57360 59480
rect 57740 59470 57750 59490
rect 57810 59470 57820 59530
rect 57740 59460 57820 59470
rect 58580 59470 58590 59530
rect 58650 59520 58660 59530
rect 58650 59490 59200 59520
rect 58650 59470 58660 59490
rect 59200 59470 59260 59480
rect 58580 59460 58660 59470
rect 58150 59440 58250 59450
rect 58150 59370 58170 59440
rect 58240 59370 58250 59440
rect 58150 59330 58250 59370
rect 58150 59260 58170 59330
rect 58240 59260 58250 59330
rect 58150 59240 58250 59260
rect 57280 59220 57360 59230
rect 57280 59160 57290 59220
rect 57350 59210 57360 59220
rect 57740 59220 57820 59230
rect 57740 59210 57750 59220
rect 57350 59180 57750 59210
rect 57350 59160 57360 59180
rect 57280 59150 57360 59160
rect 57740 59160 57750 59180
rect 57810 59160 57820 59220
rect 58580 59220 58660 59230
rect 58580 59160 58590 59220
rect 58650 59210 58660 59220
rect 59200 59220 59280 59230
rect 59200 59210 59210 59220
rect 58650 59180 59210 59210
rect 58650 59160 58660 59180
rect 57740 59150 57820 59160
rect 58160 59150 58240 59160
rect 58580 59150 58660 59160
rect 59200 59160 59210 59180
rect 59270 59160 59280 59220
rect 59200 59150 59280 59160
rect 58160 59090 58170 59150
rect 58230 59110 58240 59150
rect 58230 59100 58930 59110
rect 58230 59090 58870 59100
rect 58160 59080 58870 59090
rect 58870 59030 58930 59040
rect 54330 58030 54410 58040
rect 54330 57970 54340 58030
rect 54400 57970 54410 58030
rect 54330 57960 54410 57970
rect 57160 58030 57240 58040
rect 57160 57970 57170 58030
rect 57230 57970 57240 58030
rect 57160 57960 57240 57970
rect 59320 58040 59350 67050
rect 62440 59750 62470 67050
rect 62560 66590 62590 67050
rect 62510 66580 62590 66590
rect 62510 66520 62520 66580
rect 62580 66520 62590 66580
rect 62510 66510 62590 66520
rect 63950 66590 63980 67050
rect 63950 66580 64030 66590
rect 63950 66520 63960 66580
rect 64020 66520 64030 66580
rect 63950 66510 64030 66520
rect 63800 66470 63860 66480
rect 63150 66440 63800 66450
rect 62530 66380 62590 66390
rect 63150 66380 63160 66440
rect 63220 66420 63800 66440
rect 63220 66380 63230 66420
rect 63800 66400 63860 66410
rect 63950 66380 64010 66390
rect 62730 66370 62810 66380
rect 63150 66370 63230 66380
rect 63570 66370 63650 66380
rect 62730 66360 62740 66370
rect 62590 66330 62740 66360
rect 62530 66310 62590 66320
rect 62730 66310 62740 66330
rect 62800 66310 62810 66370
rect 62730 66300 62810 66310
rect 63570 66310 63580 66370
rect 63640 66360 63650 66370
rect 63640 66330 63950 66360
rect 63640 66310 63650 66330
rect 63950 66310 64010 66320
rect 63570 66300 63650 66310
rect 63140 66280 63240 66290
rect 63140 66210 63160 66280
rect 63230 66210 63240 66280
rect 63140 66170 63240 66210
rect 63140 66100 63160 66170
rect 63230 66100 63240 66170
rect 63140 66080 63240 66100
rect 62510 66060 62590 66070
rect 62510 66000 62520 66060
rect 62580 66050 62590 66060
rect 62730 66060 62810 66070
rect 62730 66050 62740 66060
rect 62580 66020 62740 66050
rect 62580 66000 62590 66020
rect 62510 65990 62590 66000
rect 62730 66000 62740 66020
rect 62800 66000 62810 66060
rect 63570 66060 63650 66070
rect 63570 66000 63580 66060
rect 63640 66050 63650 66060
rect 63950 66060 64030 66070
rect 63950 66050 63960 66060
rect 63640 66020 63960 66050
rect 63640 66000 63650 66020
rect 62730 65990 62810 66000
rect 63150 65990 63230 66000
rect 63570 65990 63650 66000
rect 63950 66000 63960 66020
rect 64020 66000 64030 66060
rect 63950 65990 64030 66000
rect 63150 65930 63160 65990
rect 63220 65950 63230 65990
rect 63220 65940 63920 65950
rect 63220 65930 63860 65940
rect 63150 65920 63860 65930
rect 63860 65870 63920 65880
rect 63800 64760 63860 64770
rect 63150 64730 63800 64740
rect 62530 64670 62590 64680
rect 63150 64670 63160 64730
rect 63220 64710 63800 64730
rect 63220 64670 63230 64710
rect 63800 64690 63860 64700
rect 63950 64670 64010 64680
rect 62730 64660 62810 64670
rect 63150 64660 63230 64670
rect 63570 64660 63650 64670
rect 62730 64650 62740 64660
rect 62590 64620 62740 64650
rect 62530 64600 62590 64610
rect 62730 64600 62740 64620
rect 62800 64600 62810 64660
rect 62730 64590 62810 64600
rect 63570 64600 63580 64660
rect 63640 64650 63650 64660
rect 63640 64620 63950 64650
rect 63640 64600 63650 64620
rect 63950 64600 64010 64610
rect 63570 64590 63650 64600
rect 63140 64570 63240 64580
rect 63140 64500 63160 64570
rect 63230 64500 63240 64570
rect 63140 64460 63240 64500
rect 63140 64390 63160 64460
rect 63230 64390 63240 64460
rect 63140 64370 63240 64390
rect 62510 64350 62590 64360
rect 62510 64290 62520 64350
rect 62580 64340 62590 64350
rect 62730 64350 62810 64360
rect 62730 64340 62740 64350
rect 62580 64310 62740 64340
rect 62580 64290 62590 64310
rect 62510 64280 62590 64290
rect 62730 64290 62740 64310
rect 62800 64290 62810 64350
rect 63570 64350 63650 64360
rect 63570 64290 63580 64350
rect 63640 64340 63650 64350
rect 63950 64350 64030 64360
rect 63950 64340 63960 64350
rect 63640 64310 63960 64340
rect 63640 64290 63650 64310
rect 62730 64280 62810 64290
rect 63150 64280 63230 64290
rect 63570 64280 63650 64290
rect 63950 64290 63960 64310
rect 64020 64290 64030 64350
rect 63950 64280 64030 64290
rect 63150 64220 63160 64280
rect 63220 64240 63230 64280
rect 63220 64230 63920 64240
rect 63220 64220 63860 64230
rect 63150 64210 63860 64220
rect 63860 64160 63920 64170
rect 63800 63050 63860 63060
rect 63150 63020 63800 63030
rect 62530 62960 62590 62970
rect 63150 62960 63160 63020
rect 63220 63000 63800 63020
rect 63220 62960 63230 63000
rect 63800 62980 63860 62990
rect 63950 62960 64010 62970
rect 62730 62950 62810 62960
rect 63150 62950 63230 62960
rect 63570 62950 63650 62960
rect 62730 62940 62740 62950
rect 62590 62910 62740 62940
rect 62530 62890 62590 62900
rect 62730 62890 62740 62910
rect 62800 62890 62810 62950
rect 62730 62880 62810 62890
rect 63570 62890 63580 62950
rect 63640 62940 63650 62950
rect 63640 62910 63950 62940
rect 63640 62890 63650 62910
rect 63950 62890 64010 62900
rect 63570 62880 63650 62890
rect 63140 62860 63240 62870
rect 63140 62790 63160 62860
rect 63230 62790 63240 62860
rect 63140 62750 63240 62790
rect 63140 62680 63160 62750
rect 63230 62680 63240 62750
rect 63140 62660 63240 62680
rect 62510 62640 62590 62650
rect 62510 62580 62520 62640
rect 62580 62630 62590 62640
rect 62730 62640 62810 62650
rect 62730 62630 62740 62640
rect 62580 62600 62740 62630
rect 62580 62580 62590 62600
rect 62510 62570 62590 62580
rect 62730 62580 62740 62600
rect 62800 62580 62810 62640
rect 63570 62640 63650 62650
rect 63570 62580 63580 62640
rect 63640 62630 63650 62640
rect 63950 62640 64030 62650
rect 63950 62630 63960 62640
rect 63640 62600 63960 62630
rect 63640 62580 63650 62600
rect 62730 62570 62810 62580
rect 63150 62570 63230 62580
rect 63570 62570 63650 62580
rect 63950 62580 63960 62600
rect 64020 62580 64030 62640
rect 63950 62570 64030 62580
rect 63150 62510 63160 62570
rect 63220 62530 63230 62570
rect 63220 62520 63920 62530
rect 63220 62510 63860 62520
rect 63150 62500 63860 62510
rect 63860 62450 63920 62460
rect 63800 61340 63860 61350
rect 63150 61310 63800 61320
rect 62530 61250 62590 61260
rect 63150 61250 63160 61310
rect 63220 61290 63800 61310
rect 63220 61250 63230 61290
rect 63800 61270 63860 61280
rect 63950 61250 64010 61260
rect 62730 61240 62810 61250
rect 63150 61240 63230 61250
rect 63570 61240 63650 61250
rect 62730 61230 62740 61240
rect 62590 61200 62740 61230
rect 62530 61180 62590 61190
rect 62730 61180 62740 61200
rect 62800 61180 62810 61240
rect 62730 61170 62810 61180
rect 63570 61180 63580 61240
rect 63640 61230 63650 61240
rect 63640 61200 63950 61230
rect 63640 61180 63650 61200
rect 63950 61180 64010 61190
rect 63570 61170 63650 61180
rect 63140 61150 63240 61160
rect 63140 61080 63160 61150
rect 63230 61080 63240 61150
rect 63140 61040 63240 61080
rect 63140 60970 63160 61040
rect 63230 60970 63240 61040
rect 63140 60950 63240 60970
rect 62510 60930 62590 60940
rect 62510 60870 62520 60930
rect 62580 60920 62590 60930
rect 62730 60930 62810 60940
rect 62730 60920 62740 60930
rect 62580 60890 62740 60920
rect 62580 60870 62590 60890
rect 62510 60860 62590 60870
rect 62730 60870 62740 60890
rect 62800 60870 62810 60930
rect 63570 60930 63650 60940
rect 63570 60870 63580 60930
rect 63640 60920 63650 60930
rect 63950 60930 64030 60940
rect 63950 60920 63960 60930
rect 63640 60890 63960 60920
rect 63640 60870 63650 60890
rect 62730 60860 62810 60870
rect 63150 60860 63230 60870
rect 63570 60860 63650 60870
rect 63950 60870 63960 60890
rect 64020 60870 64030 60930
rect 63950 60860 64030 60870
rect 63150 60800 63160 60860
rect 63220 60820 63230 60860
rect 63220 60810 63920 60820
rect 63220 60800 63860 60810
rect 63150 60790 63860 60800
rect 63860 60740 63920 60750
rect 62390 59740 62470 59750
rect 62390 59680 62400 59740
rect 62460 59680 62470 59740
rect 62390 59670 62470 59680
rect 64070 59750 64100 67050
rect 67430 59750 67460 67050
rect 67550 66590 67580 67050
rect 67500 66580 67580 66590
rect 67500 66520 67510 66580
rect 67570 66520 67580 66580
rect 67500 66510 67580 66520
rect 68940 66590 68970 67050
rect 68940 66580 69020 66590
rect 68940 66520 68950 66580
rect 69010 66520 69020 66580
rect 68940 66510 69020 66520
rect 68790 66470 68850 66480
rect 68140 66440 68790 66450
rect 67520 66380 67580 66390
rect 68140 66380 68150 66440
rect 68210 66420 68790 66440
rect 68210 66380 68220 66420
rect 68790 66400 68850 66410
rect 68940 66380 69000 66390
rect 67720 66370 67800 66380
rect 68140 66370 68220 66380
rect 68560 66370 68640 66380
rect 67720 66360 67730 66370
rect 67580 66330 67730 66360
rect 67520 66310 67580 66320
rect 67720 66310 67730 66330
rect 67790 66310 67800 66370
rect 67720 66300 67800 66310
rect 68560 66310 68570 66370
rect 68630 66360 68640 66370
rect 68630 66330 68940 66360
rect 68630 66310 68640 66330
rect 68940 66310 69000 66320
rect 68560 66300 68640 66310
rect 68130 66280 68230 66290
rect 68130 66210 68150 66280
rect 68220 66210 68230 66280
rect 68130 66170 68230 66210
rect 68130 66100 68150 66170
rect 68220 66100 68230 66170
rect 68130 66080 68230 66100
rect 67500 66060 67580 66070
rect 67500 66000 67510 66060
rect 67570 66050 67580 66060
rect 67720 66060 67800 66070
rect 67720 66050 67730 66060
rect 67570 66020 67730 66050
rect 67570 66000 67580 66020
rect 67500 65990 67580 66000
rect 67720 66000 67730 66020
rect 67790 66000 67800 66060
rect 68560 66060 68640 66070
rect 68560 66000 68570 66060
rect 68630 66050 68640 66060
rect 68940 66060 69020 66070
rect 68940 66050 68950 66060
rect 68630 66020 68950 66050
rect 68630 66000 68640 66020
rect 67720 65990 67800 66000
rect 68140 65990 68220 66000
rect 68560 65990 68640 66000
rect 68940 66000 68950 66020
rect 69010 66000 69020 66060
rect 68940 65990 69020 66000
rect 68140 65930 68150 65990
rect 68210 65950 68220 65990
rect 68210 65940 68910 65950
rect 68210 65930 68850 65940
rect 68140 65920 68850 65930
rect 68850 65870 68910 65880
rect 68790 64760 68850 64770
rect 68140 64730 68790 64740
rect 67520 64670 67580 64680
rect 68140 64670 68150 64730
rect 68210 64710 68790 64730
rect 68210 64670 68220 64710
rect 68790 64690 68850 64700
rect 68940 64670 69000 64680
rect 67720 64660 67800 64670
rect 68140 64660 68220 64670
rect 68560 64660 68640 64670
rect 67720 64650 67730 64660
rect 67580 64620 67730 64650
rect 67520 64600 67580 64610
rect 67720 64600 67730 64620
rect 67790 64600 67800 64660
rect 67720 64590 67800 64600
rect 68560 64600 68570 64660
rect 68630 64650 68640 64660
rect 68630 64620 68940 64650
rect 68630 64600 68640 64620
rect 68940 64600 69000 64610
rect 68560 64590 68640 64600
rect 68130 64570 68230 64580
rect 68130 64500 68150 64570
rect 68220 64500 68230 64570
rect 68130 64460 68230 64500
rect 68130 64390 68150 64460
rect 68220 64390 68230 64460
rect 68130 64370 68230 64390
rect 67500 64350 67580 64360
rect 67500 64290 67510 64350
rect 67570 64340 67580 64350
rect 67720 64350 67800 64360
rect 67720 64340 67730 64350
rect 67570 64310 67730 64340
rect 67570 64290 67580 64310
rect 67500 64280 67580 64290
rect 67720 64290 67730 64310
rect 67790 64290 67800 64350
rect 68560 64350 68640 64360
rect 68560 64290 68570 64350
rect 68630 64340 68640 64350
rect 68940 64350 69020 64360
rect 68940 64340 68950 64350
rect 68630 64310 68950 64340
rect 68630 64290 68640 64310
rect 67720 64280 67800 64290
rect 68140 64280 68220 64290
rect 68560 64280 68640 64290
rect 68940 64290 68950 64310
rect 69010 64290 69020 64350
rect 68940 64280 69020 64290
rect 68140 64220 68150 64280
rect 68210 64240 68220 64280
rect 68210 64230 68910 64240
rect 68210 64220 68850 64230
rect 68140 64210 68850 64220
rect 68850 64160 68910 64170
rect 68790 63050 68850 63060
rect 68140 63020 68790 63030
rect 67520 62960 67580 62970
rect 68140 62960 68150 63020
rect 68210 63000 68790 63020
rect 68210 62960 68220 63000
rect 68790 62980 68850 62990
rect 68940 62960 69000 62970
rect 67720 62950 67800 62960
rect 68140 62950 68220 62960
rect 68560 62950 68640 62960
rect 67720 62940 67730 62950
rect 67580 62910 67730 62940
rect 67520 62890 67580 62900
rect 67720 62890 67730 62910
rect 67790 62890 67800 62950
rect 67720 62880 67800 62890
rect 68560 62890 68570 62950
rect 68630 62940 68640 62950
rect 68630 62910 68940 62940
rect 68630 62890 68640 62910
rect 68940 62890 69000 62900
rect 68560 62880 68640 62890
rect 68130 62860 68230 62870
rect 68130 62790 68150 62860
rect 68220 62790 68230 62860
rect 68130 62750 68230 62790
rect 68130 62680 68150 62750
rect 68220 62680 68230 62750
rect 68130 62660 68230 62680
rect 67500 62640 67580 62650
rect 67500 62580 67510 62640
rect 67570 62630 67580 62640
rect 67720 62640 67800 62650
rect 67720 62630 67730 62640
rect 67570 62600 67730 62630
rect 67570 62580 67580 62600
rect 67500 62570 67580 62580
rect 67720 62580 67730 62600
rect 67790 62580 67800 62640
rect 68560 62640 68640 62650
rect 68560 62580 68570 62640
rect 68630 62630 68640 62640
rect 68940 62640 69020 62650
rect 68940 62630 68950 62640
rect 68630 62600 68950 62630
rect 68630 62580 68640 62600
rect 67720 62570 67800 62580
rect 68140 62570 68220 62580
rect 68560 62570 68640 62580
rect 68940 62580 68950 62600
rect 69010 62580 69020 62640
rect 68940 62570 69020 62580
rect 68140 62510 68150 62570
rect 68210 62530 68220 62570
rect 68210 62520 68910 62530
rect 68210 62510 68850 62520
rect 68140 62500 68850 62510
rect 68850 62450 68910 62460
rect 68790 61340 68850 61350
rect 68140 61310 68790 61320
rect 67520 61250 67580 61260
rect 68140 61250 68150 61310
rect 68210 61290 68790 61310
rect 68210 61250 68220 61290
rect 68790 61270 68850 61280
rect 68940 61250 69000 61260
rect 67720 61240 67800 61250
rect 68140 61240 68220 61250
rect 68560 61240 68640 61250
rect 67720 61230 67730 61240
rect 67580 61200 67730 61230
rect 67520 61180 67580 61190
rect 67720 61180 67730 61200
rect 67790 61180 67800 61240
rect 67720 61170 67800 61180
rect 68560 61180 68570 61240
rect 68630 61230 68640 61240
rect 68630 61200 68940 61230
rect 68630 61180 68640 61200
rect 68940 61180 69000 61190
rect 68560 61170 68640 61180
rect 68130 61150 68230 61160
rect 68130 61080 68150 61150
rect 68220 61080 68230 61150
rect 68130 61040 68230 61080
rect 68130 60970 68150 61040
rect 68220 60970 68230 61040
rect 68130 60950 68230 60970
rect 67500 60930 67580 60940
rect 67500 60870 67510 60930
rect 67570 60920 67580 60930
rect 67720 60930 67800 60940
rect 67720 60920 67730 60930
rect 67570 60890 67730 60920
rect 67570 60870 67580 60890
rect 67500 60860 67580 60870
rect 67720 60870 67730 60890
rect 67790 60870 67800 60930
rect 68560 60930 68640 60940
rect 68560 60870 68570 60930
rect 68630 60920 68640 60930
rect 68940 60930 69020 60940
rect 68940 60920 68950 60930
rect 68630 60890 68950 60920
rect 68630 60870 68640 60890
rect 67720 60860 67800 60870
rect 68140 60860 68220 60870
rect 68560 60860 68640 60870
rect 68940 60870 68950 60890
rect 69010 60870 69020 60930
rect 68940 60860 69020 60870
rect 68140 60800 68150 60860
rect 68210 60820 68220 60860
rect 68210 60810 68910 60820
rect 68210 60800 68850 60810
rect 68140 60790 68850 60800
rect 68850 60740 68910 60750
rect 64070 59740 64150 59750
rect 64070 59680 64080 59740
rect 64140 59680 64150 59740
rect 64070 59670 64150 59680
rect 67380 59740 67460 59750
rect 67380 59680 67390 59740
rect 67450 59680 67460 59740
rect 67380 59670 67460 59680
rect 69060 59750 69090 67050
rect 72540 66590 72570 67050
rect 72490 66580 72570 66590
rect 72490 66520 72500 66580
rect 72560 66520 72570 66580
rect 72490 66510 72570 66520
rect 73930 66590 73960 67050
rect 77530 66590 77560 67050
rect 73930 66580 74010 66590
rect 73930 66520 73940 66580
rect 74000 66520 74010 66580
rect 73930 66510 74010 66520
rect 77480 66580 77560 66590
rect 77480 66520 77490 66580
rect 77550 66520 77560 66580
rect 77480 66510 77560 66520
rect 78920 66590 78950 67050
rect 78920 66580 79000 66590
rect 78920 66520 78930 66580
rect 78990 66520 79000 66580
rect 78920 66510 79000 66520
rect 73780 66470 73840 66480
rect 73130 66440 73780 66450
rect 72510 66380 72570 66390
rect 73130 66380 73140 66440
rect 73200 66420 73780 66440
rect 73200 66380 73210 66420
rect 78770 66470 78830 66480
rect 73780 66400 73840 66410
rect 78120 66440 78770 66450
rect 73930 66380 73990 66390
rect 72710 66370 72790 66380
rect 73130 66370 73210 66380
rect 73550 66370 73630 66380
rect 72710 66360 72720 66370
rect 72570 66330 72720 66360
rect 72510 66310 72570 66320
rect 72710 66310 72720 66330
rect 72780 66310 72790 66370
rect 72710 66300 72790 66310
rect 73550 66310 73560 66370
rect 73620 66360 73630 66370
rect 73620 66330 73930 66360
rect 73620 66310 73630 66330
rect 73930 66310 73990 66320
rect 77500 66380 77560 66390
rect 78120 66380 78130 66440
rect 78190 66420 78770 66440
rect 78190 66380 78200 66420
rect 78770 66400 78830 66410
rect 78920 66380 78980 66390
rect 77700 66370 77780 66380
rect 78120 66370 78200 66380
rect 78540 66370 78620 66380
rect 77700 66360 77710 66370
rect 77560 66330 77710 66360
rect 77500 66310 77560 66320
rect 77700 66310 77710 66330
rect 77770 66310 77780 66370
rect 73550 66300 73630 66310
rect 77700 66300 77780 66310
rect 78540 66310 78550 66370
rect 78610 66360 78620 66370
rect 78610 66330 78920 66360
rect 78610 66310 78620 66330
rect 78920 66310 78980 66320
rect 78540 66300 78620 66310
rect 73120 66280 73220 66290
rect 73120 66210 73140 66280
rect 73210 66210 73220 66280
rect 73120 66170 73220 66210
rect 73120 66100 73140 66170
rect 73210 66100 73220 66170
rect 73120 66080 73220 66100
rect 78110 66280 78210 66290
rect 78110 66210 78130 66280
rect 78200 66210 78210 66280
rect 78110 66170 78210 66210
rect 78110 66100 78130 66170
rect 78200 66100 78210 66170
rect 78110 66080 78210 66100
rect 72490 66060 72570 66070
rect 72490 66000 72500 66060
rect 72560 66050 72570 66060
rect 72710 66060 72790 66070
rect 72710 66050 72720 66060
rect 72560 66020 72720 66050
rect 72560 66000 72570 66020
rect 72490 65990 72570 66000
rect 72710 66000 72720 66020
rect 72780 66000 72790 66060
rect 73550 66060 73630 66070
rect 73550 66000 73560 66060
rect 73620 66050 73630 66060
rect 73930 66060 74010 66070
rect 73930 66050 73940 66060
rect 73620 66020 73940 66050
rect 73620 66000 73630 66020
rect 72710 65990 72790 66000
rect 73130 65990 73210 66000
rect 73550 65990 73630 66000
rect 73930 66000 73940 66020
rect 74000 66000 74010 66060
rect 73930 65990 74010 66000
rect 77480 66060 77560 66070
rect 77480 66000 77490 66060
rect 77550 66050 77560 66060
rect 77700 66060 77780 66070
rect 77700 66050 77710 66060
rect 77550 66020 77710 66050
rect 77550 66000 77560 66020
rect 77480 65990 77560 66000
rect 77700 66000 77710 66020
rect 77770 66000 77780 66060
rect 78540 66060 78620 66070
rect 78540 66000 78550 66060
rect 78610 66050 78620 66060
rect 78920 66060 79000 66070
rect 78920 66050 78930 66060
rect 78610 66020 78930 66050
rect 78610 66000 78620 66020
rect 77700 65990 77780 66000
rect 78120 65990 78200 66000
rect 78540 65990 78620 66000
rect 78920 66000 78930 66020
rect 78990 66000 79000 66060
rect 78920 65990 79000 66000
rect 73130 65930 73140 65990
rect 73200 65950 73210 65990
rect 73200 65940 73900 65950
rect 73200 65930 73840 65940
rect 73130 65920 73840 65930
rect 78120 65930 78130 65990
rect 78190 65950 78200 65990
rect 78190 65940 78890 65950
rect 78190 65930 78830 65940
rect 78120 65920 78830 65930
rect 73840 65870 73900 65880
rect 78830 65870 78890 65880
rect 73780 64760 73840 64770
rect 73130 64730 73780 64740
rect 72510 64670 72570 64680
rect 73130 64670 73140 64730
rect 73200 64710 73780 64730
rect 73200 64670 73210 64710
rect 78770 64760 78830 64770
rect 73780 64690 73840 64700
rect 78120 64730 78770 64740
rect 73930 64670 73990 64680
rect 72710 64660 72790 64670
rect 73130 64660 73210 64670
rect 73550 64660 73630 64670
rect 72710 64650 72720 64660
rect 72570 64620 72720 64650
rect 72510 64600 72570 64610
rect 72710 64600 72720 64620
rect 72780 64600 72790 64660
rect 72710 64590 72790 64600
rect 73550 64600 73560 64660
rect 73620 64650 73630 64660
rect 73620 64620 73930 64650
rect 73620 64600 73630 64620
rect 73930 64600 73990 64610
rect 77500 64670 77560 64680
rect 78120 64670 78130 64730
rect 78190 64710 78770 64730
rect 78190 64670 78200 64710
rect 78770 64690 78830 64700
rect 78920 64670 78980 64680
rect 77700 64660 77780 64670
rect 78120 64660 78200 64670
rect 78540 64660 78620 64670
rect 77700 64650 77710 64660
rect 77560 64620 77710 64650
rect 77500 64600 77560 64610
rect 77700 64600 77710 64620
rect 77770 64600 77780 64660
rect 73550 64590 73630 64600
rect 77700 64590 77780 64600
rect 78540 64600 78550 64660
rect 78610 64650 78620 64660
rect 78610 64620 78920 64650
rect 78610 64600 78620 64620
rect 78920 64600 78980 64610
rect 78540 64590 78620 64600
rect 73120 64570 73220 64580
rect 73120 64500 73140 64570
rect 73210 64500 73220 64570
rect 73120 64460 73220 64500
rect 73120 64390 73140 64460
rect 73210 64390 73220 64460
rect 73120 64370 73220 64390
rect 78110 64570 78210 64580
rect 78110 64500 78130 64570
rect 78200 64500 78210 64570
rect 78110 64460 78210 64500
rect 78110 64390 78130 64460
rect 78200 64390 78210 64460
rect 78110 64370 78210 64390
rect 72490 64350 72570 64360
rect 72490 64290 72500 64350
rect 72560 64340 72570 64350
rect 72710 64350 72790 64360
rect 72710 64340 72720 64350
rect 72560 64310 72720 64340
rect 72560 64290 72570 64310
rect 72490 64280 72570 64290
rect 72710 64290 72720 64310
rect 72780 64290 72790 64350
rect 73550 64350 73630 64360
rect 73550 64290 73560 64350
rect 73620 64340 73630 64350
rect 73930 64350 74010 64360
rect 73930 64340 73940 64350
rect 73620 64310 73940 64340
rect 73620 64290 73630 64310
rect 72710 64280 72790 64290
rect 73130 64280 73210 64290
rect 73550 64280 73630 64290
rect 73930 64290 73940 64310
rect 74000 64290 74010 64350
rect 73930 64280 74010 64290
rect 77480 64350 77560 64360
rect 77480 64290 77490 64350
rect 77550 64340 77560 64350
rect 77700 64350 77780 64360
rect 77700 64340 77710 64350
rect 77550 64310 77710 64340
rect 77550 64290 77560 64310
rect 77480 64280 77560 64290
rect 77700 64290 77710 64310
rect 77770 64290 77780 64350
rect 78540 64350 78620 64360
rect 78540 64290 78550 64350
rect 78610 64340 78620 64350
rect 78920 64350 79000 64360
rect 78920 64340 78930 64350
rect 78610 64310 78930 64340
rect 78610 64290 78620 64310
rect 77700 64280 77780 64290
rect 78120 64280 78200 64290
rect 78540 64280 78620 64290
rect 78920 64290 78930 64310
rect 78990 64290 79000 64350
rect 78920 64280 79000 64290
rect 73130 64220 73140 64280
rect 73200 64240 73210 64280
rect 73200 64230 73900 64240
rect 73200 64220 73840 64230
rect 73130 64210 73840 64220
rect 78120 64220 78130 64280
rect 78190 64240 78200 64280
rect 78190 64230 78890 64240
rect 78190 64220 78830 64230
rect 78120 64210 78830 64220
rect 73840 64160 73900 64170
rect 78830 64160 78890 64170
rect 73780 63050 73840 63060
rect 73130 63020 73780 63030
rect 72510 62960 72570 62970
rect 73130 62960 73140 63020
rect 73200 63000 73780 63020
rect 73200 62960 73210 63000
rect 78770 63050 78830 63060
rect 73780 62980 73840 62990
rect 78120 63020 78770 63030
rect 73930 62960 73990 62970
rect 72710 62950 72790 62960
rect 73130 62950 73210 62960
rect 73550 62950 73630 62960
rect 72710 62940 72720 62950
rect 72570 62910 72720 62940
rect 72510 62890 72570 62900
rect 72710 62890 72720 62910
rect 72780 62890 72790 62950
rect 72710 62880 72790 62890
rect 73550 62890 73560 62950
rect 73620 62940 73630 62950
rect 73620 62910 73930 62940
rect 73620 62890 73630 62910
rect 73930 62890 73990 62900
rect 77500 62960 77560 62970
rect 78120 62960 78130 63020
rect 78190 63000 78770 63020
rect 78190 62960 78200 63000
rect 78770 62980 78830 62990
rect 78920 62960 78980 62970
rect 77700 62950 77780 62960
rect 78120 62950 78200 62960
rect 78540 62950 78620 62960
rect 77700 62940 77710 62950
rect 77560 62910 77710 62940
rect 77500 62890 77560 62900
rect 77700 62890 77710 62910
rect 77770 62890 77780 62950
rect 73550 62880 73630 62890
rect 77700 62880 77780 62890
rect 78540 62890 78550 62950
rect 78610 62940 78620 62950
rect 78610 62910 78920 62940
rect 78610 62890 78620 62910
rect 78920 62890 78980 62900
rect 78540 62880 78620 62890
rect 73120 62860 73220 62870
rect 73120 62790 73140 62860
rect 73210 62790 73220 62860
rect 73120 62750 73220 62790
rect 73120 62680 73140 62750
rect 73210 62680 73220 62750
rect 73120 62660 73220 62680
rect 78110 62860 78210 62870
rect 78110 62790 78130 62860
rect 78200 62790 78210 62860
rect 78110 62750 78210 62790
rect 78110 62680 78130 62750
rect 78200 62680 78210 62750
rect 78110 62660 78210 62680
rect 72490 62640 72570 62650
rect 72490 62580 72500 62640
rect 72560 62630 72570 62640
rect 72710 62640 72790 62650
rect 72710 62630 72720 62640
rect 72560 62600 72720 62630
rect 72560 62580 72570 62600
rect 72490 62570 72570 62580
rect 72710 62580 72720 62600
rect 72780 62580 72790 62640
rect 73550 62640 73630 62650
rect 73550 62580 73560 62640
rect 73620 62630 73630 62640
rect 73930 62640 74010 62650
rect 73930 62630 73940 62640
rect 73620 62600 73940 62630
rect 73620 62580 73630 62600
rect 72710 62570 72790 62580
rect 73130 62570 73210 62580
rect 73550 62570 73630 62580
rect 73930 62580 73940 62600
rect 74000 62580 74010 62640
rect 73930 62570 74010 62580
rect 77480 62640 77560 62650
rect 77480 62580 77490 62640
rect 77550 62630 77560 62640
rect 77700 62640 77780 62650
rect 77700 62630 77710 62640
rect 77550 62600 77710 62630
rect 77550 62580 77560 62600
rect 77480 62570 77560 62580
rect 77700 62580 77710 62600
rect 77770 62580 77780 62640
rect 78540 62640 78620 62650
rect 78540 62580 78550 62640
rect 78610 62630 78620 62640
rect 78920 62640 79000 62650
rect 78920 62630 78930 62640
rect 78610 62600 78930 62630
rect 78610 62580 78620 62600
rect 77700 62570 77780 62580
rect 78120 62570 78200 62580
rect 78540 62570 78620 62580
rect 78920 62580 78930 62600
rect 78990 62580 79000 62640
rect 78920 62570 79000 62580
rect 73130 62510 73140 62570
rect 73200 62530 73210 62570
rect 73200 62520 73900 62530
rect 73200 62510 73840 62520
rect 73130 62500 73840 62510
rect 78120 62510 78130 62570
rect 78190 62530 78200 62570
rect 78190 62520 78890 62530
rect 78190 62510 78830 62520
rect 78120 62500 78830 62510
rect 73840 62450 73900 62460
rect 78830 62450 78890 62460
rect 73780 61340 73840 61350
rect 73130 61310 73780 61320
rect 72510 61250 72570 61260
rect 73130 61250 73140 61310
rect 73200 61290 73780 61310
rect 73200 61250 73210 61290
rect 78770 61340 78830 61350
rect 73780 61270 73840 61280
rect 78120 61310 78770 61320
rect 73930 61250 73990 61260
rect 72710 61240 72790 61250
rect 73130 61240 73210 61250
rect 73550 61240 73630 61250
rect 72710 61230 72720 61240
rect 72570 61200 72720 61230
rect 72510 61180 72570 61190
rect 72710 61180 72720 61200
rect 72780 61180 72790 61240
rect 72710 61170 72790 61180
rect 73550 61180 73560 61240
rect 73620 61230 73630 61240
rect 73620 61200 73930 61230
rect 73620 61180 73630 61200
rect 73930 61180 73990 61190
rect 77500 61250 77560 61260
rect 78120 61250 78130 61310
rect 78190 61290 78770 61310
rect 78190 61250 78200 61290
rect 78770 61270 78830 61280
rect 78920 61250 78980 61260
rect 77700 61240 77780 61250
rect 78120 61240 78200 61250
rect 78540 61240 78620 61250
rect 77700 61230 77710 61240
rect 77560 61200 77710 61230
rect 77500 61180 77560 61190
rect 77700 61180 77710 61200
rect 77770 61180 77780 61240
rect 73550 61170 73630 61180
rect 77700 61170 77780 61180
rect 78540 61180 78550 61240
rect 78610 61230 78620 61240
rect 78610 61200 78920 61230
rect 78610 61180 78620 61200
rect 78920 61180 78980 61190
rect 78540 61170 78620 61180
rect 73120 61150 73220 61160
rect 73120 61080 73140 61150
rect 73210 61080 73220 61150
rect 73120 61040 73220 61080
rect 73120 60970 73140 61040
rect 73210 60970 73220 61040
rect 73120 60950 73220 60970
rect 78110 61150 78210 61160
rect 78110 61080 78130 61150
rect 78200 61080 78210 61150
rect 78110 61040 78210 61080
rect 78110 60970 78130 61040
rect 78200 60970 78210 61040
rect 78110 60950 78210 60970
rect 72490 60930 72570 60940
rect 72490 60870 72500 60930
rect 72560 60920 72570 60930
rect 72710 60930 72790 60940
rect 72710 60920 72720 60930
rect 72560 60890 72720 60920
rect 72560 60870 72570 60890
rect 72490 60860 72570 60870
rect 72710 60870 72720 60890
rect 72780 60870 72790 60930
rect 73550 60930 73630 60940
rect 73550 60870 73560 60930
rect 73620 60920 73630 60930
rect 73930 60930 74010 60940
rect 73930 60920 73940 60930
rect 73620 60890 73940 60920
rect 73620 60870 73630 60890
rect 72710 60860 72790 60870
rect 73130 60860 73210 60870
rect 73550 60860 73630 60870
rect 73930 60870 73940 60890
rect 74000 60870 74010 60930
rect 73930 60860 74010 60870
rect 77480 60930 77560 60940
rect 77480 60870 77490 60930
rect 77550 60920 77560 60930
rect 77700 60930 77780 60940
rect 77700 60920 77710 60930
rect 77550 60890 77710 60920
rect 77550 60870 77560 60890
rect 77480 60860 77560 60870
rect 77700 60870 77710 60890
rect 77770 60870 77780 60930
rect 78540 60930 78620 60940
rect 78540 60870 78550 60930
rect 78610 60920 78620 60930
rect 78920 60930 79000 60940
rect 78920 60920 78930 60930
rect 78610 60890 78930 60920
rect 78610 60870 78620 60890
rect 77700 60860 77780 60870
rect 78120 60860 78200 60870
rect 78540 60860 78620 60870
rect 78920 60870 78930 60890
rect 78990 60870 79000 60930
rect 78920 60860 79000 60870
rect 73130 60800 73140 60860
rect 73200 60820 73210 60860
rect 73200 60810 73900 60820
rect 73200 60800 73840 60810
rect 73130 60790 73840 60800
rect 78120 60800 78130 60860
rect 78190 60820 78200 60860
rect 78190 60810 78890 60820
rect 78190 60800 78830 60810
rect 78120 60790 78830 60800
rect 73840 60740 73900 60750
rect 78830 60740 78890 60750
rect 69060 59740 69140 59750
rect 69060 59680 69070 59740
rect 69130 59680 69140 59740
rect 69060 59670 69140 59680
rect 63800 59630 63860 59640
rect 63150 59600 63800 59610
rect 62410 59540 62470 59550
rect 63150 59540 63160 59600
rect 63220 59580 63800 59600
rect 63220 59540 63230 59580
rect 68790 59630 68850 59640
rect 63800 59560 63860 59570
rect 68140 59600 68790 59610
rect 64070 59540 64130 59550
rect 62730 59530 62810 59540
rect 63150 59530 63230 59540
rect 63570 59530 63650 59540
rect 62730 59520 62740 59530
rect 62470 59490 62740 59520
rect 62410 59470 62470 59480
rect 62730 59470 62740 59490
rect 62800 59470 62810 59530
rect 62730 59460 62810 59470
rect 63570 59470 63580 59530
rect 63640 59520 63650 59530
rect 63640 59490 64070 59520
rect 63640 59470 63650 59490
rect 64070 59470 64130 59480
rect 67400 59540 67460 59550
rect 68140 59540 68150 59600
rect 68210 59580 68790 59600
rect 68210 59540 68220 59580
rect 73780 59630 73840 59640
rect 68790 59560 68850 59570
rect 73130 59600 73780 59610
rect 69060 59540 69120 59550
rect 67720 59530 67800 59540
rect 68140 59530 68220 59540
rect 68560 59530 68640 59540
rect 67720 59520 67730 59530
rect 67460 59490 67730 59520
rect 67400 59470 67460 59480
rect 67720 59470 67730 59490
rect 67790 59470 67800 59530
rect 63570 59460 63650 59470
rect 67720 59460 67800 59470
rect 68560 59470 68570 59530
rect 68630 59520 68640 59530
rect 68630 59490 69060 59520
rect 68630 59470 68640 59490
rect 69060 59470 69120 59480
rect 72510 59540 72570 59550
rect 73130 59540 73140 59600
rect 73200 59580 73780 59600
rect 73200 59540 73210 59580
rect 78770 59630 78830 59640
rect 73780 59560 73840 59570
rect 78120 59600 78770 59610
rect 73930 59540 73990 59550
rect 72710 59530 72790 59540
rect 73130 59530 73210 59540
rect 73550 59530 73630 59540
rect 72710 59520 72720 59530
rect 72570 59490 72720 59520
rect 72510 59470 72570 59480
rect 72710 59470 72720 59490
rect 72780 59470 72790 59530
rect 68560 59460 68640 59470
rect 72710 59460 72790 59470
rect 73550 59470 73560 59530
rect 73620 59520 73630 59530
rect 73620 59490 73930 59520
rect 73620 59470 73630 59490
rect 73930 59470 73990 59480
rect 77500 59540 77560 59550
rect 78120 59540 78130 59600
rect 78190 59580 78770 59600
rect 78190 59540 78200 59580
rect 78770 59560 78830 59570
rect 78920 59540 78980 59550
rect 77700 59530 77780 59540
rect 78120 59530 78200 59540
rect 78540 59530 78620 59540
rect 77700 59520 77710 59530
rect 77560 59490 77710 59520
rect 77500 59470 77560 59480
rect 77700 59470 77710 59490
rect 77770 59470 77780 59530
rect 73550 59460 73630 59470
rect 77700 59460 77780 59470
rect 78540 59470 78550 59530
rect 78610 59520 78620 59530
rect 78610 59490 78920 59520
rect 78610 59470 78620 59490
rect 78920 59470 78980 59480
rect 78540 59460 78620 59470
rect 63140 59440 63240 59450
rect 63140 59370 63160 59440
rect 63230 59370 63240 59440
rect 63140 59330 63240 59370
rect 63140 59260 63160 59330
rect 63230 59260 63240 59330
rect 63140 59240 63240 59260
rect 68130 59440 68230 59450
rect 68130 59370 68150 59440
rect 68220 59370 68230 59440
rect 68130 59330 68230 59370
rect 68130 59260 68150 59330
rect 68220 59260 68230 59330
rect 68130 59240 68230 59260
rect 73120 59440 73220 59450
rect 73120 59370 73140 59440
rect 73210 59370 73220 59440
rect 73120 59330 73220 59370
rect 73120 59260 73140 59330
rect 73210 59260 73220 59330
rect 73120 59240 73220 59260
rect 78110 59440 78210 59450
rect 78110 59370 78130 59440
rect 78200 59370 78210 59440
rect 78110 59330 78210 59370
rect 78110 59260 78130 59330
rect 78200 59260 78210 59330
rect 78110 59240 78210 59260
rect 62390 59220 62470 59230
rect 62390 59160 62400 59220
rect 62460 59210 62470 59220
rect 62730 59220 62810 59230
rect 62730 59210 62740 59220
rect 62460 59180 62740 59210
rect 62460 59160 62470 59180
rect 62390 59150 62470 59160
rect 62730 59160 62740 59180
rect 62800 59160 62810 59220
rect 63570 59220 63650 59230
rect 63570 59160 63580 59220
rect 63640 59210 63650 59220
rect 64070 59220 64150 59230
rect 64070 59210 64080 59220
rect 63640 59180 64080 59210
rect 63640 59160 63650 59180
rect 62730 59150 62810 59160
rect 63150 59150 63230 59160
rect 63570 59150 63650 59160
rect 64070 59160 64080 59180
rect 64140 59160 64150 59220
rect 64070 59150 64150 59160
rect 67380 59220 67460 59230
rect 67380 59160 67390 59220
rect 67450 59210 67460 59220
rect 67720 59220 67800 59230
rect 67720 59210 67730 59220
rect 67450 59180 67730 59210
rect 67450 59160 67460 59180
rect 67380 59150 67460 59160
rect 67720 59160 67730 59180
rect 67790 59160 67800 59220
rect 68560 59220 68640 59230
rect 68560 59160 68570 59220
rect 68630 59210 68640 59220
rect 69060 59220 69140 59230
rect 69060 59210 69070 59220
rect 68630 59180 69070 59210
rect 68630 59160 68640 59180
rect 67720 59150 67800 59160
rect 68140 59150 68220 59160
rect 68560 59150 68640 59160
rect 69060 59160 69070 59180
rect 69130 59160 69140 59220
rect 69060 59150 69140 59160
rect 72490 59220 72570 59230
rect 72490 59160 72500 59220
rect 72560 59210 72570 59220
rect 72710 59220 72790 59230
rect 72710 59210 72720 59220
rect 72560 59180 72720 59210
rect 72560 59160 72570 59180
rect 72490 59150 72570 59160
rect 72710 59160 72720 59180
rect 72780 59160 72790 59220
rect 73550 59220 73630 59230
rect 73550 59160 73560 59220
rect 73620 59210 73630 59220
rect 73930 59220 74010 59230
rect 73930 59210 73940 59220
rect 73620 59180 73940 59210
rect 73620 59160 73630 59180
rect 72710 59150 72790 59160
rect 73130 59150 73210 59160
rect 73550 59150 73630 59160
rect 73930 59160 73940 59180
rect 74000 59160 74010 59220
rect 73930 59150 74010 59160
rect 77480 59220 77560 59230
rect 77480 59160 77490 59220
rect 77550 59210 77560 59220
rect 77700 59220 77780 59230
rect 77700 59210 77710 59220
rect 77550 59180 77710 59210
rect 77550 59160 77560 59180
rect 77480 59150 77560 59160
rect 77700 59160 77710 59180
rect 77770 59160 77780 59220
rect 78540 59220 78620 59230
rect 78540 59160 78550 59220
rect 78610 59210 78620 59220
rect 78920 59220 79000 59230
rect 78920 59210 78930 59220
rect 78610 59180 78930 59210
rect 78610 59160 78620 59180
rect 77700 59150 77780 59160
rect 78120 59150 78200 59160
rect 78540 59150 78620 59160
rect 78920 59160 78930 59180
rect 78990 59160 79000 59220
rect 78920 59150 79000 59160
rect 63150 59090 63160 59150
rect 63220 59110 63230 59150
rect 63220 59100 63920 59110
rect 63220 59090 63860 59100
rect 63150 59080 63860 59090
rect 68140 59090 68150 59150
rect 68210 59110 68220 59150
rect 68210 59100 68910 59110
rect 68210 59090 68850 59100
rect 68140 59080 68850 59090
rect 63860 59030 63920 59040
rect 73130 59090 73140 59150
rect 73200 59110 73210 59150
rect 73200 59100 73900 59110
rect 73200 59090 73840 59100
rect 73130 59080 73840 59090
rect 68850 59030 68910 59040
rect 78120 59090 78130 59150
rect 78190 59110 78200 59150
rect 78190 59100 78890 59110
rect 78190 59090 78830 59100
rect 78120 59080 78830 59090
rect 73840 59030 73900 59040
rect 78830 59030 78890 59040
rect 59320 58030 59400 58040
rect 59320 57970 59330 58030
rect 59390 57970 59400 58030
rect 59320 57960 59400 57970
rect 53820 57920 53880 57930
rect 53170 57890 53820 57900
rect 52190 57830 52250 57840
rect 53170 57830 53180 57890
rect 53240 57870 53820 57890
rect 53240 57830 53250 57870
rect 58810 57920 58870 57930
rect 53820 57850 53880 57860
rect 58160 57890 58810 57900
rect 54330 57830 54390 57840
rect 52750 57820 52830 57830
rect 53170 57820 53250 57830
rect 53590 57820 53670 57830
rect 52750 57810 52760 57820
rect 52250 57780 52760 57810
rect 52190 57760 52250 57770
rect 52750 57760 52760 57780
rect 52820 57760 52830 57820
rect 52750 57750 52830 57760
rect 53590 57760 53600 57820
rect 53660 57810 53670 57820
rect 53660 57780 54330 57810
rect 53660 57760 53670 57780
rect 54330 57760 54390 57770
rect 57180 57830 57240 57840
rect 58160 57830 58170 57890
rect 58230 57870 58810 57890
rect 58230 57830 58240 57870
rect 63800 57920 63860 57930
rect 58810 57850 58870 57860
rect 63150 57890 63800 57900
rect 59320 57830 59380 57840
rect 57740 57820 57820 57830
rect 58160 57820 58240 57830
rect 58580 57820 58660 57830
rect 57740 57810 57750 57820
rect 57240 57780 57750 57810
rect 57180 57760 57240 57770
rect 57740 57760 57750 57780
rect 57810 57760 57820 57820
rect 53590 57750 53670 57760
rect 57740 57750 57820 57760
rect 58580 57760 58590 57820
rect 58650 57810 58660 57820
rect 58650 57780 59320 57810
rect 58650 57760 58660 57780
rect 59320 57760 59380 57770
rect 62410 57830 62470 57840
rect 63150 57830 63160 57890
rect 63220 57870 63800 57890
rect 63220 57830 63230 57870
rect 68790 57920 68850 57930
rect 63800 57850 63860 57860
rect 68140 57890 68790 57900
rect 64070 57830 64130 57840
rect 62730 57820 62810 57830
rect 63150 57820 63230 57830
rect 63570 57820 63650 57830
rect 62730 57810 62740 57820
rect 62470 57780 62740 57810
rect 62410 57760 62470 57770
rect 62730 57760 62740 57780
rect 62800 57760 62810 57820
rect 58580 57750 58660 57760
rect 62730 57750 62810 57760
rect 63570 57760 63580 57820
rect 63640 57810 63650 57820
rect 63640 57780 64070 57810
rect 63640 57760 63650 57780
rect 64070 57760 64130 57770
rect 67400 57830 67460 57840
rect 68140 57830 68150 57890
rect 68210 57870 68790 57890
rect 68210 57830 68220 57870
rect 73780 57920 73840 57930
rect 68790 57850 68850 57860
rect 73130 57890 73780 57900
rect 69060 57830 69120 57840
rect 67720 57820 67800 57830
rect 68140 57820 68220 57830
rect 68560 57820 68640 57830
rect 67720 57810 67730 57820
rect 67460 57780 67730 57810
rect 67400 57760 67460 57770
rect 67720 57760 67730 57780
rect 67790 57760 67800 57820
rect 63570 57750 63650 57760
rect 67720 57750 67800 57760
rect 68560 57760 68570 57820
rect 68630 57810 68640 57820
rect 68630 57780 69060 57810
rect 68630 57760 68640 57780
rect 69060 57760 69120 57770
rect 72510 57830 72570 57840
rect 73130 57830 73140 57890
rect 73200 57870 73780 57890
rect 73200 57830 73210 57870
rect 78770 57920 78830 57930
rect 73780 57850 73840 57860
rect 78120 57890 78770 57900
rect 73930 57830 73990 57840
rect 72710 57820 72790 57830
rect 73130 57820 73210 57830
rect 73550 57820 73630 57830
rect 72710 57810 72720 57820
rect 72570 57780 72720 57810
rect 72510 57760 72570 57770
rect 72710 57760 72720 57780
rect 72780 57760 72790 57820
rect 68560 57750 68640 57760
rect 72710 57750 72790 57760
rect 73550 57760 73560 57820
rect 73620 57810 73630 57820
rect 73620 57780 73930 57810
rect 73620 57760 73630 57780
rect 73930 57760 73990 57770
rect 77500 57830 77560 57840
rect 78120 57830 78130 57890
rect 78190 57870 78770 57890
rect 78190 57830 78200 57870
rect 78770 57850 78830 57860
rect 78920 57830 78980 57840
rect 77700 57820 77780 57830
rect 78120 57820 78200 57830
rect 78540 57820 78620 57830
rect 77700 57810 77710 57820
rect 77560 57780 77710 57810
rect 77500 57760 77560 57770
rect 77700 57760 77710 57780
rect 77770 57760 77780 57820
rect 73550 57750 73630 57760
rect 77700 57750 77780 57760
rect 78540 57760 78550 57820
rect 78610 57810 78620 57820
rect 78610 57780 78920 57810
rect 78610 57760 78620 57780
rect 78920 57760 78980 57770
rect 78540 57750 78620 57760
rect 53160 57730 53260 57740
rect 53160 57660 53180 57730
rect 53250 57660 53260 57730
rect 53160 57620 53260 57660
rect 53160 57550 53180 57620
rect 53250 57550 53260 57620
rect 53160 57530 53260 57550
rect 58150 57730 58250 57740
rect 58150 57660 58170 57730
rect 58240 57660 58250 57730
rect 58150 57620 58250 57660
rect 58150 57550 58170 57620
rect 58240 57550 58250 57620
rect 58150 57530 58250 57550
rect 63140 57730 63240 57740
rect 63140 57660 63160 57730
rect 63230 57660 63240 57730
rect 63140 57620 63240 57660
rect 63140 57550 63160 57620
rect 63230 57550 63240 57620
rect 63140 57530 63240 57550
rect 68130 57730 68230 57740
rect 68130 57660 68150 57730
rect 68220 57660 68230 57730
rect 68130 57620 68230 57660
rect 68130 57550 68150 57620
rect 68220 57550 68230 57620
rect 68130 57530 68230 57550
rect 73120 57730 73220 57740
rect 73120 57660 73140 57730
rect 73210 57660 73220 57730
rect 73120 57620 73220 57660
rect 73120 57550 73140 57620
rect 73210 57550 73220 57620
rect 73120 57530 73220 57550
rect 78110 57730 78210 57740
rect 78110 57660 78130 57730
rect 78200 57660 78210 57730
rect 78110 57620 78210 57660
rect 78110 57550 78130 57620
rect 78200 57550 78210 57620
rect 78110 57530 78210 57550
rect 52170 57510 52250 57520
rect 52170 57450 52180 57510
rect 52240 57500 52250 57510
rect 52750 57510 52830 57520
rect 52750 57500 52760 57510
rect 52240 57470 52760 57500
rect 52240 57450 52250 57470
rect 52170 57440 52250 57450
rect 52750 57450 52760 57470
rect 52820 57450 52830 57510
rect 53590 57510 53670 57520
rect 53590 57450 53600 57510
rect 53660 57500 53670 57510
rect 54330 57510 54410 57520
rect 54330 57500 54340 57510
rect 53660 57470 54340 57500
rect 53660 57450 53670 57470
rect 52750 57440 52830 57450
rect 53170 57440 53250 57450
rect 53590 57440 53670 57450
rect 54330 57450 54340 57470
rect 54400 57450 54410 57510
rect 54330 57440 54410 57450
rect 57160 57510 57240 57520
rect 57160 57450 57170 57510
rect 57230 57500 57240 57510
rect 57740 57510 57820 57520
rect 57740 57500 57750 57510
rect 57230 57470 57750 57500
rect 57230 57450 57240 57470
rect 57160 57440 57240 57450
rect 57740 57450 57750 57470
rect 57810 57450 57820 57510
rect 58580 57510 58660 57520
rect 58580 57450 58590 57510
rect 58650 57500 58660 57510
rect 59320 57510 59400 57520
rect 59320 57500 59330 57510
rect 58650 57470 59330 57500
rect 58650 57450 58660 57470
rect 57740 57440 57820 57450
rect 58160 57440 58240 57450
rect 58580 57440 58660 57450
rect 59320 57450 59330 57470
rect 59390 57450 59400 57510
rect 59320 57440 59400 57450
rect 62390 57510 62470 57520
rect 62390 57450 62400 57510
rect 62460 57500 62470 57510
rect 62730 57510 62810 57520
rect 62730 57500 62740 57510
rect 62460 57470 62740 57500
rect 62460 57450 62470 57470
rect 62390 57440 62470 57450
rect 62730 57450 62740 57470
rect 62800 57450 62810 57510
rect 63570 57510 63650 57520
rect 63570 57450 63580 57510
rect 63640 57500 63650 57510
rect 64070 57510 64150 57520
rect 64070 57500 64080 57510
rect 63640 57470 64080 57500
rect 63640 57450 63650 57470
rect 62730 57440 62810 57450
rect 63150 57440 63230 57450
rect 63570 57440 63650 57450
rect 64070 57450 64080 57470
rect 64140 57450 64150 57510
rect 64070 57440 64150 57450
rect 67380 57510 67460 57520
rect 67380 57450 67390 57510
rect 67450 57500 67460 57510
rect 67720 57510 67800 57520
rect 67720 57500 67730 57510
rect 67450 57470 67730 57500
rect 67450 57450 67460 57470
rect 67380 57440 67460 57450
rect 67720 57450 67730 57470
rect 67790 57450 67800 57510
rect 68560 57510 68640 57520
rect 68560 57450 68570 57510
rect 68630 57500 68640 57510
rect 69060 57510 69140 57520
rect 69060 57500 69070 57510
rect 68630 57470 69070 57500
rect 68630 57450 68640 57470
rect 67720 57440 67800 57450
rect 68140 57440 68220 57450
rect 68560 57440 68640 57450
rect 69060 57450 69070 57470
rect 69130 57450 69140 57510
rect 69060 57440 69140 57450
rect 72490 57510 72570 57520
rect 72490 57450 72500 57510
rect 72560 57500 72570 57510
rect 72710 57510 72790 57520
rect 72710 57500 72720 57510
rect 72560 57470 72720 57500
rect 72560 57450 72570 57470
rect 72490 57440 72570 57450
rect 72710 57450 72720 57470
rect 72780 57450 72790 57510
rect 73550 57510 73630 57520
rect 73550 57450 73560 57510
rect 73620 57500 73630 57510
rect 73930 57510 74010 57520
rect 73930 57500 73940 57510
rect 73620 57470 73940 57500
rect 73620 57450 73630 57470
rect 72710 57440 72790 57450
rect 73130 57440 73210 57450
rect 73550 57440 73630 57450
rect 73930 57450 73940 57470
rect 74000 57450 74010 57510
rect 73930 57440 74010 57450
rect 77480 57510 77560 57520
rect 77480 57450 77490 57510
rect 77550 57500 77560 57510
rect 77700 57510 77780 57520
rect 77700 57500 77710 57510
rect 77550 57470 77710 57500
rect 77550 57450 77560 57470
rect 77480 57440 77560 57450
rect 77700 57450 77710 57470
rect 77770 57450 77780 57510
rect 78540 57510 78620 57520
rect 78540 57450 78550 57510
rect 78610 57500 78620 57510
rect 78920 57510 79000 57520
rect 78920 57500 78930 57510
rect 78610 57470 78930 57500
rect 78610 57450 78620 57470
rect 77700 57440 77780 57450
rect 78120 57440 78200 57450
rect 78540 57440 78620 57450
rect 78920 57450 78930 57470
rect 78990 57450 79000 57510
rect 78920 57440 79000 57450
rect 53170 57380 53180 57440
rect 53240 57400 53250 57440
rect 53240 57390 53940 57400
rect 53240 57380 53880 57390
rect 53170 57370 53880 57380
rect 58160 57380 58170 57440
rect 58230 57400 58240 57440
rect 58230 57390 58930 57400
rect 58230 57380 58870 57390
rect 58160 57370 58870 57380
rect 53880 57320 53940 57330
rect 63150 57380 63160 57440
rect 63220 57400 63230 57440
rect 63220 57390 63920 57400
rect 63220 57380 63860 57390
rect 63150 57370 63860 57380
rect 58870 57320 58930 57330
rect 68140 57380 68150 57440
rect 68210 57400 68220 57440
rect 68210 57390 68910 57400
rect 68210 57380 68850 57390
rect 68140 57370 68850 57380
rect 63860 57320 63920 57330
rect 73130 57380 73140 57440
rect 73200 57400 73210 57440
rect 73200 57390 73900 57400
rect 73200 57380 73840 57390
rect 73130 57370 73840 57380
rect 68850 57320 68910 57330
rect 78120 57380 78130 57440
rect 78190 57400 78200 57440
rect 78190 57390 78890 57400
rect 78190 57380 78830 57390
rect 78120 57370 78830 57380
rect 73840 57320 73900 57330
rect 78830 57320 78890 57330
rect 53820 56210 53880 56220
rect 53170 56180 53820 56190
rect 52190 56120 52250 56130
rect 53170 56120 53180 56180
rect 53240 56160 53820 56180
rect 53240 56120 53250 56160
rect 58810 56210 58870 56220
rect 53820 56140 53880 56150
rect 58160 56180 58810 56190
rect 54330 56120 54390 56130
rect 52750 56110 52830 56120
rect 53170 56110 53250 56120
rect 53590 56110 53670 56120
rect 52750 56100 52760 56110
rect 52250 56070 52760 56100
rect 52190 56050 52250 56060
rect 52750 56050 52760 56070
rect 52820 56050 52830 56110
rect 52750 56040 52830 56050
rect 53590 56050 53600 56110
rect 53660 56100 53670 56110
rect 53660 56070 54330 56100
rect 53660 56050 53670 56070
rect 54330 56050 54390 56060
rect 57180 56120 57240 56130
rect 58160 56120 58170 56180
rect 58230 56160 58810 56180
rect 58230 56120 58240 56160
rect 63800 56210 63860 56220
rect 58810 56140 58870 56150
rect 63150 56180 63800 56190
rect 59320 56120 59380 56130
rect 57740 56110 57820 56120
rect 58160 56110 58240 56120
rect 58580 56110 58660 56120
rect 57740 56100 57750 56110
rect 57240 56070 57750 56100
rect 57180 56050 57240 56060
rect 57740 56050 57750 56070
rect 57810 56050 57820 56110
rect 53590 56040 53670 56050
rect 57740 56040 57820 56050
rect 58580 56050 58590 56110
rect 58650 56100 58660 56110
rect 58650 56070 59320 56100
rect 58650 56050 58660 56070
rect 59320 56050 59380 56060
rect 62410 56120 62470 56130
rect 63150 56120 63160 56180
rect 63220 56160 63800 56180
rect 63220 56120 63230 56160
rect 68790 56210 68850 56220
rect 63800 56140 63860 56150
rect 68140 56180 68790 56190
rect 64070 56120 64130 56130
rect 62730 56110 62810 56120
rect 63150 56110 63230 56120
rect 63570 56110 63650 56120
rect 62730 56100 62740 56110
rect 62470 56070 62740 56100
rect 62410 56050 62470 56060
rect 62730 56050 62740 56070
rect 62800 56050 62810 56110
rect 58580 56040 58660 56050
rect 62730 56040 62810 56050
rect 63570 56050 63580 56110
rect 63640 56100 63650 56110
rect 63640 56070 64070 56100
rect 63640 56050 63650 56070
rect 64070 56050 64130 56060
rect 67400 56120 67460 56130
rect 68140 56120 68150 56180
rect 68210 56160 68790 56180
rect 68210 56120 68220 56160
rect 73780 56210 73840 56220
rect 68790 56140 68850 56150
rect 73130 56180 73780 56190
rect 69060 56120 69120 56130
rect 67720 56110 67800 56120
rect 68140 56110 68220 56120
rect 68560 56110 68640 56120
rect 67720 56100 67730 56110
rect 67460 56070 67730 56100
rect 67400 56050 67460 56060
rect 67720 56050 67730 56070
rect 67790 56050 67800 56110
rect 63570 56040 63650 56050
rect 67720 56040 67800 56050
rect 68560 56050 68570 56110
rect 68630 56100 68640 56110
rect 68630 56070 69060 56100
rect 68630 56050 68640 56070
rect 69060 56050 69120 56060
rect 72510 56120 72570 56130
rect 73130 56120 73140 56180
rect 73200 56160 73780 56180
rect 73200 56120 73210 56160
rect 78770 56210 78830 56220
rect 73780 56140 73840 56150
rect 78120 56180 78770 56190
rect 73930 56120 73990 56130
rect 72710 56110 72790 56120
rect 73130 56110 73210 56120
rect 73550 56110 73630 56120
rect 72710 56100 72720 56110
rect 72570 56070 72720 56100
rect 72510 56050 72570 56060
rect 72710 56050 72720 56070
rect 72780 56050 72790 56110
rect 68560 56040 68640 56050
rect 72710 56040 72790 56050
rect 73550 56050 73560 56110
rect 73620 56100 73630 56110
rect 73620 56070 73930 56100
rect 73620 56050 73630 56070
rect 73930 56050 73990 56060
rect 77500 56120 77560 56130
rect 78120 56120 78130 56180
rect 78190 56160 78770 56180
rect 78190 56120 78200 56160
rect 78770 56140 78830 56150
rect 78920 56120 78980 56130
rect 77700 56110 77780 56120
rect 78120 56110 78200 56120
rect 78540 56110 78620 56120
rect 77700 56100 77710 56110
rect 77560 56070 77710 56100
rect 77500 56050 77560 56060
rect 77700 56050 77710 56070
rect 77770 56050 77780 56110
rect 73550 56040 73630 56050
rect 77700 56040 77780 56050
rect 78540 56050 78550 56110
rect 78610 56100 78620 56110
rect 78610 56070 78920 56100
rect 78610 56050 78620 56070
rect 78920 56050 78980 56060
rect 78540 56040 78620 56050
rect 53160 56020 53260 56030
rect 53160 55950 53180 56020
rect 53250 55950 53260 56020
rect 53160 55910 53260 55950
rect 53160 55840 53180 55910
rect 53250 55840 53260 55910
rect 53160 55820 53260 55840
rect 58150 56020 58250 56030
rect 58150 55950 58170 56020
rect 58240 55950 58250 56020
rect 58150 55910 58250 55950
rect 58150 55840 58170 55910
rect 58240 55840 58250 55910
rect 58150 55820 58250 55840
rect 63140 56020 63240 56030
rect 63140 55950 63160 56020
rect 63230 55950 63240 56020
rect 63140 55910 63240 55950
rect 63140 55840 63160 55910
rect 63230 55840 63240 55910
rect 63140 55820 63240 55840
rect 68130 56020 68230 56030
rect 68130 55950 68150 56020
rect 68220 55950 68230 56020
rect 68130 55910 68230 55950
rect 68130 55840 68150 55910
rect 68220 55840 68230 55910
rect 68130 55820 68230 55840
rect 73120 56020 73220 56030
rect 73120 55950 73140 56020
rect 73210 55950 73220 56020
rect 73120 55910 73220 55950
rect 73120 55840 73140 55910
rect 73210 55840 73220 55910
rect 73120 55820 73220 55840
rect 78110 56020 78210 56030
rect 78110 55950 78130 56020
rect 78200 55950 78210 56020
rect 78110 55910 78210 55950
rect 78110 55840 78130 55910
rect 78200 55840 78210 55910
rect 78110 55820 78210 55840
rect 52170 55800 52250 55810
rect 52170 55740 52180 55800
rect 52240 55790 52250 55800
rect 52750 55800 52830 55810
rect 52750 55790 52760 55800
rect 52240 55760 52760 55790
rect 52240 55740 52250 55760
rect 52170 55730 52250 55740
rect 52750 55740 52760 55760
rect 52820 55740 52830 55800
rect 53590 55800 53670 55810
rect 53590 55740 53600 55800
rect 53660 55790 53670 55800
rect 54330 55800 54410 55810
rect 54330 55790 54340 55800
rect 53660 55760 54340 55790
rect 53660 55740 53670 55760
rect 52750 55730 52830 55740
rect 53170 55730 53250 55740
rect 53590 55730 53670 55740
rect 54330 55740 54340 55760
rect 54400 55740 54410 55800
rect 54330 55730 54410 55740
rect 57160 55800 57240 55810
rect 57160 55740 57170 55800
rect 57230 55790 57240 55800
rect 57740 55800 57820 55810
rect 57740 55790 57750 55800
rect 57230 55760 57750 55790
rect 57230 55740 57240 55760
rect 57160 55730 57240 55740
rect 57740 55740 57750 55760
rect 57810 55740 57820 55800
rect 58580 55800 58660 55810
rect 58580 55740 58590 55800
rect 58650 55790 58660 55800
rect 59320 55800 59400 55810
rect 59320 55790 59330 55800
rect 58650 55760 59330 55790
rect 58650 55740 58660 55760
rect 57740 55730 57820 55740
rect 58160 55730 58240 55740
rect 58580 55730 58660 55740
rect 59320 55740 59330 55760
rect 59390 55740 59400 55800
rect 59320 55730 59400 55740
rect 62390 55800 62470 55810
rect 62390 55740 62400 55800
rect 62460 55790 62470 55800
rect 62730 55800 62810 55810
rect 62730 55790 62740 55800
rect 62460 55760 62740 55790
rect 62460 55740 62470 55760
rect 62390 55730 62470 55740
rect 62730 55740 62740 55760
rect 62800 55740 62810 55800
rect 63570 55800 63650 55810
rect 63570 55740 63580 55800
rect 63640 55790 63650 55800
rect 64070 55800 64150 55810
rect 64070 55790 64080 55800
rect 63640 55760 64080 55790
rect 63640 55740 63650 55760
rect 62730 55730 62810 55740
rect 63150 55730 63230 55740
rect 63570 55730 63650 55740
rect 64070 55740 64080 55760
rect 64140 55740 64150 55800
rect 64070 55730 64150 55740
rect 67380 55800 67460 55810
rect 67380 55740 67390 55800
rect 67450 55790 67460 55800
rect 67720 55800 67800 55810
rect 67720 55790 67730 55800
rect 67450 55760 67730 55790
rect 67450 55740 67460 55760
rect 67380 55730 67460 55740
rect 67720 55740 67730 55760
rect 67790 55740 67800 55800
rect 68560 55800 68640 55810
rect 68560 55740 68570 55800
rect 68630 55790 68640 55800
rect 69060 55800 69140 55810
rect 69060 55790 69070 55800
rect 68630 55760 69070 55790
rect 68630 55740 68640 55760
rect 67720 55730 67800 55740
rect 68140 55730 68220 55740
rect 68560 55730 68640 55740
rect 69060 55740 69070 55760
rect 69130 55740 69140 55800
rect 69060 55730 69140 55740
rect 72490 55800 72570 55810
rect 72490 55740 72500 55800
rect 72560 55790 72570 55800
rect 72710 55800 72790 55810
rect 72710 55790 72720 55800
rect 72560 55760 72720 55790
rect 72560 55740 72570 55760
rect 72490 55730 72570 55740
rect 72710 55740 72720 55760
rect 72780 55740 72790 55800
rect 73550 55800 73630 55810
rect 73550 55740 73560 55800
rect 73620 55790 73630 55800
rect 73930 55800 74010 55810
rect 73930 55790 73940 55800
rect 73620 55760 73940 55790
rect 73620 55740 73630 55760
rect 72710 55730 72790 55740
rect 73130 55730 73210 55740
rect 73550 55730 73630 55740
rect 73930 55740 73940 55760
rect 74000 55740 74010 55800
rect 73930 55730 74010 55740
rect 77480 55800 77560 55810
rect 77480 55740 77490 55800
rect 77550 55790 77560 55800
rect 77700 55800 77780 55810
rect 77700 55790 77710 55800
rect 77550 55760 77710 55790
rect 77550 55740 77560 55760
rect 77480 55730 77560 55740
rect 77700 55740 77710 55760
rect 77770 55740 77780 55800
rect 78540 55800 78620 55810
rect 78540 55740 78550 55800
rect 78610 55790 78620 55800
rect 78920 55800 79000 55810
rect 78920 55790 78930 55800
rect 78610 55760 78930 55790
rect 78610 55740 78620 55760
rect 77700 55730 77780 55740
rect 78120 55730 78200 55740
rect 78540 55730 78620 55740
rect 78920 55740 78930 55760
rect 78990 55740 79000 55800
rect 78920 55730 79000 55740
rect 53170 55670 53180 55730
rect 53240 55690 53250 55730
rect 53240 55680 53940 55690
rect 53240 55670 53880 55680
rect 53170 55660 53880 55670
rect 58160 55670 58170 55730
rect 58230 55690 58240 55730
rect 58230 55680 58930 55690
rect 58230 55670 58870 55680
rect 58160 55660 58870 55670
rect 53880 55610 53940 55620
rect 63150 55670 63160 55730
rect 63220 55690 63230 55730
rect 63220 55680 63920 55690
rect 63220 55670 63860 55680
rect 63150 55660 63860 55670
rect 58870 55610 58930 55620
rect 68140 55670 68150 55730
rect 68210 55690 68220 55730
rect 68210 55680 68910 55690
rect 68210 55670 68850 55680
rect 68140 55660 68850 55670
rect 63860 55610 63920 55620
rect 73130 55670 73140 55730
rect 73200 55690 73210 55730
rect 73200 55680 73900 55690
rect 73200 55670 73840 55680
rect 73130 55660 73840 55670
rect 68850 55610 68910 55620
rect 78120 55670 78130 55730
rect 78190 55690 78200 55730
rect 78190 55680 78890 55690
rect 78190 55670 78830 55680
rect 78120 55660 78830 55670
rect 73840 55610 73900 55620
rect 78830 55610 78890 55620
rect 49580 54610 49660 54620
rect 49580 54550 49590 54610
rect 49650 54550 49660 54610
rect 49580 54540 49660 54550
rect 48830 54500 48890 54510
rect 48180 54470 48830 54480
rect 44710 54440 44830 54470
rect 43840 54430 43900 54440
rect 41850 54400 41910 54410
rect 42770 54400 42850 54410
rect 43190 54400 43270 54410
rect 43610 54400 43690 54410
rect 42770 54390 42780 54400
rect 41910 54360 42780 54390
rect 41850 54330 41910 54340
rect 42770 54340 42780 54360
rect 42840 54340 42850 54400
rect 42770 54330 42850 54340
rect 43610 54340 43620 54400
rect 43680 54390 43690 54400
rect 44710 54400 44770 54410
rect 43680 54360 44710 54390
rect 43680 54340 43690 54360
rect 43610 54330 43690 54340
rect 44710 54330 44770 54340
rect 43180 54310 43280 54320
rect 41790 54270 41910 54300
rect 37780 54090 37860 54100
rect 37780 54080 37790 54090
rect 36890 54050 37790 54080
rect 3270 53960 3280 54020
rect 3340 53980 3350 54020
rect 3340 53970 4040 53980
rect 3340 53960 3980 53970
rect 3270 53950 3980 53960
rect 8260 53960 8270 54020
rect 8330 53980 8340 54020
rect 8330 53970 9030 53980
rect 8330 53960 8970 53970
rect 8260 53950 8970 53960
rect 3980 53900 4040 53910
rect 13250 53960 13260 54020
rect 13320 53980 13330 54020
rect 13320 53970 14020 53980
rect 13320 53960 13960 53970
rect 13250 53950 13960 53960
rect 8970 53900 9030 53910
rect 18240 53960 18250 54020
rect 18310 53980 18320 54020
rect 18310 53970 19010 53980
rect 18310 53960 18950 53970
rect 18240 53950 18950 53960
rect 13960 53900 14020 53910
rect 23230 53960 23240 54020
rect 23300 53980 23310 54020
rect 23300 53970 24000 53980
rect 23300 53960 23940 53970
rect 23230 53950 23940 53960
rect 18950 53900 19010 53910
rect 28220 53960 28230 54020
rect 28290 53980 28300 54020
rect 28290 53970 28990 53980
rect 28290 53960 28930 53970
rect 28220 53950 28930 53960
rect 23940 53900 24000 53910
rect 33210 53960 33220 54020
rect 33280 53980 33290 54020
rect 33280 53970 33980 53980
rect 33280 53960 33920 53970
rect 33210 53950 33920 53960
rect 28930 53900 28990 53910
rect 33920 53900 33980 53910
rect 3920 52790 3980 52800
rect 3270 52760 3920 52770
rect 2650 52700 2710 52710
rect 3270 52700 3280 52760
rect 3340 52740 3920 52760
rect 3340 52700 3350 52740
rect 8910 52790 8970 52800
rect 3920 52720 3980 52730
rect 8260 52760 8910 52770
rect 4070 52700 4130 52710
rect 2850 52690 2930 52700
rect 3270 52690 3350 52700
rect 3690 52690 3770 52700
rect 2850 52680 2860 52690
rect 2710 52650 2860 52680
rect 2650 52630 2710 52640
rect 2850 52630 2860 52650
rect 2920 52630 2930 52690
rect 2850 52620 2930 52630
rect 3690 52630 3700 52690
rect 3760 52680 3770 52690
rect 3760 52650 4070 52680
rect 3760 52630 3770 52650
rect 4070 52630 4130 52640
rect 7640 52700 7700 52710
rect 8260 52700 8270 52760
rect 8330 52740 8910 52760
rect 8330 52700 8340 52740
rect 13900 52790 13960 52800
rect 8910 52720 8970 52730
rect 13250 52760 13900 52770
rect 9060 52700 9120 52710
rect 7840 52690 7920 52700
rect 8260 52690 8340 52700
rect 8680 52690 8760 52700
rect 7840 52680 7850 52690
rect 7700 52650 7850 52680
rect 7640 52630 7700 52640
rect 7840 52630 7850 52650
rect 7910 52630 7920 52690
rect 3690 52620 3770 52630
rect 7840 52620 7920 52630
rect 8680 52630 8690 52690
rect 8750 52680 8760 52690
rect 8750 52650 9060 52680
rect 8750 52630 8760 52650
rect 9060 52630 9120 52640
rect 12510 52700 12570 52710
rect 13250 52700 13260 52760
rect 13320 52740 13900 52760
rect 13320 52700 13330 52740
rect 18890 52790 18950 52800
rect 13900 52720 13960 52730
rect 18240 52760 18890 52770
rect 14170 52700 14230 52710
rect 12830 52690 12910 52700
rect 13250 52690 13330 52700
rect 13670 52690 13750 52700
rect 12830 52680 12840 52690
rect 12570 52650 12840 52680
rect 12510 52630 12570 52640
rect 12830 52630 12840 52650
rect 12900 52630 12910 52690
rect 8680 52620 8760 52630
rect 12830 52620 12910 52630
rect 13670 52630 13680 52690
rect 13740 52680 13750 52690
rect 13740 52650 14170 52680
rect 13740 52630 13750 52650
rect 14170 52630 14230 52640
rect 17500 52700 17560 52710
rect 18240 52700 18250 52760
rect 18310 52740 18890 52760
rect 18310 52700 18320 52740
rect 23880 52790 23940 52800
rect 18890 52720 18950 52730
rect 23230 52760 23880 52770
rect 19160 52700 19220 52710
rect 17820 52690 17900 52700
rect 18240 52690 18320 52700
rect 18660 52690 18740 52700
rect 17820 52680 17830 52690
rect 17560 52650 17830 52680
rect 17500 52630 17560 52640
rect 17820 52630 17830 52650
rect 17890 52630 17900 52690
rect 13670 52620 13750 52630
rect 17820 52620 17900 52630
rect 18660 52630 18670 52690
rect 18730 52680 18740 52690
rect 18730 52650 19160 52680
rect 18730 52630 18740 52650
rect 19160 52630 19220 52640
rect 22250 52700 22310 52710
rect 23230 52700 23240 52760
rect 23300 52740 23880 52760
rect 23300 52700 23310 52740
rect 28870 52790 28930 52800
rect 23880 52720 23940 52730
rect 28220 52760 28870 52770
rect 24390 52700 24450 52710
rect 22810 52690 22890 52700
rect 23230 52690 23310 52700
rect 23650 52690 23730 52700
rect 22810 52680 22820 52690
rect 22310 52650 22820 52680
rect 22250 52630 22310 52640
rect 22810 52630 22820 52650
rect 22880 52630 22890 52690
rect 18660 52620 18740 52630
rect 22810 52620 22890 52630
rect 23650 52630 23660 52690
rect 23720 52680 23730 52690
rect 23720 52650 24390 52680
rect 23720 52630 23730 52650
rect 24390 52630 24450 52640
rect 27240 52700 27300 52710
rect 28220 52700 28230 52760
rect 28290 52740 28870 52760
rect 28290 52700 28300 52740
rect 33860 52790 33920 52800
rect 28870 52720 28930 52730
rect 33210 52760 33860 52770
rect 29380 52700 29440 52710
rect 27800 52690 27880 52700
rect 28220 52690 28300 52700
rect 28640 52690 28720 52700
rect 27800 52680 27810 52690
rect 27300 52650 27810 52680
rect 27240 52630 27300 52640
rect 27800 52630 27810 52650
rect 27870 52630 27880 52690
rect 23650 52620 23730 52630
rect 27800 52620 27880 52630
rect 28640 52630 28650 52690
rect 28710 52680 28720 52690
rect 28710 52650 29380 52680
rect 28710 52630 28720 52650
rect 29380 52630 29440 52640
rect 31990 52700 32050 52710
rect 33210 52700 33220 52760
rect 33280 52740 33860 52760
rect 33280 52700 33290 52740
rect 33860 52720 33920 52730
rect 34610 52700 34670 52710
rect 32790 52690 32870 52700
rect 33210 52690 33290 52700
rect 33630 52690 33710 52700
rect 32790 52680 32800 52690
rect 32050 52650 32800 52680
rect 31990 52630 32050 52640
rect 32790 52630 32800 52650
rect 32860 52630 32870 52690
rect 28640 52620 28720 52630
rect 32790 52620 32870 52630
rect 33630 52630 33640 52690
rect 33700 52680 33710 52690
rect 33700 52650 34610 52680
rect 33700 52630 33710 52650
rect 34610 52630 34670 52640
rect 33630 52620 33710 52630
rect 3260 52600 3360 52610
rect 3260 52530 3280 52600
rect 3350 52530 3360 52600
rect 3260 52490 3360 52530
rect 3260 52420 3280 52490
rect 3350 52420 3360 52490
rect 3260 52400 3360 52420
rect 8250 52600 8350 52610
rect 8250 52530 8270 52600
rect 8340 52530 8350 52600
rect 8250 52490 8350 52530
rect 8250 52420 8270 52490
rect 8340 52420 8350 52490
rect 8250 52400 8350 52420
rect 13240 52600 13340 52610
rect 13240 52530 13260 52600
rect 13330 52530 13340 52600
rect 13240 52490 13340 52530
rect 13240 52420 13260 52490
rect 13330 52420 13340 52490
rect 13240 52400 13340 52420
rect 18230 52600 18330 52610
rect 18230 52530 18250 52600
rect 18320 52530 18330 52600
rect 18230 52490 18330 52530
rect 18230 52420 18250 52490
rect 18320 52420 18330 52490
rect 18230 52400 18330 52420
rect 23220 52600 23320 52610
rect 23220 52530 23240 52600
rect 23310 52530 23320 52600
rect 23220 52490 23320 52530
rect 23220 52420 23240 52490
rect 23310 52420 23320 52490
rect 23220 52400 23320 52420
rect 28210 52600 28310 52610
rect 28210 52530 28230 52600
rect 28300 52530 28310 52600
rect 28210 52490 28310 52530
rect 28210 52420 28230 52490
rect 28300 52420 28310 52490
rect 28210 52400 28310 52420
rect 33200 52600 33300 52610
rect 33200 52530 33220 52600
rect 33290 52530 33300 52600
rect 33200 52490 33300 52530
rect 33200 52420 33220 52490
rect 33290 52420 33300 52490
rect 33200 52400 33300 52420
rect 2630 52380 2710 52390
rect 2630 52320 2640 52380
rect 2700 52370 2710 52380
rect 2850 52380 2930 52390
rect 2850 52370 2860 52380
rect 2700 52340 2860 52370
rect 2700 52320 2710 52340
rect 2630 52310 2710 52320
rect 2850 52320 2860 52340
rect 2920 52320 2930 52380
rect 3690 52380 3770 52390
rect 3690 52320 3700 52380
rect 3760 52370 3770 52380
rect 4070 52380 4150 52390
rect 4070 52370 4080 52380
rect 3760 52340 4080 52370
rect 3760 52320 3770 52340
rect 2850 52310 2930 52320
rect 3270 52310 3350 52320
rect 3690 52310 3770 52320
rect 4070 52320 4080 52340
rect 4140 52320 4150 52380
rect 4070 52310 4150 52320
rect 7620 52380 7700 52390
rect 7620 52320 7630 52380
rect 7690 52370 7700 52380
rect 7840 52380 7920 52390
rect 7840 52370 7850 52380
rect 7690 52340 7850 52370
rect 7690 52320 7700 52340
rect 7620 52310 7700 52320
rect 7840 52320 7850 52340
rect 7910 52320 7920 52380
rect 8680 52380 8760 52390
rect 8680 52320 8690 52380
rect 8750 52370 8760 52380
rect 9060 52380 9140 52390
rect 9060 52370 9070 52380
rect 8750 52340 9070 52370
rect 8750 52320 8760 52340
rect 7840 52310 7920 52320
rect 8260 52310 8340 52320
rect 8680 52310 8760 52320
rect 9060 52320 9070 52340
rect 9130 52320 9140 52380
rect 9060 52310 9140 52320
rect 12490 52380 12570 52390
rect 12490 52320 12500 52380
rect 12560 52370 12570 52380
rect 12830 52380 12910 52390
rect 12830 52370 12840 52380
rect 12560 52340 12840 52370
rect 12560 52320 12570 52340
rect 12490 52310 12570 52320
rect 12830 52320 12840 52340
rect 12900 52320 12910 52380
rect 13670 52380 13750 52390
rect 13670 52320 13680 52380
rect 13740 52370 13750 52380
rect 14170 52380 14250 52390
rect 14170 52370 14180 52380
rect 13740 52340 14180 52370
rect 13740 52320 13750 52340
rect 12830 52310 12910 52320
rect 13250 52310 13330 52320
rect 13670 52310 13750 52320
rect 14170 52320 14180 52340
rect 14240 52320 14250 52380
rect 14170 52310 14250 52320
rect 17480 52380 17560 52390
rect 17480 52320 17490 52380
rect 17550 52370 17560 52380
rect 17820 52380 17900 52390
rect 17820 52370 17830 52380
rect 17550 52340 17830 52370
rect 17550 52320 17560 52340
rect 17480 52310 17560 52320
rect 17820 52320 17830 52340
rect 17890 52320 17900 52380
rect 18660 52380 18740 52390
rect 18660 52320 18670 52380
rect 18730 52370 18740 52380
rect 19160 52380 19240 52390
rect 19160 52370 19170 52380
rect 18730 52340 19170 52370
rect 18730 52320 18740 52340
rect 17820 52310 17900 52320
rect 18240 52310 18320 52320
rect 18660 52310 18740 52320
rect 19160 52320 19170 52340
rect 19230 52320 19240 52380
rect 19160 52310 19240 52320
rect 22230 52380 22310 52390
rect 22230 52320 22240 52380
rect 22300 52370 22310 52380
rect 22810 52380 22890 52390
rect 22810 52370 22820 52380
rect 22300 52340 22820 52370
rect 22300 52320 22310 52340
rect 22230 52310 22310 52320
rect 22810 52320 22820 52340
rect 22880 52320 22890 52380
rect 23650 52380 23730 52390
rect 23650 52320 23660 52380
rect 23720 52370 23730 52380
rect 24390 52380 24470 52390
rect 24390 52370 24400 52380
rect 23720 52340 24400 52370
rect 23720 52320 23730 52340
rect 22810 52310 22890 52320
rect 23230 52310 23310 52320
rect 23650 52310 23730 52320
rect 24390 52320 24400 52340
rect 24460 52320 24470 52380
rect 24390 52310 24470 52320
rect 27220 52380 27300 52390
rect 27220 52320 27230 52380
rect 27290 52370 27300 52380
rect 27800 52380 27880 52390
rect 27800 52370 27810 52380
rect 27290 52340 27810 52370
rect 27290 52320 27300 52340
rect 27220 52310 27300 52320
rect 27800 52320 27810 52340
rect 27870 52320 27880 52380
rect 28640 52380 28720 52390
rect 28640 52320 28650 52380
rect 28710 52370 28720 52380
rect 29380 52380 29460 52390
rect 29380 52370 29390 52380
rect 28710 52340 29390 52370
rect 28710 52320 28720 52340
rect 27800 52310 27880 52320
rect 28220 52310 28300 52320
rect 28640 52310 28720 52320
rect 29380 52320 29390 52340
rect 29450 52320 29460 52380
rect 29380 52310 29460 52320
rect 31970 52380 32050 52390
rect 31970 52320 31980 52380
rect 32040 52370 32050 52380
rect 32790 52380 32870 52390
rect 32790 52370 32800 52380
rect 32040 52340 32800 52370
rect 32040 52320 32050 52340
rect 31970 52310 32050 52320
rect 32790 52320 32800 52340
rect 32860 52320 32870 52380
rect 33630 52380 33710 52390
rect 33630 52320 33640 52380
rect 33700 52370 33710 52380
rect 34610 52380 34690 52390
rect 34610 52370 34620 52380
rect 33700 52340 34620 52370
rect 33700 52320 33710 52340
rect 32790 52310 32870 52320
rect 33210 52310 33290 52320
rect 33630 52310 33710 52320
rect 34610 52320 34620 52340
rect 34680 52320 34690 52380
rect 34610 52310 34690 52320
rect 3270 52250 3280 52310
rect 3340 52270 3350 52310
rect 3340 52260 4040 52270
rect 3340 52250 3980 52260
rect 3270 52240 3980 52250
rect 8260 52250 8270 52310
rect 8330 52270 8340 52310
rect 8330 52260 9030 52270
rect 8330 52250 8970 52260
rect 8260 52240 8970 52250
rect 3980 52190 4040 52200
rect 13250 52250 13260 52310
rect 13320 52270 13330 52310
rect 13320 52260 14020 52270
rect 13320 52250 13960 52260
rect 13250 52240 13960 52250
rect 8970 52190 9030 52200
rect 18240 52250 18250 52310
rect 18310 52270 18320 52310
rect 18310 52260 19010 52270
rect 18310 52250 18950 52260
rect 18240 52240 18950 52250
rect 13960 52190 14020 52200
rect 23230 52250 23240 52310
rect 23300 52270 23310 52310
rect 23300 52260 24000 52270
rect 23300 52250 23940 52260
rect 23230 52240 23940 52250
rect 18950 52190 19010 52200
rect 28220 52250 28230 52310
rect 28290 52270 28300 52310
rect 28290 52260 28990 52270
rect 28290 52250 28930 52260
rect 28220 52240 28930 52250
rect 23940 52190 24000 52200
rect 28930 52190 28990 52200
rect 3920 51080 3980 51090
rect 3270 51050 3920 51060
rect 2650 50990 2710 51000
rect 3270 50990 3280 51050
rect 3340 51030 3920 51050
rect 3340 50990 3350 51030
rect 8910 51080 8970 51090
rect 3920 51010 3980 51020
rect 8260 51050 8910 51060
rect 4070 50990 4130 51000
rect 2850 50980 2930 50990
rect 3270 50980 3350 50990
rect 3690 50980 3770 50990
rect 2850 50970 2860 50980
rect 2710 50940 2860 50970
rect 2650 50920 2710 50930
rect 2850 50920 2860 50940
rect 2920 50920 2930 50980
rect 2850 50910 2930 50920
rect 3690 50920 3700 50980
rect 3760 50970 3770 50980
rect 3760 50940 4070 50970
rect 3760 50920 3770 50940
rect 4070 50920 4130 50930
rect 7640 50990 7700 51000
rect 8260 50990 8270 51050
rect 8330 51030 8910 51050
rect 8330 50990 8340 51030
rect 13900 51080 13960 51090
rect 8910 51010 8970 51020
rect 13250 51050 13900 51060
rect 9060 50990 9120 51000
rect 7840 50980 7920 50990
rect 8260 50980 8340 50990
rect 8680 50980 8760 50990
rect 7840 50970 7850 50980
rect 7700 50940 7850 50970
rect 7640 50920 7700 50930
rect 7840 50920 7850 50940
rect 7910 50920 7920 50980
rect 3690 50910 3770 50920
rect 7840 50910 7920 50920
rect 8680 50920 8690 50980
rect 8750 50970 8760 50980
rect 8750 50940 9060 50970
rect 8750 50920 8760 50940
rect 9060 50920 9120 50930
rect 12510 50990 12570 51000
rect 13250 50990 13260 51050
rect 13320 51030 13900 51050
rect 13320 50990 13330 51030
rect 18890 51080 18950 51090
rect 13900 51010 13960 51020
rect 18240 51050 18890 51060
rect 14170 50990 14230 51000
rect 12830 50980 12910 50990
rect 13250 50980 13330 50990
rect 13670 50980 13750 50990
rect 12830 50970 12840 50980
rect 12570 50940 12840 50970
rect 12510 50920 12570 50930
rect 12830 50920 12840 50940
rect 12900 50920 12910 50980
rect 8680 50910 8760 50920
rect 12830 50910 12910 50920
rect 13670 50920 13680 50980
rect 13740 50970 13750 50980
rect 13740 50940 14170 50970
rect 13740 50920 13750 50940
rect 14170 50920 14230 50930
rect 17500 50990 17560 51000
rect 18240 50990 18250 51050
rect 18310 51030 18890 51050
rect 18310 50990 18320 51030
rect 23880 51080 23940 51090
rect 18890 51010 18950 51020
rect 23230 51050 23880 51060
rect 19160 50990 19220 51000
rect 17820 50980 17900 50990
rect 18240 50980 18320 50990
rect 18660 50980 18740 50990
rect 17820 50970 17830 50980
rect 17560 50940 17830 50970
rect 17500 50920 17560 50930
rect 17820 50920 17830 50940
rect 17890 50920 17900 50980
rect 13670 50910 13750 50920
rect 17820 50910 17900 50920
rect 18660 50920 18670 50980
rect 18730 50970 18740 50980
rect 18730 50940 19160 50970
rect 18730 50920 18740 50940
rect 19160 50920 19220 50930
rect 22250 50990 22310 51000
rect 23230 50990 23240 51050
rect 23300 51030 23880 51050
rect 23300 50990 23310 51030
rect 28870 51080 28930 51090
rect 23880 51010 23940 51020
rect 28220 51050 28870 51060
rect 24390 50990 24450 51000
rect 22810 50980 22890 50990
rect 23230 50980 23310 50990
rect 23650 50980 23730 50990
rect 22810 50970 22820 50980
rect 22310 50940 22820 50970
rect 22250 50920 22310 50930
rect 22810 50920 22820 50940
rect 22880 50920 22890 50980
rect 18660 50910 18740 50920
rect 22810 50910 22890 50920
rect 23650 50920 23660 50980
rect 23720 50970 23730 50980
rect 23720 50940 24390 50970
rect 23720 50920 23730 50940
rect 24390 50920 24450 50930
rect 27240 50990 27300 51000
rect 28220 50990 28230 51050
rect 28290 51030 28870 51050
rect 28290 50990 28300 51030
rect 28870 51010 28930 51020
rect 29380 50990 29440 51000
rect 27800 50980 27880 50990
rect 28220 50980 28300 50990
rect 28640 50980 28720 50990
rect 27800 50970 27810 50980
rect 27300 50940 27810 50970
rect 27240 50920 27300 50930
rect 27800 50920 27810 50940
rect 27870 50920 27880 50980
rect 23650 50910 23730 50920
rect 27800 50910 27880 50920
rect 28640 50920 28650 50980
rect 28710 50970 28720 50980
rect 28710 50940 29380 50970
rect 28710 50920 28720 50940
rect 29380 50920 29440 50930
rect 28640 50910 28720 50920
rect 3260 50890 3360 50900
rect 3260 50820 3280 50890
rect 3350 50820 3360 50890
rect 3260 50780 3360 50820
rect 3260 50710 3280 50780
rect 3350 50710 3360 50780
rect 3260 50690 3360 50710
rect 8250 50890 8350 50900
rect 8250 50820 8270 50890
rect 8340 50820 8350 50890
rect 8250 50780 8350 50820
rect 8250 50710 8270 50780
rect 8340 50710 8350 50780
rect 8250 50690 8350 50710
rect 13240 50890 13340 50900
rect 13240 50820 13260 50890
rect 13330 50820 13340 50890
rect 13240 50780 13340 50820
rect 13240 50710 13260 50780
rect 13330 50710 13340 50780
rect 13240 50690 13340 50710
rect 18230 50890 18330 50900
rect 18230 50820 18250 50890
rect 18320 50820 18330 50890
rect 18230 50780 18330 50820
rect 18230 50710 18250 50780
rect 18320 50710 18330 50780
rect 18230 50690 18330 50710
rect 23220 50890 23320 50900
rect 23220 50820 23240 50890
rect 23310 50820 23320 50890
rect 23220 50780 23320 50820
rect 23220 50710 23240 50780
rect 23310 50710 23320 50780
rect 23220 50690 23320 50710
rect 28210 50890 28310 50900
rect 28210 50820 28230 50890
rect 28300 50820 28310 50890
rect 28210 50780 28310 50820
rect 28210 50710 28230 50780
rect 28300 50710 28310 50780
rect 28210 50690 28310 50710
rect 2630 50670 2710 50680
rect 2630 50610 2640 50670
rect 2700 50660 2710 50670
rect 2850 50670 2930 50680
rect 2850 50660 2860 50670
rect 2700 50630 2860 50660
rect 2700 50610 2710 50630
rect 2630 50600 2710 50610
rect 2850 50610 2860 50630
rect 2920 50610 2930 50670
rect 3690 50670 3770 50680
rect 3690 50610 3700 50670
rect 3760 50660 3770 50670
rect 4070 50670 4150 50680
rect 4070 50660 4080 50670
rect 3760 50630 4080 50660
rect 3760 50610 3770 50630
rect 2850 50600 2930 50610
rect 3270 50600 3350 50610
rect 3690 50600 3770 50610
rect 4070 50610 4080 50630
rect 4140 50610 4150 50670
rect 4070 50600 4150 50610
rect 7620 50670 7700 50680
rect 7620 50610 7630 50670
rect 7690 50660 7700 50670
rect 7840 50670 7920 50680
rect 7840 50660 7850 50670
rect 7690 50630 7850 50660
rect 7690 50610 7700 50630
rect 7620 50600 7700 50610
rect 7840 50610 7850 50630
rect 7910 50610 7920 50670
rect 8680 50670 8760 50680
rect 8680 50610 8690 50670
rect 8750 50660 8760 50670
rect 9060 50670 9140 50680
rect 9060 50660 9070 50670
rect 8750 50630 9070 50660
rect 8750 50610 8760 50630
rect 7840 50600 7920 50610
rect 8260 50600 8340 50610
rect 8680 50600 8760 50610
rect 9060 50610 9070 50630
rect 9130 50610 9140 50670
rect 9060 50600 9140 50610
rect 12490 50670 12570 50680
rect 12490 50610 12500 50670
rect 12560 50660 12570 50670
rect 12830 50670 12910 50680
rect 12830 50660 12840 50670
rect 12560 50630 12840 50660
rect 12560 50610 12570 50630
rect 12490 50600 12570 50610
rect 12830 50610 12840 50630
rect 12900 50610 12910 50670
rect 13670 50670 13750 50680
rect 13670 50610 13680 50670
rect 13740 50660 13750 50670
rect 14170 50670 14250 50680
rect 14170 50660 14180 50670
rect 13740 50630 14180 50660
rect 13740 50610 13750 50630
rect 12830 50600 12910 50610
rect 13250 50600 13330 50610
rect 13670 50600 13750 50610
rect 14170 50610 14180 50630
rect 14240 50610 14250 50670
rect 14170 50600 14250 50610
rect 17480 50670 17560 50680
rect 17480 50610 17490 50670
rect 17550 50660 17560 50670
rect 17820 50670 17900 50680
rect 17820 50660 17830 50670
rect 17550 50630 17830 50660
rect 17550 50610 17560 50630
rect 17480 50600 17560 50610
rect 17820 50610 17830 50630
rect 17890 50610 17900 50670
rect 18660 50670 18740 50680
rect 18660 50610 18670 50670
rect 18730 50660 18740 50670
rect 19160 50670 19240 50680
rect 19160 50660 19170 50670
rect 18730 50630 19170 50660
rect 18730 50610 18740 50630
rect 17820 50600 17900 50610
rect 18240 50600 18320 50610
rect 18660 50600 18740 50610
rect 19160 50610 19170 50630
rect 19230 50610 19240 50670
rect 19160 50600 19240 50610
rect 22230 50670 22310 50680
rect 22230 50610 22240 50670
rect 22300 50660 22310 50670
rect 22810 50670 22890 50680
rect 22810 50660 22820 50670
rect 22300 50630 22820 50660
rect 22300 50610 22310 50630
rect 22230 50600 22310 50610
rect 22810 50610 22820 50630
rect 22880 50610 22890 50670
rect 23650 50670 23730 50680
rect 23650 50610 23660 50670
rect 23720 50660 23730 50670
rect 24390 50670 24470 50680
rect 24390 50660 24400 50670
rect 23720 50630 24400 50660
rect 23720 50610 23730 50630
rect 22810 50600 22890 50610
rect 23230 50600 23310 50610
rect 23650 50600 23730 50610
rect 24390 50610 24400 50630
rect 24460 50610 24470 50670
rect 24390 50600 24470 50610
rect 27220 50670 27300 50680
rect 27220 50610 27230 50670
rect 27290 50660 27300 50670
rect 27800 50670 27880 50680
rect 27800 50660 27810 50670
rect 27290 50630 27810 50660
rect 27290 50610 27300 50630
rect 27220 50600 27300 50610
rect 27800 50610 27810 50630
rect 27870 50610 27880 50670
rect 28640 50670 28720 50680
rect 28640 50610 28650 50670
rect 28710 50660 28720 50670
rect 29380 50670 29460 50680
rect 29380 50660 29390 50670
rect 28710 50630 29390 50660
rect 28710 50610 28720 50630
rect 27800 50600 27880 50610
rect 28220 50600 28300 50610
rect 28640 50600 28720 50610
rect 29380 50610 29390 50630
rect 29450 50610 29460 50670
rect 29380 50600 29460 50610
rect 3270 50540 3280 50600
rect 3340 50560 3350 50600
rect 3340 50550 4040 50560
rect 3340 50540 3980 50550
rect 3270 50530 3980 50540
rect 8260 50540 8270 50600
rect 8330 50560 8340 50600
rect 8330 50550 9030 50560
rect 8330 50540 8970 50550
rect 8260 50530 8970 50540
rect 3980 50480 4040 50490
rect 13250 50540 13260 50600
rect 13320 50560 13330 50600
rect 13320 50550 14020 50560
rect 13320 50540 13960 50550
rect 13250 50530 13960 50540
rect 8970 50480 9030 50490
rect 18240 50540 18250 50600
rect 18310 50560 18320 50600
rect 18310 50550 19010 50560
rect 18310 50540 18950 50550
rect 18240 50530 18950 50540
rect 13960 50480 14020 50490
rect 23230 50540 23240 50600
rect 23300 50560 23310 50600
rect 23300 50550 24000 50560
rect 23300 50540 23940 50550
rect 23230 50530 23940 50540
rect 18950 50480 19010 50490
rect 28220 50540 28230 50600
rect 28290 50560 28300 50600
rect 28290 50550 28990 50560
rect 28290 50540 28930 50550
rect 28220 50530 28930 50540
rect 23940 50480 24000 50490
rect 28930 50480 28990 50490
rect 3920 49370 3980 49380
rect 3270 49340 3920 49350
rect 2650 49280 2710 49290
rect 3270 49280 3280 49340
rect 3340 49320 3920 49340
rect 3340 49280 3350 49320
rect 8910 49370 8970 49380
rect 3920 49300 3980 49310
rect 8260 49340 8910 49350
rect 4070 49280 4130 49290
rect 2850 49270 2930 49280
rect 3270 49270 3350 49280
rect 3690 49270 3770 49280
rect 2850 49260 2860 49270
rect 2710 49230 2860 49260
rect 2650 49210 2710 49220
rect 2850 49210 2860 49230
rect 2920 49210 2930 49270
rect 2850 49200 2930 49210
rect 3690 49210 3700 49270
rect 3760 49260 3770 49270
rect 3760 49230 4070 49260
rect 3760 49210 3770 49230
rect 4070 49210 4130 49220
rect 7640 49280 7700 49290
rect 8260 49280 8270 49340
rect 8330 49320 8910 49340
rect 8330 49280 8340 49320
rect 13900 49370 13960 49380
rect 8910 49300 8970 49310
rect 13250 49340 13900 49350
rect 9060 49280 9120 49290
rect 7840 49270 7920 49280
rect 8260 49270 8340 49280
rect 8680 49270 8760 49280
rect 7840 49260 7850 49270
rect 7700 49230 7850 49260
rect 7640 49210 7700 49220
rect 7840 49210 7850 49230
rect 7910 49210 7920 49270
rect 3690 49200 3770 49210
rect 7840 49200 7920 49210
rect 8680 49210 8690 49270
rect 8750 49260 8760 49270
rect 8750 49230 9060 49260
rect 8750 49210 8760 49230
rect 9060 49210 9120 49220
rect 12510 49280 12570 49290
rect 13250 49280 13260 49340
rect 13320 49320 13900 49340
rect 13320 49280 13330 49320
rect 18890 49370 18950 49380
rect 13900 49300 13960 49310
rect 18240 49340 18890 49350
rect 14170 49280 14230 49290
rect 12830 49270 12910 49280
rect 13250 49270 13330 49280
rect 13670 49270 13750 49280
rect 12830 49260 12840 49270
rect 12570 49230 12840 49260
rect 12510 49210 12570 49220
rect 12830 49210 12840 49230
rect 12900 49210 12910 49270
rect 8680 49200 8760 49210
rect 12830 49200 12910 49210
rect 13670 49210 13680 49270
rect 13740 49260 13750 49270
rect 13740 49230 14170 49260
rect 13740 49210 13750 49230
rect 14170 49210 14230 49220
rect 17500 49280 17560 49290
rect 18240 49280 18250 49340
rect 18310 49320 18890 49340
rect 18310 49280 18320 49320
rect 23880 49370 23940 49380
rect 18890 49300 18950 49310
rect 23230 49340 23880 49350
rect 19160 49280 19220 49290
rect 17820 49270 17900 49280
rect 18240 49270 18320 49280
rect 18660 49270 18740 49280
rect 17820 49260 17830 49270
rect 17560 49230 17830 49260
rect 17500 49210 17560 49220
rect 17820 49210 17830 49230
rect 17890 49210 17900 49270
rect 13670 49200 13750 49210
rect 17820 49200 17900 49210
rect 18660 49210 18670 49270
rect 18730 49260 18740 49270
rect 18730 49230 19160 49260
rect 18730 49210 18740 49230
rect 19160 49210 19220 49220
rect 22250 49280 22310 49290
rect 23230 49280 23240 49340
rect 23300 49320 23880 49340
rect 23300 49280 23310 49320
rect 28870 49370 28930 49380
rect 23880 49300 23940 49310
rect 28220 49340 28870 49350
rect 24390 49280 24450 49290
rect 22810 49270 22890 49280
rect 23230 49270 23310 49280
rect 23650 49270 23730 49280
rect 22810 49260 22820 49270
rect 22310 49230 22820 49260
rect 22250 49210 22310 49220
rect 22810 49210 22820 49230
rect 22880 49210 22890 49270
rect 18660 49200 18740 49210
rect 22810 49200 22890 49210
rect 23650 49210 23660 49270
rect 23720 49260 23730 49270
rect 23720 49230 24390 49260
rect 23720 49210 23730 49230
rect 24390 49210 24450 49220
rect 27240 49280 27300 49290
rect 28220 49280 28230 49340
rect 28290 49320 28870 49340
rect 28290 49280 28300 49320
rect 28870 49300 28930 49310
rect 29380 49280 29440 49290
rect 27800 49270 27880 49280
rect 28220 49270 28300 49280
rect 28640 49270 28720 49280
rect 27800 49260 27810 49270
rect 27300 49230 27810 49260
rect 27240 49210 27300 49220
rect 27800 49210 27810 49230
rect 27870 49210 27880 49270
rect 23650 49200 23730 49210
rect 27800 49200 27880 49210
rect 28640 49210 28650 49270
rect 28710 49260 28720 49270
rect 28710 49230 29380 49260
rect 28710 49210 28720 49230
rect 29380 49210 29440 49220
rect 28640 49200 28720 49210
rect 3260 49180 3360 49190
rect 3260 49110 3280 49180
rect 3350 49110 3360 49180
rect 3260 49070 3360 49110
rect 3260 49000 3280 49070
rect 3350 49000 3360 49070
rect 3260 48980 3360 49000
rect 8250 49180 8350 49190
rect 8250 49110 8270 49180
rect 8340 49110 8350 49180
rect 8250 49070 8350 49110
rect 8250 49000 8270 49070
rect 8340 49000 8350 49070
rect 8250 48980 8350 49000
rect 13240 49180 13340 49190
rect 13240 49110 13260 49180
rect 13330 49110 13340 49180
rect 13240 49070 13340 49110
rect 13240 49000 13260 49070
rect 13330 49000 13340 49070
rect 13240 48980 13340 49000
rect 18230 49180 18330 49190
rect 18230 49110 18250 49180
rect 18320 49110 18330 49180
rect 18230 49070 18330 49110
rect 18230 49000 18250 49070
rect 18320 49000 18330 49070
rect 18230 48980 18330 49000
rect 23220 49180 23320 49190
rect 23220 49110 23240 49180
rect 23310 49110 23320 49180
rect 23220 49070 23320 49110
rect 23220 49000 23240 49070
rect 23310 49000 23320 49070
rect 23220 48980 23320 49000
rect 28210 49180 28310 49190
rect 28210 49110 28230 49180
rect 28300 49110 28310 49180
rect 28210 49070 28310 49110
rect 28210 49000 28230 49070
rect 28300 49000 28310 49070
rect 28210 48980 28310 49000
rect 2630 48960 2710 48970
rect 2630 48900 2640 48960
rect 2700 48950 2710 48960
rect 2850 48960 2930 48970
rect 2850 48950 2860 48960
rect 2700 48920 2860 48950
rect 2700 48900 2710 48920
rect 2630 48890 2710 48900
rect 2850 48900 2860 48920
rect 2920 48900 2930 48960
rect 3690 48960 3770 48970
rect 3690 48900 3700 48960
rect 3760 48950 3770 48960
rect 4070 48960 4150 48970
rect 4070 48950 4080 48960
rect 3760 48920 4080 48950
rect 3760 48900 3770 48920
rect 2850 48890 2930 48900
rect 3270 48890 3350 48900
rect 3690 48890 3770 48900
rect 4070 48900 4080 48920
rect 4140 48900 4150 48960
rect 4070 48890 4150 48900
rect 7620 48960 7700 48970
rect 7620 48900 7630 48960
rect 7690 48950 7700 48960
rect 7840 48960 7920 48970
rect 7840 48950 7850 48960
rect 7690 48920 7850 48950
rect 7690 48900 7700 48920
rect 7620 48890 7700 48900
rect 7840 48900 7850 48920
rect 7910 48900 7920 48960
rect 8680 48960 8760 48970
rect 8680 48900 8690 48960
rect 8750 48950 8760 48960
rect 9060 48960 9140 48970
rect 9060 48950 9070 48960
rect 8750 48920 9070 48950
rect 8750 48900 8760 48920
rect 7840 48890 7920 48900
rect 8260 48890 8340 48900
rect 8680 48890 8760 48900
rect 9060 48900 9070 48920
rect 9130 48900 9140 48960
rect 9060 48890 9140 48900
rect 12490 48960 12570 48970
rect 12490 48900 12500 48960
rect 12560 48950 12570 48960
rect 12830 48960 12910 48970
rect 12830 48950 12840 48960
rect 12560 48920 12840 48950
rect 12560 48900 12570 48920
rect 12490 48890 12570 48900
rect 12830 48900 12840 48920
rect 12900 48900 12910 48960
rect 13670 48960 13750 48970
rect 13670 48900 13680 48960
rect 13740 48950 13750 48960
rect 14170 48960 14250 48970
rect 14170 48950 14180 48960
rect 13740 48920 14180 48950
rect 13740 48900 13750 48920
rect 12830 48890 12910 48900
rect 13250 48890 13330 48900
rect 13670 48890 13750 48900
rect 14170 48900 14180 48920
rect 14240 48900 14250 48960
rect 14170 48890 14250 48900
rect 17480 48960 17560 48970
rect 17480 48900 17490 48960
rect 17550 48950 17560 48960
rect 17820 48960 17900 48970
rect 17820 48950 17830 48960
rect 17550 48920 17830 48950
rect 17550 48900 17560 48920
rect 17480 48890 17560 48900
rect 17820 48900 17830 48920
rect 17890 48900 17900 48960
rect 18660 48960 18740 48970
rect 18660 48900 18670 48960
rect 18730 48950 18740 48960
rect 19160 48960 19240 48970
rect 19160 48950 19170 48960
rect 18730 48920 19170 48950
rect 18730 48900 18740 48920
rect 17820 48890 17900 48900
rect 18240 48890 18320 48900
rect 18660 48890 18740 48900
rect 19160 48900 19170 48920
rect 19230 48900 19240 48960
rect 19160 48890 19240 48900
rect 22230 48960 22310 48970
rect 22230 48900 22240 48960
rect 22300 48950 22310 48960
rect 22810 48960 22890 48970
rect 22810 48950 22820 48960
rect 22300 48920 22820 48950
rect 22300 48900 22310 48920
rect 22230 48890 22310 48900
rect 22810 48900 22820 48920
rect 22880 48900 22890 48960
rect 23650 48960 23730 48970
rect 23650 48900 23660 48960
rect 23720 48950 23730 48960
rect 24390 48960 24470 48970
rect 24390 48950 24400 48960
rect 23720 48920 24400 48950
rect 23720 48900 23730 48920
rect 22810 48890 22890 48900
rect 23230 48890 23310 48900
rect 23650 48890 23730 48900
rect 24390 48900 24400 48920
rect 24460 48900 24470 48960
rect 24390 48890 24470 48900
rect 27220 48960 27300 48970
rect 27220 48900 27230 48960
rect 27290 48950 27300 48960
rect 27800 48960 27880 48970
rect 27800 48950 27810 48960
rect 27290 48920 27810 48950
rect 27290 48900 27300 48920
rect 27220 48890 27300 48900
rect 27800 48900 27810 48920
rect 27870 48900 27880 48960
rect 28640 48960 28720 48970
rect 28640 48900 28650 48960
rect 28710 48950 28720 48960
rect 29380 48960 29460 48970
rect 29380 48950 29390 48960
rect 28710 48920 29390 48950
rect 28710 48900 28720 48920
rect 27800 48890 27880 48900
rect 28220 48890 28300 48900
rect 28640 48890 28720 48900
rect 29380 48900 29390 48920
rect 29450 48900 29460 48960
rect 29380 48890 29460 48900
rect 3270 48830 3280 48890
rect 3340 48850 3350 48890
rect 3340 48840 4040 48850
rect 3340 48830 3980 48840
rect 3270 48820 3980 48830
rect 8260 48830 8270 48890
rect 8330 48850 8340 48890
rect 8330 48840 9030 48850
rect 8330 48830 8970 48840
rect 8260 48820 8970 48830
rect 3980 48770 4040 48780
rect 13250 48830 13260 48890
rect 13320 48850 13330 48890
rect 13320 48840 14020 48850
rect 13320 48830 13960 48840
rect 13250 48820 13960 48830
rect 8970 48770 9030 48780
rect 18240 48830 18250 48890
rect 18310 48850 18320 48890
rect 18310 48840 19010 48850
rect 18310 48830 18950 48840
rect 18240 48820 18950 48830
rect 13960 48770 14020 48780
rect 18950 48770 19010 48780
rect 3920 47660 3980 47670
rect 3270 47630 3920 47640
rect 2650 47570 2710 47580
rect 3270 47570 3280 47630
rect 3340 47610 3920 47630
rect 3340 47570 3350 47610
rect 8910 47660 8970 47670
rect 3920 47590 3980 47600
rect 8260 47630 8910 47640
rect 4070 47570 4130 47580
rect 2850 47560 2930 47570
rect 3270 47560 3350 47570
rect 3690 47560 3770 47570
rect 2850 47550 2860 47560
rect 2710 47520 2860 47550
rect 2650 47500 2710 47510
rect 2850 47500 2860 47520
rect 2920 47500 2930 47560
rect 2850 47490 2930 47500
rect 3690 47500 3700 47560
rect 3760 47550 3770 47560
rect 3760 47520 4070 47550
rect 3760 47500 3770 47520
rect 4070 47500 4130 47510
rect 7640 47570 7700 47580
rect 8260 47570 8270 47630
rect 8330 47610 8910 47630
rect 8330 47570 8340 47610
rect 13900 47660 13960 47670
rect 8910 47590 8970 47600
rect 13250 47630 13900 47640
rect 9060 47570 9120 47580
rect 7840 47560 7920 47570
rect 8260 47560 8340 47570
rect 8680 47560 8760 47570
rect 7840 47550 7850 47560
rect 7700 47520 7850 47550
rect 7640 47500 7700 47510
rect 7840 47500 7850 47520
rect 7910 47500 7920 47560
rect 3690 47490 3770 47500
rect 7840 47490 7920 47500
rect 8680 47500 8690 47560
rect 8750 47550 8760 47560
rect 8750 47520 9060 47550
rect 8750 47500 8760 47520
rect 9060 47500 9120 47510
rect 12510 47570 12570 47580
rect 13250 47570 13260 47630
rect 13320 47610 13900 47630
rect 13320 47570 13330 47610
rect 18890 47660 18950 47670
rect 13900 47590 13960 47600
rect 18240 47630 18890 47640
rect 14170 47570 14230 47580
rect 12830 47560 12910 47570
rect 13250 47560 13330 47570
rect 13670 47560 13750 47570
rect 12830 47550 12840 47560
rect 12570 47520 12840 47550
rect 12510 47500 12570 47510
rect 12830 47500 12840 47520
rect 12900 47500 12910 47560
rect 8680 47490 8760 47500
rect 12830 47490 12910 47500
rect 13670 47500 13680 47560
rect 13740 47550 13750 47560
rect 13740 47520 14170 47550
rect 13740 47500 13750 47520
rect 14170 47500 14230 47510
rect 17500 47570 17560 47580
rect 18240 47570 18250 47630
rect 18310 47610 18890 47630
rect 18310 47570 18320 47610
rect 18890 47590 18950 47600
rect 19160 47570 19220 47580
rect 17820 47560 17900 47570
rect 18240 47560 18320 47570
rect 18660 47560 18740 47570
rect 17820 47550 17830 47560
rect 17560 47520 17830 47550
rect 17500 47500 17560 47510
rect 17820 47500 17830 47520
rect 17890 47500 17900 47560
rect 13670 47490 13750 47500
rect 17820 47490 17900 47500
rect 18660 47500 18670 47560
rect 18730 47550 18740 47560
rect 18730 47520 19160 47550
rect 18730 47500 18740 47520
rect 19160 47500 19220 47510
rect 18660 47490 18740 47500
rect 3260 47470 3360 47480
rect 3260 47400 3280 47470
rect 3350 47400 3360 47470
rect 3260 47360 3360 47400
rect 3260 47290 3280 47360
rect 3350 47290 3360 47360
rect 3260 47270 3360 47290
rect 8250 47470 8350 47480
rect 8250 47400 8270 47470
rect 8340 47400 8350 47470
rect 8250 47360 8350 47400
rect 8250 47290 8270 47360
rect 8340 47290 8350 47360
rect 8250 47270 8350 47290
rect 13240 47470 13340 47480
rect 13240 47400 13260 47470
rect 13330 47400 13340 47470
rect 13240 47360 13340 47400
rect 13240 47290 13260 47360
rect 13330 47290 13340 47360
rect 13240 47270 13340 47290
rect 18230 47470 18330 47480
rect 18230 47400 18250 47470
rect 18320 47400 18330 47470
rect 18230 47360 18330 47400
rect 18230 47290 18250 47360
rect 18320 47290 18330 47360
rect 18230 47270 18330 47290
rect 2630 47250 2710 47260
rect 2630 47190 2640 47250
rect 2700 47240 2710 47250
rect 2850 47250 2930 47260
rect 2850 47240 2860 47250
rect 2700 47210 2860 47240
rect 2700 47190 2710 47210
rect 2630 47180 2710 47190
rect 2850 47190 2860 47210
rect 2920 47190 2930 47250
rect 3690 47250 3770 47260
rect 3690 47190 3700 47250
rect 3760 47240 3770 47250
rect 4070 47250 4150 47260
rect 4070 47240 4080 47250
rect 3760 47210 4080 47240
rect 3760 47190 3770 47210
rect 2850 47180 2930 47190
rect 3270 47180 3350 47190
rect 3690 47180 3770 47190
rect 4070 47190 4080 47210
rect 4140 47190 4150 47250
rect 4070 47180 4150 47190
rect 7620 47250 7700 47260
rect 7620 47190 7630 47250
rect 7690 47240 7700 47250
rect 7840 47250 7920 47260
rect 7840 47240 7850 47250
rect 7690 47210 7850 47240
rect 7690 47190 7700 47210
rect 7620 47180 7700 47190
rect 7840 47190 7850 47210
rect 7910 47190 7920 47250
rect 8680 47250 8760 47260
rect 8680 47190 8690 47250
rect 8750 47240 8760 47250
rect 9060 47250 9140 47260
rect 9060 47240 9070 47250
rect 8750 47210 9070 47240
rect 8750 47190 8760 47210
rect 7840 47180 7920 47190
rect 8260 47180 8340 47190
rect 8680 47180 8760 47190
rect 9060 47190 9070 47210
rect 9130 47190 9140 47250
rect 9060 47180 9140 47190
rect 12490 47250 12570 47260
rect 12490 47190 12500 47250
rect 12560 47240 12570 47250
rect 12830 47250 12910 47260
rect 12830 47240 12840 47250
rect 12560 47210 12840 47240
rect 12560 47190 12570 47210
rect 12490 47180 12570 47190
rect 12830 47190 12840 47210
rect 12900 47190 12910 47250
rect 13670 47250 13750 47260
rect 13670 47190 13680 47250
rect 13740 47240 13750 47250
rect 14170 47250 14250 47260
rect 14170 47240 14180 47250
rect 13740 47210 14180 47240
rect 13740 47190 13750 47210
rect 12830 47180 12910 47190
rect 13250 47180 13330 47190
rect 13670 47180 13750 47190
rect 14170 47190 14180 47210
rect 14240 47190 14250 47250
rect 14170 47180 14250 47190
rect 17480 47250 17560 47260
rect 17480 47190 17490 47250
rect 17550 47240 17560 47250
rect 17820 47250 17900 47260
rect 17820 47240 17830 47250
rect 17550 47210 17830 47240
rect 17550 47190 17560 47210
rect 17480 47180 17560 47190
rect 17820 47190 17830 47210
rect 17890 47190 17900 47250
rect 18660 47250 18740 47260
rect 18660 47190 18670 47250
rect 18730 47240 18740 47250
rect 19160 47250 19240 47260
rect 19160 47240 19170 47250
rect 18730 47210 19170 47240
rect 18730 47190 18740 47210
rect 17820 47180 17900 47190
rect 18240 47180 18320 47190
rect 18660 47180 18740 47190
rect 19160 47190 19170 47210
rect 19230 47190 19240 47250
rect 19160 47180 19240 47190
rect 3270 47120 3280 47180
rect 3340 47140 3350 47180
rect 3340 47130 4040 47140
rect 3340 47120 3980 47130
rect 3270 47110 3980 47120
rect 8260 47120 8270 47180
rect 8330 47140 8340 47180
rect 8330 47130 9030 47140
rect 8330 47120 8970 47130
rect 8260 47110 8970 47120
rect 3980 47060 4040 47070
rect 8970 47060 9030 47070
rect 3920 45950 3980 45960
rect 3270 45920 3920 45930
rect 2650 45860 2710 45870
rect 3270 45860 3280 45920
rect 3340 45900 3920 45920
rect 3340 45860 3350 45900
rect 8910 45950 8970 45960
rect 3920 45880 3980 45890
rect 8260 45920 8910 45930
rect 4070 45860 4130 45870
rect 2850 45850 2930 45860
rect 3270 45850 3350 45860
rect 3690 45850 3770 45860
rect 2850 45840 2860 45850
rect 2710 45810 2860 45840
rect 2650 45790 2710 45800
rect 2850 45790 2860 45810
rect 2920 45790 2930 45850
rect 2850 45780 2930 45790
rect 3690 45790 3700 45850
rect 3760 45840 3770 45850
rect 3760 45810 4070 45840
rect 3760 45790 3770 45810
rect 4070 45790 4130 45800
rect 7640 45860 7700 45870
rect 8260 45860 8270 45920
rect 8330 45900 8910 45920
rect 8330 45860 8340 45900
rect 8910 45880 8970 45890
rect 9060 45860 9120 45870
rect 7840 45850 7920 45860
rect 8260 45850 8340 45860
rect 8680 45850 8760 45860
rect 7840 45840 7850 45850
rect 7700 45810 7850 45840
rect 7640 45790 7700 45800
rect 7840 45790 7850 45810
rect 7910 45790 7920 45850
rect 3690 45780 3770 45790
rect 7840 45780 7920 45790
rect 8680 45790 8690 45850
rect 8750 45840 8760 45850
rect 8750 45810 9060 45840
rect 8750 45790 8760 45810
rect 9060 45790 9120 45800
rect 8680 45780 8760 45790
rect 3260 45760 3360 45770
rect 3260 45690 3280 45760
rect 3350 45690 3360 45760
rect 3260 45650 3360 45690
rect 3260 45580 3280 45650
rect 3350 45580 3360 45650
rect 3260 45560 3360 45580
rect 8250 45760 8350 45770
rect 8250 45690 8270 45760
rect 8340 45690 8350 45760
rect 8250 45650 8350 45690
rect 8250 45580 8270 45650
rect 8340 45580 8350 45650
rect 8250 45560 8350 45580
rect 2630 45540 2710 45550
rect 2630 45480 2640 45540
rect 2700 45530 2710 45540
rect 2850 45540 2930 45550
rect 2850 45530 2860 45540
rect 2700 45500 2860 45530
rect 2700 45480 2710 45500
rect 2630 45470 2710 45480
rect 2850 45480 2860 45500
rect 2920 45480 2930 45540
rect 3690 45540 3770 45550
rect 3690 45480 3700 45540
rect 3760 45530 3770 45540
rect 4070 45540 4150 45550
rect 4070 45530 4080 45540
rect 3760 45500 4080 45530
rect 3760 45480 3770 45500
rect 2850 45470 2930 45480
rect 3270 45470 3350 45480
rect 3690 45470 3770 45480
rect 4070 45480 4080 45500
rect 4140 45480 4150 45540
rect 4070 45470 4150 45480
rect 7620 45540 7700 45550
rect 7620 45480 7630 45540
rect 7690 45530 7700 45540
rect 7840 45540 7920 45550
rect 7840 45530 7850 45540
rect 7690 45500 7850 45530
rect 7690 45480 7700 45500
rect 7620 45470 7700 45480
rect 7840 45480 7850 45500
rect 7910 45480 7920 45540
rect 8680 45540 8760 45550
rect 8680 45480 8690 45540
rect 8750 45530 8760 45540
rect 9060 45540 9140 45550
rect 9060 45530 9070 45540
rect 8750 45500 9070 45530
rect 8750 45480 8760 45500
rect 7840 45470 7920 45480
rect 8260 45470 8340 45480
rect 8680 45470 8760 45480
rect 9060 45480 9070 45500
rect 9130 45480 9140 45540
rect 9060 45470 9140 45480
rect 3270 45410 3280 45470
rect 3340 45430 3350 45470
rect 3340 45420 4040 45430
rect 3340 45410 3980 45420
rect 3270 45400 3980 45410
rect 8260 45410 8270 45470
rect 8330 45430 8340 45470
rect 8330 45420 9030 45430
rect 8330 45410 8970 45420
rect 8260 45400 8970 45410
rect 3980 45350 4040 45360
rect 8970 45350 9030 45360
rect 3920 44240 3980 44250
rect 3270 44210 3920 44220
rect 2650 44150 2710 44160
rect 3270 44150 3280 44210
rect 3340 44190 3920 44210
rect 3340 44150 3350 44190
rect 8910 44240 8970 44250
rect 3920 44170 3980 44180
rect 8260 44210 8910 44220
rect 4070 44150 4130 44160
rect 2850 44140 2930 44150
rect 3270 44140 3350 44150
rect 3690 44140 3770 44150
rect 2850 44130 2860 44140
rect 2710 44100 2860 44130
rect 2650 44080 2710 44090
rect 2850 44080 2860 44100
rect 2920 44080 2930 44140
rect 2850 44070 2930 44080
rect 3690 44080 3700 44140
rect 3760 44130 3770 44140
rect 3760 44100 4070 44130
rect 3760 44080 3770 44100
rect 4070 44080 4130 44090
rect 7640 44150 7700 44160
rect 8260 44150 8270 44210
rect 8330 44190 8910 44210
rect 8330 44150 8340 44190
rect 8910 44170 8970 44180
rect 9060 44150 9120 44160
rect 7840 44140 7920 44150
rect 8260 44140 8340 44150
rect 8680 44140 8760 44150
rect 7840 44130 7850 44140
rect 7700 44100 7850 44130
rect 7640 44080 7700 44090
rect 7840 44080 7850 44100
rect 7910 44080 7920 44140
rect 3690 44070 3770 44080
rect 7840 44070 7920 44080
rect 8680 44080 8690 44140
rect 8750 44130 8760 44140
rect 8750 44100 9060 44130
rect 8750 44080 8760 44100
rect 9060 44080 9120 44090
rect 8680 44070 8760 44080
rect 3260 44050 3360 44060
rect 3260 43980 3280 44050
rect 3350 43980 3360 44050
rect 3260 43940 3360 43980
rect 3260 43870 3280 43940
rect 3350 43870 3360 43940
rect 3260 43850 3360 43870
rect 8250 44050 8350 44060
rect 8250 43980 8270 44050
rect 8340 43980 8350 44050
rect 8250 43940 8350 43980
rect 8250 43870 8270 43940
rect 8340 43870 8350 43940
rect 8250 43850 8350 43870
rect 2630 43830 2710 43840
rect 2630 43770 2640 43830
rect 2700 43820 2710 43830
rect 2850 43830 2930 43840
rect 2850 43820 2860 43830
rect 2700 43790 2860 43820
rect 2700 43770 2710 43790
rect 2630 43760 2710 43770
rect 2850 43770 2860 43790
rect 2920 43770 2930 43830
rect 3690 43830 3770 43840
rect 3690 43770 3700 43830
rect 3760 43820 3770 43830
rect 4070 43830 4150 43840
rect 4070 43820 4080 43830
rect 3760 43790 4080 43820
rect 3760 43770 3770 43790
rect 2850 43760 2930 43770
rect 3270 43760 3350 43770
rect 3690 43760 3770 43770
rect 4070 43770 4080 43790
rect 4140 43770 4150 43830
rect 4070 43760 4150 43770
rect 7620 43830 7700 43840
rect 7620 43770 7630 43830
rect 7690 43820 7700 43830
rect 7840 43830 7920 43840
rect 7840 43820 7850 43830
rect 7690 43790 7850 43820
rect 7690 43770 7700 43790
rect 7620 43760 7700 43770
rect 7840 43770 7850 43790
rect 7910 43770 7920 43830
rect 8680 43830 8760 43840
rect 8680 43770 8690 43830
rect 8750 43820 8760 43830
rect 9060 43830 9140 43840
rect 9060 43820 9070 43830
rect 8750 43790 9070 43820
rect 8750 43770 8760 43790
rect 7840 43760 7920 43770
rect 8260 43760 8340 43770
rect 8680 43760 8760 43770
rect 9060 43770 9070 43790
rect 9130 43770 9140 43830
rect 9060 43760 9140 43770
rect 3270 43700 3280 43760
rect 3340 43720 3350 43760
rect 3340 43710 4040 43720
rect 3340 43700 3980 43710
rect 3270 43690 3980 43700
rect 8260 43700 8270 43760
rect 8330 43720 8340 43760
rect 8330 43710 9030 43720
rect 8330 43700 8970 43710
rect 8260 43690 8970 43700
rect 3980 43640 4040 43650
rect 8970 43640 9030 43650
rect 3920 42530 3980 42540
rect 3270 42500 3920 42510
rect 2650 42440 2710 42450
rect 3270 42440 3280 42500
rect 3340 42480 3920 42500
rect 3340 42440 3350 42480
rect 8910 42530 8970 42540
rect 3920 42460 3980 42470
rect 8260 42500 8910 42510
rect 4070 42440 4130 42450
rect 2850 42430 2930 42440
rect 3270 42430 3350 42440
rect 3690 42430 3770 42440
rect 2850 42420 2860 42430
rect 2710 42390 2860 42420
rect 2650 42370 2710 42380
rect 2850 42370 2860 42390
rect 2920 42370 2930 42430
rect 2850 42360 2930 42370
rect 3690 42370 3700 42430
rect 3760 42420 3770 42430
rect 3760 42390 4070 42420
rect 3760 42370 3770 42390
rect 4070 42370 4130 42380
rect 7640 42440 7700 42450
rect 8260 42440 8270 42500
rect 8330 42480 8910 42500
rect 8330 42440 8340 42480
rect 8910 42460 8970 42470
rect 9060 42440 9120 42450
rect 7840 42430 7920 42440
rect 8260 42430 8340 42440
rect 8680 42430 8760 42440
rect 7840 42420 7850 42430
rect 7700 42390 7850 42420
rect 7640 42370 7700 42380
rect 7840 42370 7850 42390
rect 7910 42370 7920 42430
rect 3690 42360 3770 42370
rect 7840 42360 7920 42370
rect 8680 42370 8690 42430
rect 8750 42420 8760 42430
rect 8750 42390 9060 42420
rect 8750 42370 8760 42390
rect 9060 42370 9120 42380
rect 8680 42360 8760 42370
rect 3260 42340 3360 42350
rect 3260 42270 3280 42340
rect 3350 42270 3360 42340
rect 3260 42230 3360 42270
rect 3260 42160 3280 42230
rect 3350 42160 3360 42230
rect 3260 42140 3360 42160
rect 8250 42340 8350 42350
rect 8250 42270 8270 42340
rect 8340 42270 8350 42340
rect 8250 42230 8350 42270
rect 8250 42160 8270 42230
rect 8340 42160 8350 42230
rect 8250 42140 8350 42160
rect 2630 42120 2710 42130
rect 2630 42060 2640 42120
rect 2700 42110 2710 42120
rect 2850 42120 2930 42130
rect 2850 42110 2860 42120
rect 2700 42080 2860 42110
rect 2700 42060 2710 42080
rect 2630 42050 2710 42060
rect 2850 42060 2860 42080
rect 2920 42060 2930 42120
rect 3690 42120 3770 42130
rect 3690 42060 3700 42120
rect 3760 42110 3770 42120
rect 4070 42120 4150 42130
rect 4070 42110 4080 42120
rect 3760 42080 4080 42110
rect 3760 42060 3770 42080
rect 2850 42050 2930 42060
rect 3270 42050 3350 42060
rect 3690 42050 3770 42060
rect 4070 42060 4080 42080
rect 4140 42060 4150 42120
rect 4070 42050 4150 42060
rect 7620 42120 7700 42130
rect 7620 42060 7630 42120
rect 7690 42110 7700 42120
rect 7840 42120 7920 42130
rect 7840 42110 7850 42120
rect 7690 42080 7850 42110
rect 7690 42060 7700 42080
rect 7620 42050 7700 42060
rect 7840 42060 7850 42080
rect 7910 42060 7920 42120
rect 8680 42120 8760 42130
rect 8680 42060 8690 42120
rect 8750 42110 8760 42120
rect 9060 42120 9140 42130
rect 9060 42110 9070 42120
rect 8750 42080 9070 42110
rect 8750 42060 8760 42080
rect 7840 42050 7920 42060
rect 8260 42050 8340 42060
rect 8680 42050 8760 42060
rect 9060 42060 9070 42080
rect 9130 42060 9140 42120
rect 9060 42050 9140 42060
rect 3270 41990 3280 42050
rect 3340 42010 3350 42050
rect 3340 42000 4040 42010
rect 3340 41990 3980 42000
rect 3270 41980 3980 41990
rect 8260 41990 8270 42050
rect 8330 42010 8340 42050
rect 8330 42000 9030 42010
rect 8330 41990 8970 42000
rect 8260 41980 8970 41990
rect 3980 41930 4040 41940
rect 8970 41930 9030 41940
rect 3920 40820 3980 40830
rect 3270 40790 3920 40800
rect 2650 40730 2710 40740
rect 3270 40730 3280 40790
rect 3340 40770 3920 40790
rect 3340 40730 3350 40770
rect 8910 40820 8970 40830
rect 3920 40750 3980 40760
rect 8260 40790 8910 40800
rect 4070 40730 4130 40740
rect 2850 40720 2930 40730
rect 3270 40720 3350 40730
rect 3690 40720 3770 40730
rect 2850 40710 2860 40720
rect 2710 40680 2860 40710
rect 2650 40660 2710 40670
rect 2850 40660 2860 40680
rect 2920 40660 2930 40720
rect 2850 40650 2930 40660
rect 3690 40660 3700 40720
rect 3760 40710 3770 40720
rect 3760 40680 4070 40710
rect 3760 40660 3770 40680
rect 4070 40660 4130 40670
rect 7640 40730 7700 40740
rect 8260 40730 8270 40790
rect 8330 40770 8910 40790
rect 8330 40730 8340 40770
rect 8910 40750 8970 40760
rect 9060 40730 9120 40740
rect 7840 40720 7920 40730
rect 8260 40720 8340 40730
rect 8680 40720 8760 40730
rect 7840 40710 7850 40720
rect 7700 40680 7850 40710
rect 7640 40660 7700 40670
rect 7840 40660 7850 40680
rect 7910 40660 7920 40720
rect 3690 40650 3770 40660
rect 7840 40650 7920 40660
rect 8680 40660 8690 40720
rect 8750 40710 8760 40720
rect 8750 40680 9060 40710
rect 8750 40660 8760 40680
rect 9060 40660 9120 40670
rect 8680 40650 8760 40660
rect 3260 40630 3360 40640
rect 3260 40560 3280 40630
rect 3350 40560 3360 40630
rect 3260 40520 3360 40560
rect 3260 40450 3280 40520
rect 3350 40450 3360 40520
rect 3260 40430 3360 40450
rect 8250 40630 8350 40640
rect 8250 40560 8270 40630
rect 8340 40560 8350 40630
rect 8250 40520 8350 40560
rect 8250 40450 8270 40520
rect 8340 40450 8350 40520
rect 8250 40430 8350 40450
rect 2630 40410 2710 40420
rect 2630 40350 2640 40410
rect 2700 40400 2710 40410
rect 2850 40410 2930 40420
rect 2850 40400 2860 40410
rect 2700 40370 2860 40400
rect 2700 40350 2710 40370
rect 2630 40340 2710 40350
rect 2850 40350 2860 40370
rect 2920 40350 2930 40410
rect 3690 40410 3770 40420
rect 3690 40350 3700 40410
rect 3760 40400 3770 40410
rect 4070 40410 4150 40420
rect 4070 40400 4080 40410
rect 3760 40370 4080 40400
rect 3760 40350 3770 40370
rect 2850 40340 2930 40350
rect 3270 40340 3350 40350
rect 3690 40340 3770 40350
rect 4070 40350 4080 40370
rect 4140 40350 4150 40410
rect 4070 40340 4150 40350
rect 7620 40410 7700 40420
rect 7620 40350 7630 40410
rect 7690 40400 7700 40410
rect 7840 40410 7920 40420
rect 7840 40400 7850 40410
rect 7690 40370 7850 40400
rect 7690 40350 7700 40370
rect 7620 40340 7700 40350
rect 7840 40350 7850 40370
rect 7910 40350 7920 40410
rect 8680 40410 8760 40420
rect 8680 40350 8690 40410
rect 8750 40400 8760 40410
rect 9060 40410 9140 40420
rect 9060 40400 9070 40410
rect 8750 40370 9070 40400
rect 8750 40350 8760 40370
rect 7840 40340 7920 40350
rect 8260 40340 8340 40350
rect 8680 40340 8760 40350
rect 9060 40350 9070 40370
rect 9130 40350 9140 40410
rect 9060 40340 9140 40350
rect 2680 39240 2710 40340
rect 3270 40280 3280 40340
rect 3340 40300 3350 40340
rect 3340 40290 4040 40300
rect 3340 40280 3980 40290
rect 3270 40270 3980 40280
rect 3980 40220 4040 40230
rect 2450 39230 2510 39240
rect 2450 39160 2510 39170
rect 2540 39210 2710 39240
rect 2740 39680 2820 39690
rect 2740 39620 2750 39680
rect 2810 39620 2820 39680
rect 3810 39680 3890 39690
rect 3810 39620 3820 39680
rect 3880 39620 3890 39680
rect 2450 36180 2480 39160
rect 2540 36320 2570 39210
rect 2740 38840 2810 39620
rect 3810 39610 3890 39620
rect 3980 39680 4040 39690
rect 3980 39610 4040 39620
rect 2740 38830 2820 38840
rect 2740 38770 2750 38830
rect 2810 38770 2820 38830
rect 2740 38760 2820 38770
rect 3820 38700 3890 39610
rect 4010 38700 4040 39610
rect 4070 39240 4100 40340
rect 7670 39240 7700 40340
rect 8260 40280 8270 40340
rect 8330 40300 8340 40340
rect 8330 40290 9030 40300
rect 8330 40280 8970 40290
rect 8260 40270 8970 40280
rect 8970 40220 9030 40230
rect 4070 39210 4240 39240
rect 3810 38690 3890 38700
rect 3810 38630 3820 38690
rect 3880 38630 3890 38690
rect 3960 38640 3970 38700
rect 4030 38640 4040 38700
rect 3810 38620 3890 38630
rect 4210 36320 4240 39210
rect 4270 39230 4330 39240
rect 4270 39160 4330 39170
rect 2510 36310 2590 36320
rect 2510 36250 2520 36310
rect 2580 36250 2590 36310
rect 4190 36260 4200 36320
rect 4260 36260 4270 36320
rect 2510 36240 2590 36250
rect 4300 36180 4330 39160
rect 2450 36170 2530 36180
rect 2450 36110 2460 36170
rect 2520 36110 2530 36170
rect 4250 36120 4260 36180
rect 4320 36120 4330 36180
rect 7440 39230 7500 39240
rect 7440 39160 7500 39170
rect 7530 39210 7700 39240
rect 7730 39680 7810 39690
rect 7730 39620 7740 39680
rect 7800 39620 7810 39680
rect 8800 39680 8880 39690
rect 8800 39620 8810 39680
rect 8870 39620 8880 39680
rect 7440 36180 7470 39160
rect 7530 36320 7560 39210
rect 7730 38840 7800 39620
rect 8800 39610 8880 39620
rect 8970 39680 9030 39690
rect 8970 39610 9030 39620
rect 7730 38830 7810 38840
rect 7730 38770 7740 38830
rect 7800 38770 7810 38830
rect 7730 38760 7810 38770
rect 8810 38700 8880 39610
rect 9000 38700 9030 39610
rect 9060 39240 9090 40340
rect 12540 39300 12570 47180
rect 13250 47120 13260 47180
rect 13320 47140 13330 47180
rect 13320 47130 14020 47140
rect 13320 47120 13960 47130
rect 13250 47110 13960 47120
rect 13960 47060 14020 47070
rect 13900 45950 13960 45960
rect 13250 45920 13900 45930
rect 12630 45860 12690 45870
rect 13250 45860 13260 45920
rect 13320 45900 13900 45920
rect 13320 45860 13330 45900
rect 13900 45880 13960 45890
rect 14050 45860 14110 45870
rect 12830 45850 12910 45860
rect 13250 45850 13330 45860
rect 13670 45850 13750 45860
rect 12830 45840 12840 45850
rect 12690 45810 12840 45840
rect 12630 45790 12690 45800
rect 12830 45790 12840 45810
rect 12900 45790 12910 45850
rect 12830 45780 12910 45790
rect 13670 45790 13680 45850
rect 13740 45840 13750 45850
rect 13740 45810 14050 45840
rect 13740 45790 13750 45810
rect 14050 45790 14110 45800
rect 13670 45780 13750 45790
rect 13240 45760 13340 45770
rect 13240 45690 13260 45760
rect 13330 45690 13340 45760
rect 13240 45650 13340 45690
rect 13240 45580 13260 45650
rect 13330 45580 13340 45650
rect 13240 45560 13340 45580
rect 12610 45540 12690 45550
rect 12610 45480 12620 45540
rect 12680 45530 12690 45540
rect 12830 45540 12910 45550
rect 12830 45530 12840 45540
rect 12680 45500 12840 45530
rect 12680 45480 12690 45500
rect 12610 45470 12690 45480
rect 12830 45480 12840 45500
rect 12900 45480 12910 45540
rect 13670 45540 13750 45550
rect 13670 45480 13680 45540
rect 13740 45530 13750 45540
rect 14050 45540 14130 45550
rect 14050 45530 14060 45540
rect 13740 45500 14060 45530
rect 13740 45480 13750 45500
rect 12830 45470 12910 45480
rect 13250 45470 13330 45480
rect 13670 45470 13750 45480
rect 14050 45480 14060 45500
rect 14120 45480 14130 45540
rect 14050 45470 14130 45480
rect 13250 45410 13260 45470
rect 13320 45430 13330 45470
rect 13320 45420 14020 45430
rect 13320 45410 13960 45420
rect 13250 45400 13960 45410
rect 13960 45350 14020 45360
rect 13900 44240 13960 44250
rect 13250 44210 13900 44220
rect 12630 44150 12690 44160
rect 13250 44150 13260 44210
rect 13320 44190 13900 44210
rect 13320 44150 13330 44190
rect 13900 44170 13960 44180
rect 14050 44150 14110 44160
rect 12830 44140 12910 44150
rect 13250 44140 13330 44150
rect 13670 44140 13750 44150
rect 12830 44130 12840 44140
rect 12690 44100 12840 44130
rect 12630 44080 12690 44090
rect 12830 44080 12840 44100
rect 12900 44080 12910 44140
rect 12830 44070 12910 44080
rect 13670 44080 13680 44140
rect 13740 44130 13750 44140
rect 13740 44100 14050 44130
rect 13740 44080 13750 44100
rect 14050 44080 14110 44090
rect 13670 44070 13750 44080
rect 13240 44050 13340 44060
rect 13240 43980 13260 44050
rect 13330 43980 13340 44050
rect 13240 43940 13340 43980
rect 13240 43870 13260 43940
rect 13330 43870 13340 43940
rect 13240 43850 13340 43870
rect 12610 43830 12690 43840
rect 12610 43770 12620 43830
rect 12680 43820 12690 43830
rect 12830 43830 12910 43840
rect 12830 43820 12840 43830
rect 12680 43790 12840 43820
rect 12680 43770 12690 43790
rect 12610 43760 12690 43770
rect 12830 43770 12840 43790
rect 12900 43770 12910 43830
rect 13670 43830 13750 43840
rect 13670 43770 13680 43830
rect 13740 43820 13750 43830
rect 14050 43830 14130 43840
rect 14050 43820 14060 43830
rect 13740 43790 14060 43820
rect 13740 43770 13750 43790
rect 12830 43760 12910 43770
rect 13250 43760 13330 43770
rect 13670 43760 13750 43770
rect 14050 43770 14060 43790
rect 14120 43770 14130 43830
rect 14050 43760 14130 43770
rect 13250 43700 13260 43760
rect 13320 43720 13330 43760
rect 13320 43710 14020 43720
rect 13320 43700 13960 43710
rect 13250 43690 13960 43700
rect 13960 43640 14020 43650
rect 13900 42530 13960 42540
rect 13250 42500 13900 42510
rect 12630 42440 12690 42450
rect 13250 42440 13260 42500
rect 13320 42480 13900 42500
rect 13320 42440 13330 42480
rect 13900 42460 13960 42470
rect 14050 42440 14110 42450
rect 12830 42430 12910 42440
rect 13250 42430 13330 42440
rect 13670 42430 13750 42440
rect 12830 42420 12840 42430
rect 12690 42390 12840 42420
rect 12630 42370 12690 42380
rect 12830 42370 12840 42390
rect 12900 42370 12910 42430
rect 12830 42360 12910 42370
rect 13670 42370 13680 42430
rect 13740 42420 13750 42430
rect 13740 42390 14050 42420
rect 13740 42370 13750 42390
rect 14050 42370 14110 42380
rect 13670 42360 13750 42370
rect 13240 42340 13340 42350
rect 13240 42270 13260 42340
rect 13330 42270 13340 42340
rect 13240 42230 13340 42270
rect 13240 42160 13260 42230
rect 13330 42160 13340 42230
rect 13240 42140 13340 42160
rect 12610 42120 12690 42130
rect 12610 42060 12620 42120
rect 12680 42110 12690 42120
rect 12830 42120 12910 42130
rect 12830 42110 12840 42120
rect 12680 42080 12840 42110
rect 12680 42060 12690 42080
rect 12610 42050 12690 42060
rect 12830 42060 12840 42080
rect 12900 42060 12910 42120
rect 13670 42120 13750 42130
rect 13670 42060 13680 42120
rect 13740 42110 13750 42120
rect 14050 42120 14130 42130
rect 14050 42110 14060 42120
rect 13740 42080 14060 42110
rect 13740 42060 13750 42080
rect 12830 42050 12910 42060
rect 13250 42050 13330 42060
rect 13670 42050 13750 42060
rect 14050 42060 14060 42080
rect 14120 42060 14130 42120
rect 14050 42050 14130 42060
rect 13250 41990 13260 42050
rect 13320 42010 13330 42050
rect 13320 42000 14020 42010
rect 13320 41990 13960 42000
rect 13250 41980 13960 41990
rect 13960 41930 14020 41940
rect 13900 40820 13960 40830
rect 13250 40790 13900 40800
rect 12630 40730 12690 40740
rect 13250 40730 13260 40790
rect 13320 40770 13900 40790
rect 13320 40730 13330 40770
rect 13900 40750 13960 40760
rect 14050 40730 14110 40740
rect 12830 40720 12910 40730
rect 13250 40720 13330 40730
rect 13670 40720 13750 40730
rect 12830 40710 12840 40720
rect 12690 40680 12840 40710
rect 12630 40660 12690 40670
rect 12830 40660 12840 40680
rect 12900 40660 12910 40720
rect 12830 40650 12910 40660
rect 13670 40660 13680 40720
rect 13740 40710 13750 40720
rect 13740 40680 14050 40710
rect 13740 40660 13750 40680
rect 14050 40660 14110 40670
rect 13670 40650 13750 40660
rect 13240 40630 13340 40640
rect 13240 40560 13260 40630
rect 13330 40560 13340 40630
rect 13240 40520 13340 40560
rect 13240 40450 13260 40520
rect 13330 40450 13340 40520
rect 13240 40430 13340 40450
rect 12610 40410 12690 40420
rect 12610 40350 12620 40410
rect 12680 40400 12690 40410
rect 12830 40410 12910 40420
rect 12830 40400 12840 40410
rect 12680 40370 12840 40400
rect 12680 40350 12690 40370
rect 12610 40340 12690 40350
rect 12830 40350 12840 40370
rect 12900 40350 12910 40410
rect 13670 40410 13750 40420
rect 13670 40350 13680 40410
rect 13740 40400 13750 40410
rect 14050 40410 14130 40420
rect 14050 40400 14060 40410
rect 13740 40370 14060 40400
rect 13740 40350 13750 40370
rect 12830 40340 12910 40350
rect 13250 40340 13330 40350
rect 13670 40340 13750 40350
rect 14050 40350 14060 40370
rect 14120 40350 14130 40410
rect 14050 40340 14130 40350
rect 12250 39290 12310 39300
rect 9060 39210 9230 39240
rect 8800 38690 8880 38700
rect 8800 38630 8810 38690
rect 8870 38630 8880 38690
rect 8950 38640 8960 38700
rect 9020 38640 9030 38700
rect 8800 38620 8880 38630
rect 9200 36320 9230 39210
rect 9260 39230 9320 39240
rect 9260 39160 9320 39170
rect 7500 36310 7580 36320
rect 7500 36250 7510 36310
rect 7570 36250 7580 36310
rect 9180 36260 9190 36320
rect 9250 36260 9260 36320
rect 7500 36240 7580 36250
rect 9290 36180 9320 39160
rect 12250 39220 12310 39230
rect 12340 39270 12570 39300
rect 12250 36460 12280 39220
rect 12340 36600 12370 39270
rect 12660 39240 12690 40340
rect 13250 40280 13260 40340
rect 13320 40300 13330 40340
rect 13320 40290 14020 40300
rect 13320 40280 13960 40290
rect 13250 40270 13960 40280
rect 13960 40220 14020 40230
rect 12430 39230 12490 39240
rect 12430 39160 12490 39170
rect 12520 39210 12690 39240
rect 12720 39680 12800 39690
rect 12720 39620 12730 39680
rect 12790 39620 12800 39680
rect 13790 39680 13870 39690
rect 13790 39620 13800 39680
rect 13860 39620 13870 39680
rect 12310 36590 12390 36600
rect 12310 36530 12320 36590
rect 12380 36530 12390 36590
rect 12310 36520 12390 36530
rect 12250 36450 12330 36460
rect 12250 36390 12260 36450
rect 12320 36390 12330 36450
rect 12250 36380 12330 36390
rect 7440 36170 7520 36180
rect 2450 36100 2530 36110
rect 7440 36110 7450 36170
rect 7510 36110 7520 36170
rect 9240 36120 9250 36180
rect 9310 36120 9320 36180
rect 12430 36180 12460 39160
rect 12520 36320 12550 39210
rect 12720 38840 12790 39620
rect 13790 39610 13870 39620
rect 13960 39680 14020 39690
rect 13960 39610 14020 39620
rect 12720 38830 12800 38840
rect 12720 38770 12730 38830
rect 12790 38770 12800 38830
rect 12720 38760 12800 38770
rect 13800 38700 13870 39610
rect 13990 38700 14020 39610
rect 14050 39240 14080 40340
rect 14170 39300 14200 47180
rect 17530 39300 17560 47180
rect 18240 47120 18250 47180
rect 18310 47140 18320 47180
rect 18310 47130 19010 47140
rect 18310 47120 18950 47130
rect 18240 47110 18950 47120
rect 18950 47060 19010 47070
rect 18890 45950 18950 45960
rect 18240 45920 18890 45930
rect 17620 45860 17680 45870
rect 18240 45860 18250 45920
rect 18310 45900 18890 45920
rect 18310 45860 18320 45900
rect 18890 45880 18950 45890
rect 19040 45860 19100 45870
rect 17820 45850 17900 45860
rect 18240 45850 18320 45860
rect 18660 45850 18740 45860
rect 17820 45840 17830 45850
rect 17680 45810 17830 45840
rect 17620 45790 17680 45800
rect 17820 45790 17830 45810
rect 17890 45790 17900 45850
rect 17820 45780 17900 45790
rect 18660 45790 18670 45850
rect 18730 45840 18740 45850
rect 18730 45810 19040 45840
rect 18730 45790 18740 45810
rect 19040 45790 19100 45800
rect 18660 45780 18740 45790
rect 18230 45760 18330 45770
rect 18230 45690 18250 45760
rect 18320 45690 18330 45760
rect 18230 45650 18330 45690
rect 18230 45580 18250 45650
rect 18320 45580 18330 45650
rect 18230 45560 18330 45580
rect 17600 45540 17680 45550
rect 17600 45480 17610 45540
rect 17670 45530 17680 45540
rect 17820 45540 17900 45550
rect 17820 45530 17830 45540
rect 17670 45500 17830 45530
rect 17670 45480 17680 45500
rect 17600 45470 17680 45480
rect 17820 45480 17830 45500
rect 17890 45480 17900 45540
rect 18660 45540 18740 45550
rect 18660 45480 18670 45540
rect 18730 45530 18740 45540
rect 19040 45540 19120 45550
rect 19040 45530 19050 45540
rect 18730 45500 19050 45530
rect 18730 45480 18740 45500
rect 17820 45470 17900 45480
rect 18240 45470 18320 45480
rect 18660 45470 18740 45480
rect 19040 45480 19050 45500
rect 19110 45480 19120 45540
rect 19040 45470 19120 45480
rect 18240 45410 18250 45470
rect 18310 45430 18320 45470
rect 18310 45420 19010 45430
rect 18310 45410 18950 45420
rect 18240 45400 18950 45410
rect 18950 45350 19010 45360
rect 18890 44240 18950 44250
rect 18240 44210 18890 44220
rect 17620 44150 17680 44160
rect 18240 44150 18250 44210
rect 18310 44190 18890 44210
rect 18310 44150 18320 44190
rect 18890 44170 18950 44180
rect 19040 44150 19100 44160
rect 17820 44140 17900 44150
rect 18240 44140 18320 44150
rect 18660 44140 18740 44150
rect 17820 44130 17830 44140
rect 17680 44100 17830 44130
rect 17620 44080 17680 44090
rect 17820 44080 17830 44100
rect 17890 44080 17900 44140
rect 17820 44070 17900 44080
rect 18660 44080 18670 44140
rect 18730 44130 18740 44140
rect 18730 44100 19040 44130
rect 18730 44080 18740 44100
rect 19040 44080 19100 44090
rect 18660 44070 18740 44080
rect 18230 44050 18330 44060
rect 18230 43980 18250 44050
rect 18320 43980 18330 44050
rect 18230 43940 18330 43980
rect 18230 43870 18250 43940
rect 18320 43870 18330 43940
rect 18230 43850 18330 43870
rect 17600 43830 17680 43840
rect 17600 43770 17610 43830
rect 17670 43820 17680 43830
rect 17820 43830 17900 43840
rect 17820 43820 17830 43830
rect 17670 43790 17830 43820
rect 17670 43770 17680 43790
rect 17600 43760 17680 43770
rect 17820 43770 17830 43790
rect 17890 43770 17900 43830
rect 18660 43830 18740 43840
rect 18660 43770 18670 43830
rect 18730 43820 18740 43830
rect 19040 43830 19120 43840
rect 19040 43820 19050 43830
rect 18730 43790 19050 43820
rect 18730 43770 18740 43790
rect 17820 43760 17900 43770
rect 18240 43760 18320 43770
rect 18660 43760 18740 43770
rect 19040 43770 19050 43790
rect 19110 43770 19120 43830
rect 19040 43760 19120 43770
rect 18240 43700 18250 43760
rect 18310 43720 18320 43760
rect 18310 43710 19010 43720
rect 18310 43700 18950 43710
rect 18240 43690 18950 43700
rect 18950 43640 19010 43650
rect 18890 42530 18950 42540
rect 18240 42500 18890 42510
rect 17620 42440 17680 42450
rect 18240 42440 18250 42500
rect 18310 42480 18890 42500
rect 18310 42440 18320 42480
rect 18890 42460 18950 42470
rect 19040 42440 19100 42450
rect 17820 42430 17900 42440
rect 18240 42430 18320 42440
rect 18660 42430 18740 42440
rect 17820 42420 17830 42430
rect 17680 42390 17830 42420
rect 17620 42370 17680 42380
rect 17820 42370 17830 42390
rect 17890 42370 17900 42430
rect 17820 42360 17900 42370
rect 18660 42370 18670 42430
rect 18730 42420 18740 42430
rect 18730 42390 19040 42420
rect 18730 42370 18740 42390
rect 19040 42370 19100 42380
rect 18660 42360 18740 42370
rect 18230 42340 18330 42350
rect 18230 42270 18250 42340
rect 18320 42270 18330 42340
rect 18230 42230 18330 42270
rect 18230 42160 18250 42230
rect 18320 42160 18330 42230
rect 18230 42140 18330 42160
rect 17600 42120 17680 42130
rect 17600 42060 17610 42120
rect 17670 42110 17680 42120
rect 17820 42120 17900 42130
rect 17820 42110 17830 42120
rect 17670 42080 17830 42110
rect 17670 42060 17680 42080
rect 17600 42050 17680 42060
rect 17820 42060 17830 42080
rect 17890 42060 17900 42120
rect 18660 42120 18740 42130
rect 18660 42060 18670 42120
rect 18730 42110 18740 42120
rect 19040 42120 19120 42130
rect 19040 42110 19050 42120
rect 18730 42080 19050 42110
rect 18730 42060 18740 42080
rect 17820 42050 17900 42060
rect 18240 42050 18320 42060
rect 18660 42050 18740 42060
rect 19040 42060 19050 42080
rect 19110 42060 19120 42120
rect 19040 42050 19120 42060
rect 18240 41990 18250 42050
rect 18310 42010 18320 42050
rect 18310 42000 19010 42010
rect 18310 41990 18950 42000
rect 18240 41980 18950 41990
rect 18950 41930 19010 41940
rect 18890 40820 18950 40830
rect 18240 40790 18890 40800
rect 17620 40730 17680 40740
rect 18240 40730 18250 40790
rect 18310 40770 18890 40790
rect 18310 40730 18320 40770
rect 18890 40750 18950 40760
rect 19040 40730 19100 40740
rect 17820 40720 17900 40730
rect 18240 40720 18320 40730
rect 18660 40720 18740 40730
rect 17820 40710 17830 40720
rect 17680 40680 17830 40710
rect 17620 40660 17680 40670
rect 17820 40660 17830 40680
rect 17890 40660 17900 40720
rect 17820 40650 17900 40660
rect 18660 40660 18670 40720
rect 18730 40710 18740 40720
rect 18730 40680 19040 40710
rect 18730 40660 18740 40680
rect 19040 40660 19100 40670
rect 18660 40650 18740 40660
rect 18230 40630 18330 40640
rect 18230 40560 18250 40630
rect 18320 40560 18330 40630
rect 18230 40520 18330 40560
rect 18230 40450 18250 40520
rect 18320 40450 18330 40520
rect 18230 40430 18330 40450
rect 17600 40410 17680 40420
rect 17600 40350 17610 40410
rect 17670 40400 17680 40410
rect 17820 40410 17900 40420
rect 17820 40400 17830 40410
rect 17670 40370 17830 40400
rect 17670 40350 17680 40370
rect 17600 40340 17680 40350
rect 17820 40350 17830 40370
rect 17890 40350 17900 40410
rect 18660 40410 18740 40420
rect 18660 40350 18670 40410
rect 18730 40400 18740 40410
rect 19040 40410 19120 40420
rect 19040 40400 19050 40410
rect 18730 40370 19050 40400
rect 18730 40350 18740 40370
rect 17820 40340 17900 40350
rect 18240 40340 18320 40350
rect 18660 40340 18740 40350
rect 19040 40350 19050 40370
rect 19110 40350 19120 40410
rect 19040 40340 19120 40350
rect 14170 39270 14400 39300
rect 14050 39210 14220 39240
rect 13790 38690 13870 38700
rect 13790 38630 13800 38690
rect 13860 38630 13870 38690
rect 13940 38640 13950 38700
rect 14010 38640 14020 38700
rect 13790 38620 13870 38630
rect 14190 36320 14220 39210
rect 14250 39230 14310 39240
rect 14250 39160 14310 39170
rect 12490 36310 12570 36320
rect 12490 36250 12500 36310
rect 12560 36250 12570 36310
rect 14170 36260 14180 36320
rect 14240 36260 14250 36320
rect 12490 36240 12570 36250
rect 14280 36180 14310 39160
rect 14370 36600 14400 39270
rect 14430 39290 14490 39300
rect 14430 39220 14490 39230
rect 14350 36540 14360 36600
rect 14420 36540 14430 36600
rect 14460 36460 14490 39220
rect 14410 36400 14420 36460
rect 14480 36400 14490 36460
rect 17240 39290 17300 39300
rect 17240 39220 17300 39230
rect 17330 39270 17560 39300
rect 17240 36460 17270 39220
rect 17330 36600 17360 39270
rect 17650 39240 17680 40340
rect 18240 40280 18250 40340
rect 18310 40300 18320 40340
rect 18310 40290 19010 40300
rect 18310 40280 18950 40290
rect 18240 40270 18950 40280
rect 18950 40220 19010 40230
rect 17420 39230 17480 39240
rect 17420 39160 17480 39170
rect 17510 39210 17680 39240
rect 17710 39680 17790 39690
rect 17710 39620 17720 39680
rect 17780 39620 17790 39680
rect 18780 39680 18860 39690
rect 18780 39620 18790 39680
rect 18850 39620 18860 39680
rect 17300 36590 17380 36600
rect 17300 36530 17310 36590
rect 17370 36530 17380 36590
rect 17300 36520 17380 36530
rect 17240 36450 17320 36460
rect 17240 36390 17250 36450
rect 17310 36390 17320 36450
rect 17240 36380 17320 36390
rect 12430 36170 12510 36180
rect 7440 36100 7520 36110
rect 12430 36110 12440 36170
rect 12500 36110 12510 36170
rect 14230 36120 14240 36180
rect 14300 36120 14310 36180
rect 17420 36180 17450 39160
rect 17510 36320 17540 39210
rect 17710 38840 17780 39620
rect 18780 39610 18860 39620
rect 18950 39680 19010 39690
rect 18950 39610 19010 39620
rect 17710 38830 17790 38840
rect 17710 38770 17720 38830
rect 17780 38770 17790 38830
rect 17710 38760 17790 38770
rect 18790 38700 18860 39610
rect 18980 38700 19010 39610
rect 19040 39240 19070 40340
rect 19160 39300 19190 47180
rect 22280 39420 22310 48890
rect 23230 48830 23240 48890
rect 23300 48850 23310 48890
rect 23300 48840 24000 48850
rect 23300 48830 23940 48840
rect 23230 48820 23940 48830
rect 23940 48770 24000 48780
rect 23880 47660 23940 47670
rect 23230 47630 23880 47640
rect 22370 47570 22430 47580
rect 23230 47570 23240 47630
rect 23300 47610 23880 47630
rect 23300 47570 23310 47610
rect 23880 47590 23940 47600
rect 24270 47570 24330 47580
rect 22810 47560 22890 47570
rect 23230 47560 23310 47570
rect 23650 47560 23730 47570
rect 22810 47550 22820 47560
rect 22430 47520 22820 47550
rect 22370 47500 22430 47510
rect 22810 47500 22820 47520
rect 22880 47500 22890 47560
rect 22810 47490 22890 47500
rect 23650 47500 23660 47560
rect 23720 47550 23730 47560
rect 23720 47520 24270 47550
rect 23720 47500 23730 47520
rect 24270 47500 24330 47510
rect 23650 47490 23730 47500
rect 23220 47470 23320 47480
rect 23220 47400 23240 47470
rect 23310 47400 23320 47470
rect 23220 47360 23320 47400
rect 23220 47290 23240 47360
rect 23310 47290 23320 47360
rect 23220 47270 23320 47290
rect 22350 47250 22430 47260
rect 22350 47190 22360 47250
rect 22420 47240 22430 47250
rect 22810 47250 22890 47260
rect 22810 47240 22820 47250
rect 22420 47210 22820 47240
rect 22420 47190 22430 47210
rect 22350 47180 22430 47190
rect 22810 47190 22820 47210
rect 22880 47190 22890 47250
rect 23650 47250 23730 47260
rect 23650 47190 23660 47250
rect 23720 47240 23730 47250
rect 24270 47250 24350 47260
rect 24270 47240 24280 47250
rect 23720 47210 24280 47240
rect 23720 47190 23730 47210
rect 22810 47180 22890 47190
rect 23230 47180 23310 47190
rect 23650 47180 23730 47190
rect 24270 47190 24280 47210
rect 24340 47190 24350 47250
rect 24270 47180 24350 47190
rect 21870 39410 21930 39420
rect 21870 39340 21930 39350
rect 21960 39390 22310 39420
rect 19160 39270 19390 39300
rect 19040 39210 19210 39240
rect 18780 38690 18860 38700
rect 18780 38630 18790 38690
rect 18850 38630 18860 38690
rect 18930 38640 18940 38700
rect 19000 38640 19010 38700
rect 18780 38620 18860 38630
rect 19180 36320 19210 39210
rect 19240 39230 19300 39240
rect 19240 39160 19300 39170
rect 17480 36310 17560 36320
rect 17480 36250 17490 36310
rect 17550 36250 17560 36310
rect 19160 36260 19170 36320
rect 19230 36260 19240 36320
rect 17480 36240 17560 36250
rect 19270 36180 19300 39160
rect 19360 36600 19390 39270
rect 19420 39290 19480 39300
rect 19420 39220 19480 39230
rect 19340 36540 19350 36600
rect 19410 36540 19420 36600
rect 19450 36460 19480 39220
rect 21870 36740 21900 39340
rect 21960 36880 21990 39390
rect 22400 39360 22430 47180
rect 23230 47120 23240 47180
rect 23300 47140 23310 47180
rect 23300 47130 24000 47140
rect 23300 47120 23940 47130
rect 23230 47110 23940 47120
rect 23940 47060 24000 47070
rect 23880 45950 23940 45960
rect 23230 45920 23880 45930
rect 22490 45860 22550 45870
rect 23230 45860 23240 45920
rect 23300 45900 23880 45920
rect 23300 45860 23310 45900
rect 23880 45880 23940 45890
rect 24150 45860 24210 45870
rect 22810 45850 22890 45860
rect 23230 45850 23310 45860
rect 23650 45850 23730 45860
rect 22810 45840 22820 45850
rect 22550 45810 22820 45840
rect 22490 45790 22550 45800
rect 22810 45790 22820 45810
rect 22880 45790 22890 45850
rect 22810 45780 22890 45790
rect 23650 45790 23660 45850
rect 23720 45840 23730 45850
rect 23720 45810 24150 45840
rect 23720 45790 23730 45810
rect 24150 45790 24210 45800
rect 23650 45780 23730 45790
rect 23220 45760 23320 45770
rect 23220 45690 23240 45760
rect 23310 45690 23320 45760
rect 23220 45650 23320 45690
rect 23220 45580 23240 45650
rect 23310 45580 23320 45650
rect 23220 45560 23320 45580
rect 22470 45540 22550 45550
rect 22470 45480 22480 45540
rect 22540 45530 22550 45540
rect 22810 45540 22890 45550
rect 22810 45530 22820 45540
rect 22540 45500 22820 45530
rect 22540 45480 22550 45500
rect 22470 45470 22550 45480
rect 22810 45480 22820 45500
rect 22880 45480 22890 45540
rect 23650 45540 23730 45550
rect 23650 45480 23660 45540
rect 23720 45530 23730 45540
rect 24150 45540 24230 45550
rect 24150 45530 24160 45540
rect 23720 45500 24160 45530
rect 23720 45480 23730 45500
rect 22810 45470 22890 45480
rect 23230 45470 23310 45480
rect 23650 45470 23730 45480
rect 24150 45480 24160 45500
rect 24220 45480 24230 45540
rect 24150 45470 24230 45480
rect 23230 45410 23240 45470
rect 23300 45430 23310 45470
rect 23300 45420 24000 45430
rect 23300 45410 23940 45420
rect 23230 45400 23940 45410
rect 23940 45350 24000 45360
rect 23880 44240 23940 44250
rect 23230 44210 23880 44220
rect 22490 44150 22550 44160
rect 23230 44150 23240 44210
rect 23300 44190 23880 44210
rect 23300 44150 23310 44190
rect 23880 44170 23940 44180
rect 24150 44150 24210 44160
rect 22810 44140 22890 44150
rect 23230 44140 23310 44150
rect 23650 44140 23730 44150
rect 22810 44130 22820 44140
rect 22550 44100 22820 44130
rect 22490 44080 22550 44090
rect 22810 44080 22820 44100
rect 22880 44080 22890 44140
rect 22810 44070 22890 44080
rect 23650 44080 23660 44140
rect 23720 44130 23730 44140
rect 23720 44100 24150 44130
rect 23720 44080 23730 44100
rect 24150 44080 24210 44090
rect 23650 44070 23730 44080
rect 23220 44050 23320 44060
rect 23220 43980 23240 44050
rect 23310 43980 23320 44050
rect 23220 43940 23320 43980
rect 23220 43870 23240 43940
rect 23310 43870 23320 43940
rect 23220 43850 23320 43870
rect 22470 43830 22550 43840
rect 22470 43770 22480 43830
rect 22540 43820 22550 43830
rect 22810 43830 22890 43840
rect 22810 43820 22820 43830
rect 22540 43790 22820 43820
rect 22540 43770 22550 43790
rect 22470 43760 22550 43770
rect 22810 43770 22820 43790
rect 22880 43770 22890 43830
rect 23650 43830 23730 43840
rect 23650 43770 23660 43830
rect 23720 43820 23730 43830
rect 24150 43830 24230 43840
rect 24150 43820 24160 43830
rect 23720 43790 24160 43820
rect 23720 43770 23730 43790
rect 22810 43760 22890 43770
rect 23230 43760 23310 43770
rect 23650 43760 23730 43770
rect 24150 43770 24160 43790
rect 24220 43770 24230 43830
rect 24150 43760 24230 43770
rect 22050 39350 22110 39360
rect 22050 39280 22110 39290
rect 22140 39330 22430 39360
rect 22050 37020 22080 39280
rect 22140 37160 22170 39330
rect 22520 39300 22550 43760
rect 23230 43700 23240 43760
rect 23300 43720 23310 43760
rect 23300 43710 24000 43720
rect 23300 43700 23940 43710
rect 23230 43690 23940 43700
rect 23940 43640 24000 43650
rect 23880 42530 23940 42540
rect 23230 42500 23880 42510
rect 22610 42440 22670 42450
rect 23230 42440 23240 42500
rect 23300 42480 23880 42500
rect 23300 42440 23310 42480
rect 23880 42460 23940 42470
rect 24030 42440 24090 42450
rect 22810 42430 22890 42440
rect 23230 42430 23310 42440
rect 23650 42430 23730 42440
rect 22810 42420 22820 42430
rect 22670 42390 22820 42420
rect 22610 42370 22670 42380
rect 22810 42370 22820 42390
rect 22880 42370 22890 42430
rect 22810 42360 22890 42370
rect 23650 42370 23660 42430
rect 23720 42420 23730 42430
rect 23720 42390 24030 42420
rect 23720 42370 23730 42390
rect 24030 42370 24090 42380
rect 23650 42360 23730 42370
rect 23220 42340 23320 42350
rect 23220 42270 23240 42340
rect 23310 42270 23320 42340
rect 23220 42230 23320 42270
rect 23220 42160 23240 42230
rect 23310 42160 23320 42230
rect 23220 42140 23320 42160
rect 22590 42120 22670 42130
rect 22590 42060 22600 42120
rect 22660 42110 22670 42120
rect 22810 42120 22890 42130
rect 22810 42110 22820 42120
rect 22660 42080 22820 42110
rect 22660 42060 22670 42080
rect 22590 42050 22670 42060
rect 22810 42060 22820 42080
rect 22880 42060 22890 42120
rect 23650 42120 23730 42130
rect 23650 42060 23660 42120
rect 23720 42110 23730 42120
rect 24030 42120 24110 42130
rect 24030 42110 24040 42120
rect 23720 42080 24040 42110
rect 23720 42060 23730 42080
rect 22810 42050 22890 42060
rect 23230 42050 23310 42060
rect 23650 42050 23730 42060
rect 24030 42060 24040 42080
rect 24100 42060 24110 42120
rect 24030 42050 24110 42060
rect 23230 41990 23240 42050
rect 23300 42010 23310 42050
rect 23300 42000 24000 42010
rect 23300 41990 23940 42000
rect 23230 41980 23940 41990
rect 23940 41930 24000 41940
rect 23880 40820 23940 40830
rect 23230 40790 23880 40800
rect 22610 40730 22670 40740
rect 23230 40730 23240 40790
rect 23300 40770 23880 40790
rect 23300 40730 23310 40770
rect 23880 40750 23940 40760
rect 24030 40730 24090 40740
rect 22810 40720 22890 40730
rect 23230 40720 23310 40730
rect 23650 40720 23730 40730
rect 22810 40710 22820 40720
rect 22670 40680 22820 40710
rect 22610 40660 22670 40670
rect 22810 40660 22820 40680
rect 22880 40660 22890 40720
rect 22810 40650 22890 40660
rect 23650 40660 23660 40720
rect 23720 40710 23730 40720
rect 23720 40680 24030 40710
rect 23720 40660 23730 40680
rect 24030 40660 24090 40670
rect 23650 40650 23730 40660
rect 23220 40630 23320 40640
rect 23220 40560 23240 40630
rect 23310 40560 23320 40630
rect 23220 40520 23320 40560
rect 23220 40450 23240 40520
rect 23310 40450 23320 40520
rect 23220 40430 23320 40450
rect 22590 40410 22670 40420
rect 22590 40350 22600 40410
rect 22660 40400 22670 40410
rect 22810 40410 22890 40420
rect 22810 40400 22820 40410
rect 22660 40370 22820 40400
rect 22660 40350 22670 40370
rect 22590 40340 22670 40350
rect 22810 40350 22820 40370
rect 22880 40350 22890 40410
rect 23650 40410 23730 40420
rect 23650 40350 23660 40410
rect 23720 40400 23730 40410
rect 24030 40410 24110 40420
rect 24030 40400 24040 40410
rect 23720 40370 24040 40400
rect 23720 40350 23730 40370
rect 22810 40340 22890 40350
rect 23230 40340 23310 40350
rect 23650 40340 23730 40350
rect 24030 40350 24040 40370
rect 24100 40350 24110 40410
rect 24030 40340 24110 40350
rect 22230 39290 22290 39300
rect 22230 39220 22290 39230
rect 22320 39270 22550 39300
rect 22110 37150 22190 37160
rect 22110 37090 22120 37150
rect 22180 37090 22190 37150
rect 22110 37080 22190 37090
rect 22050 37010 22130 37020
rect 22050 36950 22060 37010
rect 22120 36950 22130 37010
rect 22050 36940 22130 36950
rect 21930 36870 22010 36880
rect 21930 36810 21940 36870
rect 22000 36810 22010 36870
rect 21930 36800 22010 36810
rect 21870 36730 21950 36740
rect 21870 36670 21880 36730
rect 21940 36670 21950 36730
rect 21870 36660 21950 36670
rect 19400 36400 19410 36460
rect 19470 36400 19480 36460
rect 22230 36460 22260 39220
rect 22320 36600 22350 39270
rect 22640 39240 22670 40340
rect 23230 40280 23240 40340
rect 23300 40300 23310 40340
rect 23300 40290 24000 40300
rect 23300 40280 23940 40290
rect 23230 40270 23940 40280
rect 23940 40220 24000 40230
rect 22410 39230 22470 39240
rect 22410 39160 22470 39170
rect 22500 39210 22670 39240
rect 22700 39680 22780 39690
rect 22700 39620 22710 39680
rect 22770 39620 22780 39680
rect 23770 39680 23850 39690
rect 23770 39620 23780 39680
rect 23840 39620 23850 39680
rect 22290 36590 22370 36600
rect 22290 36530 22300 36590
rect 22360 36530 22370 36590
rect 22290 36520 22370 36530
rect 22230 36450 22310 36460
rect 22230 36390 22240 36450
rect 22300 36390 22310 36450
rect 22230 36380 22310 36390
rect 17420 36170 17500 36180
rect 12430 36100 12510 36110
rect 17420 36110 17430 36170
rect 17490 36110 17500 36170
rect 19220 36120 19230 36180
rect 19290 36120 19300 36180
rect 22410 36180 22440 39160
rect 22500 36320 22530 39210
rect 22700 38840 22770 39620
rect 23770 39610 23850 39620
rect 23940 39680 24000 39690
rect 23940 39610 24000 39620
rect 22700 38830 22780 38840
rect 22700 38770 22710 38830
rect 22770 38770 22780 38830
rect 22700 38760 22780 38770
rect 23780 38700 23850 39610
rect 23970 38700 24000 39610
rect 24030 39240 24060 40340
rect 24150 39300 24180 43760
rect 24270 39360 24300 47180
rect 24390 39420 24420 48890
rect 27270 39420 27300 48890
rect 28220 48830 28230 48890
rect 28290 48850 28300 48890
rect 28290 48840 28990 48850
rect 28290 48830 28930 48840
rect 28220 48820 28930 48830
rect 28930 48770 28990 48780
rect 28870 47660 28930 47670
rect 28220 47630 28870 47640
rect 27360 47570 27420 47580
rect 28220 47570 28230 47630
rect 28290 47610 28870 47630
rect 28290 47570 28300 47610
rect 28870 47590 28930 47600
rect 29260 47570 29320 47580
rect 27800 47560 27880 47570
rect 28220 47560 28300 47570
rect 28640 47560 28720 47570
rect 27800 47550 27810 47560
rect 27420 47520 27810 47550
rect 27360 47500 27420 47510
rect 27800 47500 27810 47520
rect 27870 47500 27880 47560
rect 27800 47490 27880 47500
rect 28640 47500 28650 47560
rect 28710 47550 28720 47560
rect 28710 47520 29260 47550
rect 28710 47500 28720 47520
rect 29260 47500 29320 47510
rect 28640 47490 28720 47500
rect 28210 47470 28310 47480
rect 28210 47400 28230 47470
rect 28300 47400 28310 47470
rect 28210 47360 28310 47400
rect 28210 47290 28230 47360
rect 28300 47290 28310 47360
rect 28210 47270 28310 47290
rect 27340 47250 27420 47260
rect 27340 47190 27350 47250
rect 27410 47240 27420 47250
rect 27800 47250 27880 47260
rect 27800 47240 27810 47250
rect 27410 47210 27810 47240
rect 27410 47190 27420 47210
rect 27340 47180 27420 47190
rect 27800 47190 27810 47210
rect 27870 47190 27880 47250
rect 28640 47250 28720 47260
rect 28640 47190 28650 47250
rect 28710 47240 28720 47250
rect 29260 47250 29340 47260
rect 29260 47240 29270 47250
rect 28710 47210 29270 47240
rect 28710 47190 28720 47210
rect 27800 47180 27880 47190
rect 28220 47180 28300 47190
rect 28640 47180 28720 47190
rect 29260 47190 29270 47210
rect 29330 47190 29340 47250
rect 29260 47180 29340 47190
rect 24390 39390 24740 39420
rect 24270 39330 24560 39360
rect 24150 39270 24380 39300
rect 24030 39210 24200 39240
rect 23770 38690 23850 38700
rect 23770 38630 23780 38690
rect 23840 38630 23850 38690
rect 23920 38640 23930 38700
rect 23990 38640 24000 38700
rect 23770 38620 23850 38630
rect 24170 36320 24200 39210
rect 24230 39230 24290 39240
rect 24230 39160 24290 39170
rect 22470 36310 22550 36320
rect 22470 36250 22480 36310
rect 22540 36250 22550 36310
rect 24150 36260 24160 36320
rect 24220 36260 24230 36320
rect 22470 36240 22550 36250
rect 24260 36180 24290 39160
rect 24350 36600 24380 39270
rect 24410 39290 24470 39300
rect 24410 39220 24470 39230
rect 24330 36540 24340 36600
rect 24400 36540 24410 36600
rect 24440 36460 24470 39220
rect 24530 37160 24560 39330
rect 24590 39350 24650 39360
rect 24590 39280 24650 39290
rect 24510 37100 24520 37160
rect 24580 37100 24590 37160
rect 24620 37020 24650 39280
rect 24570 36960 24580 37020
rect 24640 36960 24650 37020
rect 24710 36880 24740 39390
rect 24770 39410 24830 39420
rect 24770 39340 24830 39350
rect 24690 36820 24700 36880
rect 24760 36820 24770 36880
rect 24800 36740 24830 39340
rect 24750 36680 24760 36740
rect 24820 36680 24830 36740
rect 26860 39410 26920 39420
rect 26860 39340 26920 39350
rect 26950 39390 27300 39420
rect 26860 36740 26890 39340
rect 26950 36880 26980 39390
rect 27390 39360 27420 47180
rect 28220 47120 28230 47180
rect 28290 47140 28300 47180
rect 28290 47130 28990 47140
rect 28290 47120 28930 47130
rect 28220 47110 28930 47120
rect 28930 47060 28990 47070
rect 28870 45950 28930 45960
rect 28220 45920 28870 45930
rect 27480 45860 27540 45870
rect 28220 45860 28230 45920
rect 28290 45900 28870 45920
rect 28290 45860 28300 45900
rect 28870 45880 28930 45890
rect 29140 45860 29200 45870
rect 27800 45850 27880 45860
rect 28220 45850 28300 45860
rect 28640 45850 28720 45860
rect 27800 45840 27810 45850
rect 27540 45810 27810 45840
rect 27480 45790 27540 45800
rect 27800 45790 27810 45810
rect 27870 45790 27880 45850
rect 27800 45780 27880 45790
rect 28640 45790 28650 45850
rect 28710 45840 28720 45850
rect 28710 45810 29140 45840
rect 28710 45790 28720 45810
rect 29140 45790 29200 45800
rect 28640 45780 28720 45790
rect 28210 45760 28310 45770
rect 28210 45690 28230 45760
rect 28300 45690 28310 45760
rect 28210 45650 28310 45690
rect 28210 45580 28230 45650
rect 28300 45580 28310 45650
rect 28210 45560 28310 45580
rect 27460 45540 27540 45550
rect 27460 45480 27470 45540
rect 27530 45530 27540 45540
rect 27800 45540 27880 45550
rect 27800 45530 27810 45540
rect 27530 45500 27810 45530
rect 27530 45480 27540 45500
rect 27460 45470 27540 45480
rect 27800 45480 27810 45500
rect 27870 45480 27880 45540
rect 28640 45540 28720 45550
rect 28640 45480 28650 45540
rect 28710 45530 28720 45540
rect 29140 45540 29220 45550
rect 29140 45530 29150 45540
rect 28710 45500 29150 45530
rect 28710 45480 28720 45500
rect 27800 45470 27880 45480
rect 28220 45470 28300 45480
rect 28640 45470 28720 45480
rect 29140 45480 29150 45500
rect 29210 45480 29220 45540
rect 29140 45470 29220 45480
rect 28220 45410 28230 45470
rect 28290 45430 28300 45470
rect 28290 45420 28990 45430
rect 28290 45410 28930 45420
rect 28220 45400 28930 45410
rect 28930 45350 28990 45360
rect 28870 44240 28930 44250
rect 28220 44210 28870 44220
rect 27480 44150 27540 44160
rect 28220 44150 28230 44210
rect 28290 44190 28870 44210
rect 28290 44150 28300 44190
rect 28870 44170 28930 44180
rect 29140 44150 29200 44160
rect 27800 44140 27880 44150
rect 28220 44140 28300 44150
rect 28640 44140 28720 44150
rect 27800 44130 27810 44140
rect 27540 44100 27810 44130
rect 27480 44080 27540 44090
rect 27800 44080 27810 44100
rect 27870 44080 27880 44140
rect 27800 44070 27880 44080
rect 28640 44080 28650 44140
rect 28710 44130 28720 44140
rect 28710 44100 29140 44130
rect 28710 44080 28720 44100
rect 29140 44080 29200 44090
rect 28640 44070 28720 44080
rect 28210 44050 28310 44060
rect 28210 43980 28230 44050
rect 28300 43980 28310 44050
rect 28210 43940 28310 43980
rect 28210 43870 28230 43940
rect 28300 43870 28310 43940
rect 28210 43850 28310 43870
rect 27460 43830 27540 43840
rect 27460 43770 27470 43830
rect 27530 43820 27540 43830
rect 27800 43830 27880 43840
rect 27800 43820 27810 43830
rect 27530 43790 27810 43820
rect 27530 43770 27540 43790
rect 27460 43760 27540 43770
rect 27800 43770 27810 43790
rect 27870 43770 27880 43830
rect 28640 43830 28720 43840
rect 28640 43770 28650 43830
rect 28710 43820 28720 43830
rect 29140 43830 29220 43840
rect 29140 43820 29150 43830
rect 28710 43790 29150 43820
rect 28710 43770 28720 43790
rect 27800 43760 27880 43770
rect 28220 43760 28300 43770
rect 28640 43760 28720 43770
rect 29140 43770 29150 43790
rect 29210 43770 29220 43830
rect 29140 43760 29220 43770
rect 27040 39350 27100 39360
rect 27040 39280 27100 39290
rect 27130 39330 27420 39360
rect 27040 37020 27070 39280
rect 27130 37160 27160 39330
rect 27510 39300 27540 43760
rect 28220 43700 28230 43760
rect 28290 43720 28300 43760
rect 28290 43710 28990 43720
rect 28290 43700 28930 43710
rect 28220 43690 28930 43700
rect 28930 43640 28990 43650
rect 28870 42530 28930 42540
rect 28220 42500 28870 42510
rect 27600 42440 27660 42450
rect 28220 42440 28230 42500
rect 28290 42480 28870 42500
rect 28290 42440 28300 42480
rect 28870 42460 28930 42470
rect 29020 42440 29080 42450
rect 27800 42430 27880 42440
rect 28220 42430 28300 42440
rect 28640 42430 28720 42440
rect 27800 42420 27810 42430
rect 27660 42390 27810 42420
rect 27600 42370 27660 42380
rect 27800 42370 27810 42390
rect 27870 42370 27880 42430
rect 27800 42360 27880 42370
rect 28640 42370 28650 42430
rect 28710 42420 28720 42430
rect 28710 42390 29020 42420
rect 28710 42370 28720 42390
rect 29020 42370 29080 42380
rect 28640 42360 28720 42370
rect 28210 42340 28310 42350
rect 28210 42270 28230 42340
rect 28300 42270 28310 42340
rect 28210 42230 28310 42270
rect 28210 42160 28230 42230
rect 28300 42160 28310 42230
rect 28210 42140 28310 42160
rect 27580 42120 27660 42130
rect 27580 42060 27590 42120
rect 27650 42110 27660 42120
rect 27800 42120 27880 42130
rect 27800 42110 27810 42120
rect 27650 42080 27810 42110
rect 27650 42060 27660 42080
rect 27580 42050 27660 42060
rect 27800 42060 27810 42080
rect 27870 42060 27880 42120
rect 28640 42120 28720 42130
rect 28640 42060 28650 42120
rect 28710 42110 28720 42120
rect 29020 42120 29100 42130
rect 29020 42110 29030 42120
rect 28710 42080 29030 42110
rect 28710 42060 28720 42080
rect 27800 42050 27880 42060
rect 28220 42050 28300 42060
rect 28640 42050 28720 42060
rect 29020 42060 29030 42080
rect 29090 42060 29100 42120
rect 29020 42050 29100 42060
rect 28220 41990 28230 42050
rect 28290 42010 28300 42050
rect 28290 42000 28990 42010
rect 28290 41990 28930 42000
rect 28220 41980 28930 41990
rect 28930 41930 28990 41940
rect 28870 40820 28930 40830
rect 28220 40790 28870 40800
rect 27600 40730 27660 40740
rect 28220 40730 28230 40790
rect 28290 40770 28870 40790
rect 28290 40730 28300 40770
rect 28870 40750 28930 40760
rect 29020 40730 29080 40740
rect 27800 40720 27880 40730
rect 28220 40720 28300 40730
rect 28640 40720 28720 40730
rect 27800 40710 27810 40720
rect 27660 40680 27810 40710
rect 27600 40660 27660 40670
rect 27800 40660 27810 40680
rect 27870 40660 27880 40720
rect 27800 40650 27880 40660
rect 28640 40660 28650 40720
rect 28710 40710 28720 40720
rect 28710 40680 29020 40710
rect 28710 40660 28720 40680
rect 29020 40660 29080 40670
rect 28640 40650 28720 40660
rect 28210 40630 28310 40640
rect 28210 40560 28230 40630
rect 28300 40560 28310 40630
rect 28210 40520 28310 40560
rect 28210 40450 28230 40520
rect 28300 40450 28310 40520
rect 28210 40430 28310 40450
rect 27580 40410 27660 40420
rect 27580 40350 27590 40410
rect 27650 40400 27660 40410
rect 27800 40410 27880 40420
rect 27800 40400 27810 40410
rect 27650 40370 27810 40400
rect 27650 40350 27660 40370
rect 27580 40340 27660 40350
rect 27800 40350 27810 40370
rect 27870 40350 27880 40410
rect 28640 40410 28720 40420
rect 28640 40350 28650 40410
rect 28710 40400 28720 40410
rect 29020 40410 29100 40420
rect 29020 40400 29030 40410
rect 28710 40370 29030 40400
rect 28710 40350 28720 40370
rect 27800 40340 27880 40350
rect 28220 40340 28300 40350
rect 28640 40340 28720 40350
rect 29020 40350 29030 40370
rect 29090 40350 29100 40410
rect 29020 40340 29100 40350
rect 27220 39290 27280 39300
rect 27220 39220 27280 39230
rect 27310 39270 27540 39300
rect 27100 37150 27180 37160
rect 27100 37090 27110 37150
rect 27170 37090 27180 37150
rect 27100 37080 27180 37090
rect 27040 37010 27120 37020
rect 27040 36950 27050 37010
rect 27110 36950 27120 37010
rect 27040 36940 27120 36950
rect 26920 36870 27000 36880
rect 26920 36810 26930 36870
rect 26990 36810 27000 36870
rect 26920 36800 27000 36810
rect 26860 36730 26940 36740
rect 26860 36670 26870 36730
rect 26930 36670 26940 36730
rect 26860 36660 26940 36670
rect 24390 36400 24400 36460
rect 24460 36400 24470 36460
rect 27220 36460 27250 39220
rect 27310 36600 27340 39270
rect 27630 39240 27660 40340
rect 28220 40280 28230 40340
rect 28290 40300 28300 40340
rect 28290 40290 28990 40300
rect 28290 40280 28930 40290
rect 28220 40270 28930 40280
rect 28930 40220 28990 40230
rect 27400 39230 27460 39240
rect 27400 39160 27460 39170
rect 27490 39210 27660 39240
rect 27690 39680 27770 39690
rect 27690 39620 27700 39680
rect 27760 39620 27770 39680
rect 28760 39680 28840 39690
rect 28760 39620 28770 39680
rect 28830 39620 28840 39680
rect 27280 36590 27360 36600
rect 27280 36530 27290 36590
rect 27350 36530 27360 36590
rect 27280 36520 27360 36530
rect 27220 36450 27300 36460
rect 27220 36390 27230 36450
rect 27290 36390 27300 36450
rect 27220 36380 27300 36390
rect 22410 36170 22490 36180
rect 17420 36100 17500 36110
rect 22410 36110 22420 36170
rect 22480 36110 22490 36170
rect 24210 36120 24220 36180
rect 24280 36120 24290 36180
rect 27400 36180 27430 39160
rect 27490 36320 27520 39210
rect 27690 38840 27760 39620
rect 28760 39610 28840 39620
rect 28930 39680 28990 39690
rect 28930 39610 28990 39620
rect 27690 38830 27770 38840
rect 27690 38770 27700 38830
rect 27760 38770 27770 38830
rect 27690 38760 27770 38770
rect 28770 38700 28840 39610
rect 28960 38700 28990 39610
rect 29020 39240 29050 40340
rect 29140 39300 29170 43760
rect 29260 39360 29290 47180
rect 29380 39420 29410 48890
rect 32020 39540 32050 52310
rect 33210 52250 33220 52310
rect 33280 52270 33290 52310
rect 33280 52260 33980 52270
rect 33280 52250 33920 52260
rect 33210 52240 33920 52250
rect 33920 52190 33980 52200
rect 33860 51080 33920 51090
rect 33210 51050 33860 51060
rect 32110 50990 32170 51000
rect 33210 50990 33220 51050
rect 33280 51030 33860 51050
rect 33280 50990 33290 51030
rect 33860 51010 33920 51020
rect 34490 50990 34550 51000
rect 32790 50980 32870 50990
rect 33210 50980 33290 50990
rect 33630 50980 33710 50990
rect 32790 50970 32800 50980
rect 32170 50940 32800 50970
rect 32110 50920 32170 50930
rect 32790 50920 32800 50940
rect 32860 50920 32870 50980
rect 32790 50910 32870 50920
rect 33630 50920 33640 50980
rect 33700 50970 33710 50980
rect 33700 50940 34490 50970
rect 33700 50920 33710 50940
rect 34490 50920 34550 50930
rect 33630 50910 33710 50920
rect 33200 50890 33300 50900
rect 33200 50820 33220 50890
rect 33290 50820 33300 50890
rect 33200 50780 33300 50820
rect 33200 50710 33220 50780
rect 33290 50710 33300 50780
rect 33200 50690 33300 50710
rect 32090 50670 32170 50680
rect 32090 50610 32100 50670
rect 32160 50660 32170 50670
rect 32790 50670 32870 50680
rect 32790 50660 32800 50670
rect 32160 50630 32800 50660
rect 32160 50610 32170 50630
rect 32090 50600 32170 50610
rect 32790 50610 32800 50630
rect 32860 50610 32870 50670
rect 33630 50670 33710 50680
rect 33630 50610 33640 50670
rect 33700 50660 33710 50670
rect 34490 50670 34570 50680
rect 34490 50660 34500 50670
rect 33700 50630 34500 50660
rect 33700 50610 33710 50630
rect 32790 50600 32870 50610
rect 33210 50600 33290 50610
rect 33630 50600 33710 50610
rect 34490 50610 34500 50630
rect 34560 50610 34570 50670
rect 34490 50600 34570 50610
rect 31490 39530 31550 39540
rect 31490 39460 31550 39470
rect 31580 39510 32050 39540
rect 29380 39390 29730 39420
rect 29260 39330 29550 39360
rect 29140 39270 29370 39300
rect 29020 39210 29190 39240
rect 28760 38690 28840 38700
rect 28760 38630 28770 38690
rect 28830 38630 28840 38690
rect 28910 38640 28920 38700
rect 28980 38640 28990 38700
rect 28760 38620 28840 38630
rect 29160 36320 29190 39210
rect 29220 39230 29280 39240
rect 29220 39160 29280 39170
rect 27460 36310 27540 36320
rect 27460 36250 27470 36310
rect 27530 36250 27540 36310
rect 29140 36260 29150 36320
rect 29210 36260 29220 36320
rect 27460 36240 27540 36250
rect 29250 36180 29280 39160
rect 29340 36600 29370 39270
rect 29400 39290 29460 39300
rect 29400 39220 29460 39230
rect 29320 36540 29330 36600
rect 29390 36540 29400 36600
rect 29430 36460 29460 39220
rect 29520 37160 29550 39330
rect 29580 39350 29640 39360
rect 29580 39280 29640 39290
rect 29500 37100 29510 37160
rect 29570 37100 29580 37160
rect 29610 37020 29640 39280
rect 29560 36960 29570 37020
rect 29630 36960 29640 37020
rect 29700 36880 29730 39390
rect 29760 39410 29820 39420
rect 29760 39340 29820 39350
rect 29680 36820 29690 36880
rect 29750 36820 29760 36880
rect 29790 36740 29820 39340
rect 31490 37300 31520 39460
rect 31580 37440 31610 39510
rect 32140 39480 32170 50600
rect 33210 50540 33220 50600
rect 33280 50560 33290 50600
rect 33280 50550 33980 50560
rect 33280 50540 33920 50550
rect 33210 50530 33920 50540
rect 33920 50480 33980 50490
rect 33860 49370 33920 49380
rect 33210 49340 33860 49350
rect 32230 49280 32290 49290
rect 33210 49280 33220 49340
rect 33280 49320 33860 49340
rect 33280 49280 33290 49320
rect 33860 49300 33920 49310
rect 34370 49280 34430 49290
rect 32790 49270 32870 49280
rect 33210 49270 33290 49280
rect 33630 49270 33710 49280
rect 32790 49260 32800 49270
rect 32290 49230 32800 49260
rect 32230 49210 32290 49220
rect 32790 49210 32800 49230
rect 32860 49210 32870 49270
rect 32790 49200 32870 49210
rect 33630 49210 33640 49270
rect 33700 49260 33710 49270
rect 33700 49230 34370 49260
rect 33700 49210 33710 49230
rect 34370 49210 34430 49220
rect 33630 49200 33710 49210
rect 33200 49180 33300 49190
rect 33200 49110 33220 49180
rect 33290 49110 33300 49180
rect 33200 49070 33300 49110
rect 33200 49000 33220 49070
rect 33290 49000 33300 49070
rect 33200 48980 33300 49000
rect 32210 48960 32290 48970
rect 32210 48900 32220 48960
rect 32280 48950 32290 48960
rect 32790 48960 32870 48970
rect 32790 48950 32800 48960
rect 32280 48920 32800 48950
rect 32280 48900 32290 48920
rect 32210 48890 32290 48900
rect 32790 48900 32800 48920
rect 32860 48900 32870 48960
rect 33630 48960 33710 48970
rect 33630 48900 33640 48960
rect 33700 48950 33710 48960
rect 34370 48960 34450 48970
rect 34370 48950 34380 48960
rect 33700 48920 34380 48950
rect 33700 48900 33710 48920
rect 32790 48890 32870 48900
rect 33210 48890 33290 48900
rect 33630 48890 33710 48900
rect 34370 48900 34380 48920
rect 34440 48900 34450 48960
rect 34370 48890 34450 48900
rect 31670 39470 31730 39480
rect 31670 39400 31730 39410
rect 31760 39450 32170 39480
rect 31670 37580 31700 39400
rect 31760 37720 31790 39450
rect 32260 39420 32290 48890
rect 33210 48830 33220 48890
rect 33280 48850 33290 48890
rect 33280 48840 33980 48850
rect 33280 48830 33920 48840
rect 33210 48820 33920 48830
rect 33920 48770 33980 48780
rect 33860 47660 33920 47670
rect 33210 47630 33860 47640
rect 32350 47570 32410 47580
rect 33210 47570 33220 47630
rect 33280 47610 33860 47630
rect 33280 47570 33290 47610
rect 33860 47590 33920 47600
rect 34250 47570 34310 47580
rect 32790 47560 32870 47570
rect 33210 47560 33290 47570
rect 33630 47560 33710 47570
rect 32790 47550 32800 47560
rect 32410 47520 32800 47550
rect 32350 47500 32410 47510
rect 32790 47500 32800 47520
rect 32860 47500 32870 47560
rect 32790 47490 32870 47500
rect 33630 47500 33640 47560
rect 33700 47550 33710 47560
rect 33700 47520 34250 47550
rect 33700 47500 33710 47520
rect 34250 47500 34310 47510
rect 33630 47490 33710 47500
rect 33200 47470 33300 47480
rect 33200 47400 33220 47470
rect 33290 47400 33300 47470
rect 33200 47360 33300 47400
rect 33200 47290 33220 47360
rect 33290 47290 33300 47360
rect 33200 47270 33300 47290
rect 32330 47250 32410 47260
rect 32330 47190 32340 47250
rect 32400 47240 32410 47250
rect 32790 47250 32870 47260
rect 32790 47240 32800 47250
rect 32400 47210 32800 47240
rect 32400 47190 32410 47210
rect 32330 47180 32410 47190
rect 32790 47190 32800 47210
rect 32860 47190 32870 47250
rect 33630 47250 33710 47260
rect 33630 47190 33640 47250
rect 33700 47240 33710 47250
rect 34250 47250 34330 47260
rect 34250 47240 34260 47250
rect 33700 47210 34260 47240
rect 33700 47190 33710 47210
rect 32790 47180 32870 47190
rect 33210 47180 33290 47190
rect 33630 47180 33710 47190
rect 34250 47190 34260 47210
rect 34320 47190 34330 47250
rect 34250 47180 34330 47190
rect 31850 39410 31910 39420
rect 31850 39340 31910 39350
rect 31940 39390 32290 39420
rect 31730 37710 31810 37720
rect 31730 37650 31740 37710
rect 31800 37650 31810 37710
rect 31730 37640 31810 37650
rect 31670 37570 31750 37580
rect 31670 37510 31680 37570
rect 31740 37510 31750 37570
rect 31670 37500 31750 37510
rect 31550 37430 31630 37440
rect 31550 37370 31560 37430
rect 31620 37370 31630 37430
rect 31550 37360 31630 37370
rect 31490 37290 31570 37300
rect 31490 37230 31500 37290
rect 31560 37230 31570 37290
rect 31490 37220 31570 37230
rect 31850 37020 31880 39340
rect 31940 37160 31970 39390
rect 32380 39360 32410 47180
rect 33210 47120 33220 47180
rect 33280 47140 33290 47180
rect 33280 47130 33980 47140
rect 33280 47120 33920 47130
rect 33210 47110 33920 47120
rect 33920 47060 33980 47070
rect 33860 45950 33920 45960
rect 33210 45920 33860 45930
rect 32470 45860 32530 45870
rect 33210 45860 33220 45920
rect 33280 45900 33860 45920
rect 33280 45860 33290 45900
rect 33860 45880 33920 45890
rect 34130 45860 34190 45870
rect 32790 45850 32870 45860
rect 33210 45850 33290 45860
rect 33630 45850 33710 45860
rect 32790 45840 32800 45850
rect 32530 45810 32800 45840
rect 32470 45790 32530 45800
rect 32790 45790 32800 45810
rect 32860 45790 32870 45850
rect 32790 45780 32870 45790
rect 33630 45790 33640 45850
rect 33700 45840 33710 45850
rect 33700 45810 34130 45840
rect 33700 45790 33710 45810
rect 34130 45790 34190 45800
rect 33630 45780 33710 45790
rect 33200 45760 33300 45770
rect 33200 45690 33220 45760
rect 33290 45690 33300 45760
rect 33200 45650 33300 45690
rect 33200 45580 33220 45650
rect 33290 45580 33300 45650
rect 33200 45560 33300 45580
rect 32450 45540 32530 45550
rect 32450 45480 32460 45540
rect 32520 45530 32530 45540
rect 32790 45540 32870 45550
rect 32790 45530 32800 45540
rect 32520 45500 32800 45530
rect 32520 45480 32530 45500
rect 32450 45470 32530 45480
rect 32790 45480 32800 45500
rect 32860 45480 32870 45540
rect 33630 45540 33710 45550
rect 33630 45480 33640 45540
rect 33700 45530 33710 45540
rect 34130 45540 34210 45550
rect 34130 45530 34140 45540
rect 33700 45500 34140 45530
rect 33700 45480 33710 45500
rect 32790 45470 32870 45480
rect 33210 45470 33290 45480
rect 33630 45470 33710 45480
rect 34130 45480 34140 45500
rect 34200 45480 34210 45540
rect 34130 45470 34210 45480
rect 33210 45410 33220 45470
rect 33280 45430 33290 45470
rect 33280 45420 33980 45430
rect 33280 45410 33920 45420
rect 33210 45400 33920 45410
rect 33920 45350 33980 45360
rect 33860 44240 33920 44250
rect 33210 44210 33860 44220
rect 32470 44150 32530 44160
rect 33210 44150 33220 44210
rect 33280 44190 33860 44210
rect 33280 44150 33290 44190
rect 33860 44170 33920 44180
rect 34130 44150 34190 44160
rect 32790 44140 32870 44150
rect 33210 44140 33290 44150
rect 33630 44140 33710 44150
rect 32790 44130 32800 44140
rect 32530 44100 32800 44130
rect 32470 44080 32530 44090
rect 32790 44080 32800 44100
rect 32860 44080 32870 44140
rect 32790 44070 32870 44080
rect 33630 44080 33640 44140
rect 33700 44130 33710 44140
rect 33700 44100 34130 44130
rect 33700 44080 33710 44100
rect 34130 44080 34190 44090
rect 33630 44070 33710 44080
rect 33200 44050 33300 44060
rect 33200 43980 33220 44050
rect 33290 43980 33300 44050
rect 33200 43940 33300 43980
rect 33200 43870 33220 43940
rect 33290 43870 33300 43940
rect 33200 43850 33300 43870
rect 32450 43830 32530 43840
rect 32450 43770 32460 43830
rect 32520 43820 32530 43830
rect 32790 43830 32870 43840
rect 32790 43820 32800 43830
rect 32520 43790 32800 43820
rect 32520 43770 32530 43790
rect 32450 43760 32530 43770
rect 32790 43770 32800 43790
rect 32860 43770 32870 43830
rect 33630 43830 33710 43840
rect 33630 43770 33640 43830
rect 33700 43820 33710 43830
rect 34130 43830 34210 43840
rect 34130 43820 34140 43830
rect 33700 43790 34140 43820
rect 33700 43770 33710 43790
rect 32790 43760 32870 43770
rect 33210 43760 33290 43770
rect 33630 43760 33710 43770
rect 34130 43770 34140 43790
rect 34200 43770 34210 43830
rect 34130 43760 34210 43770
rect 32030 39350 32090 39360
rect 32030 39280 32090 39290
rect 32120 39330 32410 39360
rect 31910 37150 31990 37160
rect 31910 37090 31920 37150
rect 31980 37090 31990 37150
rect 31910 37080 31990 37090
rect 31850 37010 31930 37020
rect 31850 36950 31860 37010
rect 31920 36950 31930 37010
rect 31850 36940 31930 36950
rect 29740 36680 29750 36740
rect 29810 36680 29820 36740
rect 32030 36740 32060 39280
rect 32120 36880 32150 39330
rect 32500 39300 32530 43760
rect 33210 43700 33220 43760
rect 33280 43720 33290 43760
rect 33280 43710 33980 43720
rect 33280 43700 33920 43710
rect 33210 43690 33920 43700
rect 33920 43640 33980 43650
rect 33860 42530 33920 42540
rect 33210 42500 33860 42510
rect 32590 42440 32650 42450
rect 33210 42440 33220 42500
rect 33280 42480 33860 42500
rect 33280 42440 33290 42480
rect 33860 42460 33920 42470
rect 34010 42440 34070 42450
rect 32790 42430 32870 42440
rect 33210 42430 33290 42440
rect 33630 42430 33710 42440
rect 32790 42420 32800 42430
rect 32650 42390 32800 42420
rect 32590 42370 32650 42380
rect 32790 42370 32800 42390
rect 32860 42370 32870 42430
rect 32790 42360 32870 42370
rect 33630 42370 33640 42430
rect 33700 42420 33710 42430
rect 33700 42390 34010 42420
rect 33700 42370 33710 42390
rect 34010 42370 34070 42380
rect 33630 42360 33710 42370
rect 33200 42340 33300 42350
rect 33200 42270 33220 42340
rect 33290 42270 33300 42340
rect 33200 42230 33300 42270
rect 33200 42160 33220 42230
rect 33290 42160 33300 42230
rect 33200 42140 33300 42160
rect 32570 42120 32650 42130
rect 32570 42060 32580 42120
rect 32640 42110 32650 42120
rect 32790 42120 32870 42130
rect 32790 42110 32800 42120
rect 32640 42080 32800 42110
rect 32640 42060 32650 42080
rect 32570 42050 32650 42060
rect 32790 42060 32800 42080
rect 32860 42060 32870 42120
rect 33630 42120 33710 42130
rect 33630 42060 33640 42120
rect 33700 42110 33710 42120
rect 34010 42120 34090 42130
rect 34010 42110 34020 42120
rect 33700 42080 34020 42110
rect 33700 42060 33710 42080
rect 32790 42050 32870 42060
rect 33210 42050 33290 42060
rect 33630 42050 33710 42060
rect 34010 42060 34020 42080
rect 34080 42060 34090 42120
rect 34010 42050 34090 42060
rect 33210 41990 33220 42050
rect 33280 42010 33290 42050
rect 33280 42000 33980 42010
rect 33280 41990 33920 42000
rect 33210 41980 33920 41990
rect 33920 41930 33980 41940
rect 33860 40820 33920 40830
rect 33210 40790 33860 40800
rect 32590 40730 32650 40740
rect 33210 40730 33220 40790
rect 33280 40770 33860 40790
rect 33280 40730 33290 40770
rect 33860 40750 33920 40760
rect 34010 40730 34070 40740
rect 32790 40720 32870 40730
rect 33210 40720 33290 40730
rect 33630 40720 33710 40730
rect 32790 40710 32800 40720
rect 32650 40680 32800 40710
rect 32590 40660 32650 40670
rect 32790 40660 32800 40680
rect 32860 40660 32870 40720
rect 32790 40650 32870 40660
rect 33630 40660 33640 40720
rect 33700 40710 33710 40720
rect 33700 40680 34010 40710
rect 33700 40660 33710 40680
rect 34010 40660 34070 40670
rect 33630 40650 33710 40660
rect 33200 40630 33300 40640
rect 33200 40560 33220 40630
rect 33290 40560 33300 40630
rect 33200 40520 33300 40560
rect 33200 40450 33220 40520
rect 33290 40450 33300 40520
rect 33200 40430 33300 40450
rect 32570 40410 32650 40420
rect 32570 40350 32580 40410
rect 32640 40400 32650 40410
rect 32790 40410 32870 40420
rect 32790 40400 32800 40410
rect 32640 40370 32800 40400
rect 32640 40350 32650 40370
rect 32570 40340 32650 40350
rect 32790 40350 32800 40370
rect 32860 40350 32870 40410
rect 33630 40410 33710 40420
rect 33630 40350 33640 40410
rect 33700 40400 33710 40410
rect 34010 40410 34090 40420
rect 34010 40400 34020 40410
rect 33700 40370 34020 40400
rect 33700 40350 33710 40370
rect 32790 40340 32870 40350
rect 33210 40340 33290 40350
rect 33630 40340 33710 40350
rect 34010 40350 34020 40370
rect 34080 40350 34090 40410
rect 34010 40340 34090 40350
rect 32210 39290 32270 39300
rect 32210 39220 32270 39230
rect 32300 39270 32530 39300
rect 32090 36870 32170 36880
rect 32090 36810 32100 36870
rect 32160 36810 32170 36870
rect 32090 36800 32170 36810
rect 32030 36730 32110 36740
rect 32030 36670 32040 36730
rect 32100 36670 32110 36730
rect 32030 36660 32110 36670
rect 29380 36400 29390 36460
rect 29450 36400 29460 36460
rect 32210 36460 32240 39220
rect 32300 36600 32330 39270
rect 32620 39240 32650 40340
rect 33210 40280 33220 40340
rect 33280 40300 33290 40340
rect 33280 40290 33980 40300
rect 33280 40280 33920 40290
rect 33210 40270 33920 40280
rect 33920 40220 33980 40230
rect 32390 39230 32450 39240
rect 32390 39160 32450 39170
rect 32480 39210 32650 39240
rect 32680 39680 32760 39690
rect 32680 39620 32690 39680
rect 32750 39620 32760 39680
rect 33750 39680 33830 39690
rect 33750 39620 33760 39680
rect 33820 39620 33830 39680
rect 32270 36590 32350 36600
rect 32270 36530 32280 36590
rect 32340 36530 32350 36590
rect 32270 36520 32350 36530
rect 32210 36450 32290 36460
rect 32210 36390 32220 36450
rect 32280 36390 32290 36450
rect 32210 36380 32290 36390
rect 27400 36170 27480 36180
rect 22410 36100 22490 36110
rect 27400 36110 27410 36170
rect 27470 36110 27480 36170
rect 29200 36120 29210 36180
rect 29270 36120 29280 36180
rect 32390 36180 32420 39160
rect 32480 36320 32510 39210
rect 32680 38840 32750 39620
rect 33750 39610 33830 39620
rect 33920 39680 33980 39690
rect 33920 39610 33980 39620
rect 32680 38830 32760 38840
rect 32680 38770 32690 38830
rect 32750 38770 32760 38830
rect 32680 38760 32760 38770
rect 33760 38700 33830 39610
rect 33950 38700 33980 39610
rect 34010 39240 34040 40340
rect 34130 39300 34160 43760
rect 34250 39360 34280 47180
rect 34370 39420 34400 48890
rect 34490 39480 34520 50600
rect 34610 39540 34640 52310
rect 36890 39600 36920 54050
rect 37780 54030 37790 54050
rect 37850 54030 37860 54090
rect 38620 54090 38700 54100
rect 38620 54030 38630 54090
rect 38690 54080 38700 54090
rect 39720 54080 39750 54270
rect 38690 54050 39750 54080
rect 38690 54030 38700 54050
rect 37780 54020 37860 54030
rect 38200 54020 38280 54030
rect 38620 54020 38700 54030
rect 38200 53960 38210 54020
rect 38270 53980 38280 54020
rect 38270 53970 38970 53980
rect 38270 53960 38910 53970
rect 38200 53950 38910 53960
rect 38910 53900 38970 53910
rect 38850 52790 38910 52800
rect 38200 52760 38850 52770
rect 36980 52700 37040 52710
rect 38200 52700 38210 52760
rect 38270 52740 38850 52760
rect 38270 52700 38280 52740
rect 38850 52720 38910 52730
rect 39600 52700 39660 52710
rect 37780 52690 37860 52700
rect 38200 52690 38280 52700
rect 38620 52690 38700 52700
rect 37780 52680 37790 52690
rect 37040 52650 37790 52680
rect 36980 52630 37040 52640
rect 37780 52630 37790 52650
rect 37850 52630 37860 52690
rect 37780 52620 37860 52630
rect 38620 52630 38630 52690
rect 38690 52680 38700 52690
rect 38690 52650 39600 52680
rect 38690 52630 38700 52650
rect 39600 52630 39660 52640
rect 38620 52620 38700 52630
rect 38190 52600 38290 52610
rect 38190 52530 38210 52600
rect 38280 52530 38290 52600
rect 38190 52490 38290 52530
rect 38190 52420 38210 52490
rect 38280 52420 38290 52490
rect 38190 52400 38290 52420
rect 36960 52390 37040 52400
rect 39600 52390 39680 52400
rect 36960 52330 36970 52390
rect 37030 52370 37040 52390
rect 37780 52380 37860 52390
rect 37780 52370 37790 52380
rect 37030 52340 37790 52370
rect 37030 52330 37040 52340
rect 36960 52320 37040 52330
rect 36300 39590 36360 39600
rect 34610 39510 35080 39540
rect 34490 39450 34900 39480
rect 34370 39390 34720 39420
rect 34250 39330 34540 39360
rect 34130 39270 34360 39300
rect 34010 39210 34180 39240
rect 33750 38690 33830 38700
rect 33750 38630 33760 38690
rect 33820 38630 33830 38690
rect 33900 38640 33910 38700
rect 33970 38640 33980 38700
rect 33750 38620 33830 38630
rect 34150 36320 34180 39210
rect 34210 39230 34270 39240
rect 34210 39160 34270 39170
rect 32450 36310 32530 36320
rect 32450 36250 32460 36310
rect 32520 36250 32530 36310
rect 34130 36260 34140 36320
rect 34200 36260 34210 36320
rect 32450 36240 32530 36250
rect 34240 36180 34270 39160
rect 34330 36600 34360 39270
rect 34390 39290 34450 39300
rect 34390 39220 34450 39230
rect 34310 36540 34320 36600
rect 34380 36540 34390 36600
rect 34420 36460 34450 39220
rect 34510 36880 34540 39330
rect 34570 39350 34630 39360
rect 34570 39280 34630 39290
rect 34490 36820 34500 36880
rect 34560 36820 34570 36880
rect 34600 36740 34630 39280
rect 34690 37160 34720 39390
rect 34750 39410 34810 39420
rect 34750 39340 34810 39350
rect 34670 37100 34680 37160
rect 34740 37100 34750 37160
rect 34780 37020 34810 39340
rect 34870 37720 34900 39450
rect 34930 39470 34990 39480
rect 34930 39400 34990 39410
rect 34850 37660 34860 37720
rect 34920 37660 34930 37720
rect 34960 37580 34990 39400
rect 34910 37520 34920 37580
rect 34980 37520 34990 37580
rect 35050 37440 35080 39510
rect 35110 39530 35170 39540
rect 35110 39460 35170 39470
rect 35030 37380 35040 37440
rect 35100 37380 35110 37440
rect 35140 37300 35170 39460
rect 36300 39520 36360 39530
rect 36390 39570 36920 39600
rect 36300 38420 36330 39520
rect 36390 38560 36420 39570
rect 37010 39540 37040 52320
rect 37780 52320 37790 52340
rect 37850 52320 37860 52380
rect 38620 52380 38700 52390
rect 38620 52320 38630 52380
rect 38690 52370 38700 52380
rect 39600 52370 39610 52390
rect 38690 52340 39610 52370
rect 38690 52320 38700 52340
rect 37780 52310 37860 52320
rect 38200 52310 38280 52320
rect 38620 52310 38700 52320
rect 39600 52330 39610 52340
rect 39670 52330 39680 52390
rect 39600 52320 39680 52330
rect 38200 52250 38210 52310
rect 38270 52270 38280 52310
rect 38270 52260 38970 52270
rect 38270 52250 38910 52260
rect 38200 52240 38910 52250
rect 38910 52190 38970 52200
rect 38850 51080 38910 51090
rect 38200 51050 38850 51060
rect 37100 50990 37160 51000
rect 38200 50990 38210 51050
rect 38270 51030 38850 51050
rect 38270 50990 38280 51030
rect 38850 51010 38910 51020
rect 39480 50990 39540 51000
rect 37780 50980 37860 50990
rect 38200 50980 38280 50990
rect 38620 50980 38700 50990
rect 37780 50970 37790 50980
rect 37160 50940 37790 50970
rect 37100 50920 37160 50930
rect 37780 50920 37790 50940
rect 37850 50920 37860 50980
rect 37780 50910 37860 50920
rect 38620 50920 38630 50980
rect 38690 50970 38700 50980
rect 38690 50940 39480 50970
rect 38690 50920 38700 50940
rect 39480 50920 39540 50930
rect 38620 50910 38700 50920
rect 38190 50890 38290 50900
rect 38190 50820 38210 50890
rect 38280 50820 38290 50890
rect 38190 50780 38290 50820
rect 38190 50710 38210 50780
rect 38280 50710 38290 50780
rect 38190 50690 38290 50710
rect 37080 50680 37160 50690
rect 39480 50680 39560 50690
rect 37080 50620 37090 50680
rect 37150 50660 37160 50680
rect 37780 50670 37860 50680
rect 37780 50660 37790 50670
rect 37150 50630 37790 50660
rect 37150 50620 37160 50630
rect 37080 50610 37160 50620
rect 36480 39530 36540 39540
rect 36480 39460 36540 39470
rect 36570 39510 37040 39540
rect 36360 38550 36440 38560
rect 36360 38490 36370 38550
rect 36430 38490 36440 38550
rect 36360 38480 36440 38490
rect 36300 38410 36380 38420
rect 36300 38350 36310 38410
rect 36370 38350 36380 38410
rect 36300 38340 36380 38350
rect 36480 37860 36510 39460
rect 36570 38000 36600 39510
rect 37130 39480 37160 50610
rect 37780 50610 37790 50630
rect 37850 50610 37860 50670
rect 38620 50670 38700 50680
rect 38620 50610 38630 50670
rect 38690 50660 38700 50670
rect 39480 50660 39490 50680
rect 38690 50630 39490 50660
rect 38690 50610 38700 50630
rect 37780 50600 37860 50610
rect 38200 50600 38280 50610
rect 38620 50600 38700 50610
rect 39480 50620 39490 50630
rect 39550 50620 39560 50680
rect 39480 50610 39560 50620
rect 38200 50540 38210 50600
rect 38270 50560 38280 50600
rect 38270 50550 38970 50560
rect 38270 50540 38910 50550
rect 38200 50530 38910 50540
rect 38910 50480 38970 50490
rect 38850 49370 38910 49380
rect 38200 49340 38850 49350
rect 37220 49280 37280 49290
rect 38200 49280 38210 49340
rect 38270 49320 38850 49340
rect 38270 49280 38280 49320
rect 38850 49300 38910 49310
rect 39360 49280 39420 49290
rect 37780 49270 37860 49280
rect 38200 49270 38280 49280
rect 38620 49270 38700 49280
rect 37780 49260 37790 49270
rect 37280 49230 37790 49260
rect 37220 49210 37280 49220
rect 37780 49210 37790 49230
rect 37850 49210 37860 49270
rect 37780 49200 37860 49210
rect 38620 49210 38630 49270
rect 38690 49260 38700 49270
rect 38690 49230 39360 49260
rect 38690 49210 38700 49230
rect 39360 49210 39420 49220
rect 38620 49200 38700 49210
rect 38190 49180 38290 49190
rect 38190 49110 38210 49180
rect 38280 49110 38290 49180
rect 38190 49070 38290 49110
rect 38190 49000 38210 49070
rect 38280 49000 38290 49070
rect 38190 48980 38290 49000
rect 37200 48970 37280 48980
rect 39360 48970 39440 48980
rect 37200 48910 37210 48970
rect 37270 48950 37280 48970
rect 37780 48960 37860 48970
rect 37780 48950 37790 48960
rect 37270 48920 37790 48950
rect 37270 48910 37280 48920
rect 37200 48900 37280 48910
rect 36660 39470 36720 39480
rect 36660 39400 36720 39410
rect 36750 39450 37160 39480
rect 36540 37990 36620 38000
rect 36540 37930 36550 37990
rect 36610 37930 36620 37990
rect 36540 37920 36620 37930
rect 36480 37850 36560 37860
rect 36480 37790 36490 37850
rect 36550 37790 36560 37850
rect 36480 37780 36560 37790
rect 35090 37240 35100 37300
rect 35160 37240 35170 37300
rect 36660 37300 36690 39400
rect 36750 37440 36780 39450
rect 37250 39420 37280 48900
rect 37780 48900 37790 48920
rect 37850 48900 37860 48960
rect 38620 48960 38700 48970
rect 38620 48900 38630 48960
rect 38690 48950 38700 48960
rect 39360 48950 39370 48970
rect 38690 48920 39370 48950
rect 38690 48900 38700 48920
rect 37780 48890 37860 48900
rect 38200 48890 38280 48900
rect 38620 48890 38700 48900
rect 39360 48910 39370 48920
rect 39430 48910 39440 48970
rect 39360 48900 39440 48910
rect 38200 48830 38210 48890
rect 38270 48850 38280 48890
rect 38270 48840 38970 48850
rect 38270 48830 38910 48840
rect 38200 48820 38910 48830
rect 38910 48770 38970 48780
rect 38850 47660 38910 47670
rect 38200 47630 38850 47640
rect 37340 47570 37400 47580
rect 38200 47570 38210 47630
rect 38270 47610 38850 47630
rect 38270 47570 38280 47610
rect 38850 47590 38910 47600
rect 39240 47570 39300 47580
rect 37780 47560 37860 47570
rect 38200 47560 38280 47570
rect 38620 47560 38700 47570
rect 37780 47550 37790 47560
rect 37400 47520 37790 47550
rect 37340 47500 37400 47510
rect 37780 47500 37790 47520
rect 37850 47500 37860 47560
rect 37780 47490 37860 47500
rect 38620 47500 38630 47560
rect 38690 47550 38700 47560
rect 38690 47520 39240 47550
rect 38690 47500 38700 47520
rect 39240 47500 39300 47510
rect 38620 47490 38700 47500
rect 38190 47470 38290 47480
rect 38190 47400 38210 47470
rect 38280 47400 38290 47470
rect 38190 47360 38290 47400
rect 38190 47290 38210 47360
rect 38280 47290 38290 47360
rect 38190 47270 38290 47290
rect 37320 47260 37400 47270
rect 39240 47260 39320 47270
rect 37320 47200 37330 47260
rect 37390 47240 37400 47260
rect 37780 47250 37860 47260
rect 37780 47240 37790 47250
rect 37390 47210 37790 47240
rect 37390 47200 37400 47210
rect 37320 47190 37400 47200
rect 36840 39410 36900 39420
rect 36840 39340 36900 39350
rect 36930 39390 37280 39420
rect 36720 37430 36800 37440
rect 36720 37370 36730 37430
rect 36790 37370 36800 37430
rect 36720 37360 36800 37370
rect 36660 37290 36740 37300
rect 36660 37230 36670 37290
rect 36730 37230 36740 37290
rect 36660 37220 36740 37230
rect 34730 36960 34740 37020
rect 34800 36960 34810 37020
rect 36840 37020 36870 39340
rect 36930 37160 36960 39390
rect 37370 39360 37400 47190
rect 37780 47190 37790 47210
rect 37850 47190 37860 47250
rect 38620 47250 38700 47260
rect 38620 47190 38630 47250
rect 38690 47240 38700 47250
rect 39240 47240 39250 47260
rect 38690 47210 39250 47240
rect 38690 47190 38700 47210
rect 37780 47180 37860 47190
rect 38200 47180 38280 47190
rect 38620 47180 38700 47190
rect 39240 47200 39250 47210
rect 39310 47200 39320 47260
rect 39240 47190 39320 47200
rect 38200 47120 38210 47180
rect 38270 47140 38280 47180
rect 38270 47130 38970 47140
rect 38270 47120 38910 47130
rect 38200 47110 38910 47120
rect 38910 47060 38970 47070
rect 38850 45950 38910 45960
rect 38200 45920 38850 45930
rect 37460 45860 37520 45870
rect 38200 45860 38210 45920
rect 38270 45900 38850 45920
rect 38270 45860 38280 45900
rect 38850 45880 38910 45890
rect 39120 45860 39180 45870
rect 37780 45850 37860 45860
rect 38200 45850 38280 45860
rect 38620 45850 38700 45860
rect 37780 45840 37790 45850
rect 37520 45810 37790 45840
rect 37460 45790 37520 45800
rect 37780 45790 37790 45810
rect 37850 45790 37860 45850
rect 37780 45780 37860 45790
rect 38620 45790 38630 45850
rect 38690 45840 38700 45850
rect 38690 45810 39120 45840
rect 38690 45790 38700 45810
rect 39120 45790 39180 45800
rect 38620 45780 38700 45790
rect 38190 45760 38290 45770
rect 38190 45690 38210 45760
rect 38280 45690 38290 45760
rect 38190 45650 38290 45690
rect 38190 45580 38210 45650
rect 38280 45580 38290 45650
rect 38190 45560 38290 45580
rect 37440 45550 37520 45560
rect 39120 45550 39200 45560
rect 37440 45490 37450 45550
rect 37510 45530 37520 45550
rect 37780 45540 37860 45550
rect 37780 45530 37790 45540
rect 37510 45500 37790 45530
rect 37510 45490 37520 45500
rect 37440 45480 37520 45490
rect 37780 45480 37790 45500
rect 37850 45480 37860 45540
rect 38620 45540 38700 45550
rect 38620 45480 38630 45540
rect 38690 45530 38700 45540
rect 39120 45530 39130 45550
rect 38690 45500 39130 45530
rect 38690 45480 38700 45500
rect 39120 45490 39130 45500
rect 39190 45490 39200 45550
rect 39120 45480 39200 45490
rect 37780 45470 37860 45480
rect 38200 45470 38280 45480
rect 38620 45470 38700 45480
rect 38200 45410 38210 45470
rect 38270 45430 38280 45470
rect 38270 45420 38970 45430
rect 38270 45410 38910 45420
rect 38200 45400 38910 45410
rect 38910 45350 38970 45360
rect 38850 44240 38910 44250
rect 38200 44210 38850 44220
rect 37460 44150 37520 44160
rect 38200 44150 38210 44210
rect 38270 44190 38850 44210
rect 38270 44150 38280 44190
rect 38850 44170 38910 44180
rect 37780 44140 37860 44150
rect 38200 44140 38280 44150
rect 38620 44140 38700 44150
rect 37780 44130 37790 44140
rect 37520 44100 37790 44130
rect 37460 44080 37520 44090
rect 37780 44080 37790 44100
rect 37850 44080 37860 44140
rect 37780 44070 37860 44080
rect 38620 44080 38630 44140
rect 38690 44130 38700 44140
rect 39120 44140 39180 44150
rect 38690 44100 39120 44130
rect 38690 44080 38700 44100
rect 38620 44070 38700 44080
rect 39120 44070 39180 44080
rect 38190 44050 38290 44060
rect 38190 43980 38210 44050
rect 38280 43980 38290 44050
rect 38190 43940 38290 43980
rect 38190 43870 38210 43940
rect 38280 43870 38290 43940
rect 38190 43850 38290 43870
rect 37440 43840 37520 43850
rect 37440 43780 37450 43840
rect 37510 43820 37520 43840
rect 37780 43830 37860 43840
rect 37780 43820 37790 43830
rect 37510 43790 37790 43820
rect 37510 43780 37520 43790
rect 37440 43770 37520 43780
rect 37020 39350 37080 39360
rect 37020 39280 37080 39290
rect 37110 39330 37400 39360
rect 36900 37150 36980 37160
rect 36900 37090 36910 37150
rect 36970 37090 36980 37150
rect 36900 37080 36980 37090
rect 36840 37010 36920 37020
rect 36840 36950 36850 37010
rect 36910 36950 36920 37010
rect 36840 36940 36920 36950
rect 34550 36680 34560 36740
rect 34620 36680 34630 36740
rect 37020 36740 37050 39280
rect 37110 36880 37140 39330
rect 37490 39300 37520 43770
rect 37780 43770 37790 43790
rect 37850 43770 37860 43830
rect 38620 43830 38700 43840
rect 38620 43770 38630 43830
rect 38690 43820 38700 43830
rect 39120 43830 39200 43840
rect 39120 43820 39130 43830
rect 38690 43790 39130 43820
rect 38690 43770 38700 43790
rect 37780 43760 37860 43770
rect 38200 43760 38280 43770
rect 38620 43760 38700 43770
rect 39120 43770 39130 43790
rect 39190 43770 39200 43830
rect 39120 43760 39200 43770
rect 38200 43700 38210 43760
rect 38270 43720 38280 43760
rect 38270 43710 38970 43720
rect 38270 43700 38910 43710
rect 38200 43690 38910 43700
rect 38910 43640 38970 43650
rect 38850 42530 38910 42540
rect 38200 42500 38850 42510
rect 37580 42440 37640 42450
rect 38200 42440 38210 42500
rect 38270 42480 38850 42500
rect 38270 42440 38280 42480
rect 38850 42460 38910 42470
rect 37780 42430 37860 42440
rect 38200 42430 38280 42440
rect 38620 42430 38700 42440
rect 37780 42420 37790 42430
rect 37640 42390 37790 42420
rect 37580 42370 37640 42380
rect 37780 42370 37790 42390
rect 37850 42370 37860 42430
rect 37780 42360 37860 42370
rect 38620 42370 38630 42430
rect 38690 42420 38700 42430
rect 39000 42430 39060 42440
rect 38690 42390 39000 42420
rect 38690 42370 38700 42390
rect 38620 42360 38700 42370
rect 39000 42360 39060 42370
rect 38190 42340 38290 42350
rect 38190 42270 38210 42340
rect 38280 42270 38290 42340
rect 38190 42230 38290 42270
rect 38190 42160 38210 42230
rect 38280 42160 38290 42230
rect 38190 42140 38290 42160
rect 37560 42130 37640 42140
rect 37560 42070 37570 42130
rect 37630 42110 37640 42130
rect 37780 42120 37860 42130
rect 37780 42110 37790 42120
rect 37630 42080 37790 42110
rect 37630 42070 37640 42080
rect 37560 42060 37640 42070
rect 37780 42060 37790 42080
rect 37850 42060 37860 42120
rect 38620 42120 38700 42130
rect 38620 42060 38630 42120
rect 38690 42110 38700 42120
rect 39000 42120 39080 42130
rect 39000 42110 39010 42120
rect 38690 42080 39010 42110
rect 38690 42060 38700 42080
rect 37780 42050 37860 42060
rect 38200 42050 38280 42060
rect 38620 42050 38700 42060
rect 39000 42060 39010 42080
rect 39070 42060 39080 42120
rect 39000 42050 39080 42060
rect 38200 41990 38210 42050
rect 38270 42010 38280 42050
rect 38270 42000 38970 42010
rect 38270 41990 38910 42000
rect 38200 41980 38910 41990
rect 38910 41930 38970 41940
rect 38850 40820 38910 40830
rect 38200 40790 38850 40800
rect 37580 40730 37640 40740
rect 38200 40730 38210 40790
rect 38270 40770 38850 40790
rect 38270 40730 38280 40770
rect 38850 40750 38910 40760
rect 39000 40730 39060 40740
rect 37780 40720 37860 40730
rect 38200 40720 38280 40730
rect 38620 40720 38700 40730
rect 37780 40710 37790 40720
rect 37640 40680 37790 40710
rect 37580 40660 37640 40670
rect 37780 40660 37790 40680
rect 37850 40660 37860 40720
rect 37780 40650 37860 40660
rect 38620 40660 38630 40720
rect 38690 40710 38700 40720
rect 38690 40680 39000 40710
rect 38690 40660 38700 40680
rect 39000 40660 39060 40670
rect 38620 40650 38700 40660
rect 38190 40630 38290 40640
rect 38190 40560 38210 40630
rect 38280 40560 38290 40630
rect 38190 40520 38290 40560
rect 38190 40450 38210 40520
rect 38280 40450 38290 40520
rect 38190 40430 38290 40450
rect 37560 40420 37640 40430
rect 39000 40420 39080 40430
rect 37560 40360 37570 40420
rect 37630 40400 37640 40420
rect 37780 40410 37860 40420
rect 37780 40400 37790 40410
rect 37630 40370 37790 40400
rect 37630 40360 37640 40370
rect 37560 40350 37640 40360
rect 37200 39290 37260 39300
rect 37200 39220 37260 39230
rect 37290 39270 37520 39300
rect 37080 36870 37160 36880
rect 37080 36810 37090 36870
rect 37150 36810 37160 36870
rect 37080 36800 37160 36810
rect 37020 36730 37100 36740
rect 37020 36670 37030 36730
rect 37090 36670 37100 36730
rect 37020 36660 37100 36670
rect 34370 36400 34380 36460
rect 34440 36400 34450 36460
rect 37200 36460 37230 39220
rect 37290 36600 37320 39270
rect 37610 39240 37640 40350
rect 37780 40350 37790 40370
rect 37850 40350 37860 40410
rect 38620 40410 38700 40420
rect 38620 40350 38630 40410
rect 38690 40400 38700 40410
rect 39000 40400 39010 40420
rect 38690 40370 39010 40400
rect 38690 40350 38700 40370
rect 39000 40360 39010 40370
rect 39070 40360 39080 40420
rect 39000 40350 39080 40360
rect 37780 40340 37860 40350
rect 38200 40340 38280 40350
rect 38620 40340 38700 40350
rect 38200 40280 38210 40340
rect 38270 40300 38280 40340
rect 38270 40290 38970 40300
rect 38270 40280 38910 40290
rect 38200 40270 38910 40280
rect 38910 40220 38970 40230
rect 39000 40210 39080 40220
rect 39000 40150 39010 40210
rect 39070 40150 39080 40210
rect 39000 40140 39080 40150
rect 37380 39230 37440 39240
rect 37380 39160 37440 39170
rect 37470 39210 37640 39240
rect 37670 39680 37750 39690
rect 37670 39620 37680 39680
rect 37740 39620 37750 39680
rect 38740 39680 38820 39690
rect 38740 39620 38750 39680
rect 38810 39620 38820 39680
rect 37260 36590 37340 36600
rect 37260 36530 37270 36590
rect 37330 36530 37340 36590
rect 37260 36520 37340 36530
rect 37200 36450 37280 36460
rect 37200 36390 37210 36450
rect 37270 36390 37280 36450
rect 37200 36380 37280 36390
rect 32390 36170 32470 36180
rect 27400 36100 27480 36110
rect 32390 36110 32400 36170
rect 32460 36110 32470 36170
rect 34190 36120 34200 36180
rect 34260 36120 34270 36180
rect 37380 36180 37410 39160
rect 37470 36320 37500 39210
rect 37670 38840 37740 39620
rect 38740 39610 38820 39620
rect 38910 39680 38970 39690
rect 38910 39610 38970 39620
rect 37670 38830 37750 38840
rect 37670 38770 37680 38830
rect 37740 38770 37750 38830
rect 37670 38760 37750 38770
rect 38750 38700 38820 39610
rect 38940 38700 38970 39610
rect 39000 39240 39030 40140
rect 39120 39300 39150 43760
rect 39240 39360 39270 47190
rect 39360 39420 39390 48900
rect 39480 39480 39510 50610
rect 39600 39540 39630 52320
rect 39720 39600 39750 54050
rect 41880 54080 41910 54270
rect 43180 54240 43200 54310
rect 43270 54240 43280 54310
rect 44800 54300 44830 54440
rect 46960 54410 47020 54420
rect 48180 54410 48190 54470
rect 48250 54450 48830 54470
rect 48250 54410 48260 54450
rect 53820 54500 53880 54510
rect 48830 54430 48890 54440
rect 53170 54470 53820 54480
rect 49580 54410 49640 54420
rect 47760 54400 47840 54410
rect 48180 54400 48260 54410
rect 48600 54400 48680 54410
rect 47760 54390 47770 54400
rect 47020 54360 47770 54390
rect 46960 54340 47020 54350
rect 47760 54340 47770 54360
rect 47830 54340 47840 54400
rect 47760 54330 47840 54340
rect 48600 54340 48610 54400
rect 48670 54390 48680 54400
rect 48670 54360 49580 54390
rect 48670 54340 48680 54360
rect 49580 54340 49640 54350
rect 52190 54410 52250 54420
rect 53170 54410 53180 54470
rect 53240 54450 53820 54470
rect 53240 54410 53250 54450
rect 58810 54500 58870 54510
rect 53820 54430 53880 54440
rect 58160 54470 58810 54480
rect 54330 54410 54390 54420
rect 52750 54400 52830 54410
rect 53170 54400 53250 54410
rect 53590 54400 53670 54410
rect 52750 54390 52760 54400
rect 52250 54360 52760 54390
rect 52190 54340 52250 54350
rect 52750 54340 52760 54360
rect 52820 54340 52830 54400
rect 48600 54330 48680 54340
rect 52750 54330 52830 54340
rect 53590 54340 53600 54400
rect 53660 54390 53670 54400
rect 53660 54360 54330 54390
rect 53660 54340 53670 54360
rect 54330 54340 54390 54350
rect 57180 54410 57240 54420
rect 58160 54410 58170 54470
rect 58230 54450 58810 54470
rect 58230 54410 58240 54450
rect 63800 54500 63860 54510
rect 58810 54430 58870 54440
rect 63150 54470 63800 54480
rect 59320 54410 59380 54420
rect 57740 54400 57820 54410
rect 58160 54400 58240 54410
rect 58580 54400 58660 54410
rect 57740 54390 57750 54400
rect 57240 54360 57750 54390
rect 57180 54340 57240 54350
rect 57740 54340 57750 54360
rect 57810 54340 57820 54400
rect 53590 54330 53670 54340
rect 57740 54330 57820 54340
rect 58580 54340 58590 54400
rect 58650 54390 58660 54400
rect 58650 54360 59320 54390
rect 58650 54340 58660 54360
rect 59320 54340 59380 54350
rect 62410 54410 62470 54420
rect 63150 54410 63160 54470
rect 63220 54450 63800 54470
rect 63220 54410 63230 54450
rect 68790 54500 68850 54510
rect 63800 54430 63860 54440
rect 68140 54470 68790 54480
rect 64070 54410 64130 54420
rect 62730 54400 62810 54410
rect 63150 54400 63230 54410
rect 63570 54400 63650 54410
rect 62730 54390 62740 54400
rect 62470 54360 62740 54390
rect 62410 54340 62470 54350
rect 62730 54340 62740 54360
rect 62800 54340 62810 54400
rect 58580 54330 58660 54340
rect 62730 54330 62810 54340
rect 63570 54340 63580 54400
rect 63640 54390 63650 54400
rect 63640 54360 64070 54390
rect 63640 54340 63650 54360
rect 64070 54340 64130 54350
rect 67400 54410 67460 54420
rect 68140 54410 68150 54470
rect 68210 54450 68790 54470
rect 68210 54410 68220 54450
rect 73780 54500 73840 54510
rect 68790 54430 68850 54440
rect 73130 54470 73780 54480
rect 69060 54410 69120 54420
rect 67720 54400 67800 54410
rect 68140 54400 68220 54410
rect 68560 54400 68640 54410
rect 67720 54390 67730 54400
rect 67460 54360 67730 54390
rect 67400 54340 67460 54350
rect 67720 54340 67730 54360
rect 67790 54340 67800 54400
rect 63570 54330 63650 54340
rect 67720 54330 67800 54340
rect 68560 54340 68570 54400
rect 68630 54390 68640 54400
rect 68630 54360 69060 54390
rect 68630 54340 68640 54360
rect 69060 54340 69120 54350
rect 72510 54410 72570 54420
rect 73130 54410 73140 54470
rect 73200 54450 73780 54470
rect 73200 54410 73210 54450
rect 78770 54500 78830 54510
rect 73780 54430 73840 54440
rect 78120 54470 78770 54480
rect 73930 54410 73990 54420
rect 72710 54400 72790 54410
rect 73130 54400 73210 54410
rect 73550 54400 73630 54410
rect 72710 54390 72720 54400
rect 72570 54360 72720 54390
rect 72510 54340 72570 54350
rect 72710 54340 72720 54360
rect 72780 54340 72790 54400
rect 68560 54330 68640 54340
rect 72710 54330 72790 54340
rect 73550 54340 73560 54400
rect 73620 54390 73630 54400
rect 73620 54360 73930 54390
rect 73620 54340 73630 54360
rect 73930 54340 73990 54350
rect 77500 54410 77560 54420
rect 78120 54410 78130 54470
rect 78190 54450 78770 54470
rect 78190 54410 78200 54450
rect 78770 54430 78830 54440
rect 78920 54410 78980 54420
rect 77700 54400 77780 54410
rect 78120 54400 78200 54410
rect 78540 54400 78620 54410
rect 77700 54390 77710 54400
rect 77560 54360 77710 54390
rect 77500 54340 77560 54350
rect 77700 54340 77710 54360
rect 77770 54340 77780 54400
rect 73550 54330 73630 54340
rect 77700 54330 77780 54340
rect 78540 54340 78550 54400
rect 78610 54390 78620 54400
rect 78610 54360 78920 54390
rect 78610 54340 78620 54360
rect 78920 54340 78980 54350
rect 78540 54330 78620 54340
rect 43180 54200 43280 54240
rect 43180 54130 43200 54200
rect 43270 54130 43280 54200
rect 43180 54110 43280 54130
rect 44710 54270 44830 54300
rect 48170 54310 48270 54320
rect 42770 54090 42850 54100
rect 42770 54080 42780 54090
rect 41880 54050 42780 54080
rect 41880 39600 41910 54050
rect 42770 54030 42780 54050
rect 42840 54030 42850 54090
rect 43610 54090 43690 54100
rect 43610 54030 43620 54090
rect 43680 54080 43690 54090
rect 44710 54080 44740 54270
rect 48170 54240 48190 54310
rect 48260 54240 48270 54310
rect 48170 54200 48270 54240
rect 48170 54130 48190 54200
rect 48260 54130 48270 54200
rect 48170 54110 48270 54130
rect 53160 54310 53260 54320
rect 53160 54240 53180 54310
rect 53250 54240 53260 54310
rect 53160 54200 53260 54240
rect 53160 54130 53180 54200
rect 53250 54130 53260 54200
rect 53160 54110 53260 54130
rect 58150 54310 58250 54320
rect 58150 54240 58170 54310
rect 58240 54240 58250 54310
rect 58150 54200 58250 54240
rect 58150 54130 58170 54200
rect 58240 54130 58250 54200
rect 58150 54110 58250 54130
rect 63140 54310 63240 54320
rect 63140 54240 63160 54310
rect 63230 54240 63240 54310
rect 63140 54200 63240 54240
rect 63140 54130 63160 54200
rect 63230 54130 63240 54200
rect 63140 54110 63240 54130
rect 68130 54310 68230 54320
rect 68130 54240 68150 54310
rect 68220 54240 68230 54310
rect 68130 54200 68230 54240
rect 68130 54130 68150 54200
rect 68220 54130 68230 54200
rect 68130 54110 68230 54130
rect 73120 54310 73220 54320
rect 73120 54240 73140 54310
rect 73210 54240 73220 54310
rect 73120 54200 73220 54240
rect 73120 54130 73140 54200
rect 73210 54130 73220 54200
rect 73120 54110 73220 54130
rect 78110 54310 78210 54320
rect 78110 54240 78130 54310
rect 78200 54240 78210 54310
rect 78110 54200 78210 54240
rect 78110 54130 78130 54200
rect 78200 54130 78210 54200
rect 78110 54110 78210 54130
rect 43680 54050 44740 54080
rect 43680 54030 43690 54050
rect 42770 54020 42850 54030
rect 43190 54020 43270 54030
rect 43610 54020 43690 54030
rect 43190 53960 43200 54020
rect 43260 53980 43270 54020
rect 43260 53970 43960 53980
rect 43260 53960 43900 53970
rect 43190 53950 43900 53960
rect 43900 53900 43960 53910
rect 43840 52790 43900 52800
rect 43190 52760 43840 52770
rect 41970 52700 42030 52710
rect 43190 52700 43200 52760
rect 43260 52740 43840 52760
rect 43260 52700 43270 52740
rect 43840 52720 43900 52730
rect 44590 52700 44650 52710
rect 42770 52690 42850 52700
rect 43190 52690 43270 52700
rect 43610 52690 43690 52700
rect 42770 52680 42780 52690
rect 42030 52650 42780 52680
rect 41970 52630 42030 52640
rect 42770 52630 42780 52650
rect 42840 52630 42850 52690
rect 42770 52620 42850 52630
rect 43610 52630 43620 52690
rect 43680 52680 43690 52690
rect 43680 52650 44590 52680
rect 43680 52630 43690 52650
rect 44590 52630 44650 52640
rect 43610 52620 43690 52630
rect 43180 52600 43280 52610
rect 43180 52530 43200 52600
rect 43270 52530 43280 52600
rect 43180 52490 43280 52530
rect 43180 52420 43200 52490
rect 43270 52420 43280 52490
rect 43180 52400 43280 52420
rect 41950 52390 42030 52400
rect 44590 52390 44670 52400
rect 41950 52330 41960 52390
rect 42020 52370 42030 52390
rect 42770 52380 42850 52390
rect 42770 52370 42780 52380
rect 42020 52340 42780 52370
rect 42020 52330 42030 52340
rect 41950 52320 42030 52330
rect 39720 39570 40250 39600
rect 39600 39510 40070 39540
rect 39480 39450 39890 39480
rect 39360 39390 39710 39420
rect 39240 39330 39530 39360
rect 39120 39270 39350 39300
rect 39000 39210 39170 39240
rect 38740 38690 38820 38700
rect 38740 38630 38750 38690
rect 38810 38630 38820 38690
rect 38890 38640 38900 38700
rect 38960 38640 38970 38700
rect 38740 38620 38820 38630
rect 39140 36320 39170 39210
rect 39200 39230 39260 39240
rect 39200 39160 39260 39170
rect 37440 36310 37520 36320
rect 37440 36250 37450 36310
rect 37510 36250 37520 36310
rect 39120 36260 39130 36320
rect 39190 36260 39200 36320
rect 37440 36240 37520 36250
rect 39230 36180 39260 39160
rect 39320 36600 39350 39270
rect 39380 39290 39440 39300
rect 39380 39220 39440 39230
rect 39300 36540 39310 36600
rect 39370 36540 39380 36600
rect 39410 36460 39440 39220
rect 39500 36880 39530 39330
rect 39560 39350 39620 39360
rect 39560 39280 39620 39290
rect 39480 36820 39490 36880
rect 39550 36820 39560 36880
rect 39590 36740 39620 39280
rect 39680 37160 39710 39390
rect 39740 39410 39800 39420
rect 39740 39340 39800 39350
rect 39660 37100 39670 37160
rect 39730 37100 39740 37160
rect 39770 37020 39800 39340
rect 39860 37440 39890 39450
rect 39920 39470 39980 39480
rect 39920 39400 39980 39410
rect 39840 37380 39850 37440
rect 39910 37380 39920 37440
rect 39950 37300 39980 39400
rect 40040 38000 40070 39510
rect 40100 39530 40160 39540
rect 40100 39460 40160 39470
rect 40020 37940 40030 38000
rect 40090 37940 40100 38000
rect 40130 37860 40160 39460
rect 40220 38560 40250 39570
rect 40280 39590 40340 39600
rect 40280 39520 40340 39530
rect 40190 38500 40200 38560
rect 40260 38500 40270 38560
rect 40310 38420 40340 39520
rect 40260 38360 40270 38420
rect 40330 38360 40340 38420
rect 41290 39590 41350 39600
rect 41290 39520 41350 39530
rect 41380 39570 41910 39600
rect 40080 37800 40090 37860
rect 40150 37800 40160 37860
rect 41290 37860 41320 39520
rect 41380 38000 41410 39570
rect 42000 39540 42030 52320
rect 42770 52320 42780 52340
rect 42840 52320 42850 52380
rect 43610 52380 43690 52390
rect 43610 52320 43620 52380
rect 43680 52370 43690 52380
rect 44590 52370 44600 52390
rect 43680 52340 44600 52370
rect 43680 52320 43690 52340
rect 42770 52310 42850 52320
rect 43190 52310 43270 52320
rect 43610 52310 43690 52320
rect 44590 52330 44600 52340
rect 44660 52330 44670 52390
rect 44590 52320 44670 52330
rect 43190 52250 43200 52310
rect 43260 52270 43270 52310
rect 43260 52260 43960 52270
rect 43260 52250 43900 52260
rect 43190 52240 43900 52250
rect 43900 52190 43960 52200
rect 43840 51080 43900 51090
rect 43190 51050 43840 51060
rect 42090 50990 42150 51000
rect 43190 50990 43200 51050
rect 43260 51030 43840 51050
rect 43260 50990 43270 51030
rect 43840 51010 43900 51020
rect 44470 50990 44530 51000
rect 42770 50980 42850 50990
rect 43190 50980 43270 50990
rect 43610 50980 43690 50990
rect 42770 50970 42780 50980
rect 42150 50940 42780 50970
rect 42090 50920 42150 50930
rect 42770 50920 42780 50940
rect 42840 50920 42850 50980
rect 42770 50910 42850 50920
rect 43610 50920 43620 50980
rect 43680 50970 43690 50980
rect 43680 50940 44470 50970
rect 43680 50920 43690 50940
rect 44470 50920 44530 50930
rect 43610 50910 43690 50920
rect 43180 50890 43280 50900
rect 43180 50820 43200 50890
rect 43270 50820 43280 50890
rect 43180 50780 43280 50820
rect 43180 50710 43200 50780
rect 43270 50710 43280 50780
rect 43180 50690 43280 50710
rect 42070 50680 42150 50690
rect 44470 50680 44550 50690
rect 42070 50620 42080 50680
rect 42140 50660 42150 50680
rect 42770 50670 42850 50680
rect 42770 50660 42780 50670
rect 42140 50630 42780 50660
rect 42140 50620 42150 50630
rect 42070 50610 42150 50620
rect 41470 39530 41530 39540
rect 41470 39460 41530 39470
rect 41560 39510 42030 39540
rect 41470 38140 41500 39460
rect 41560 38280 41590 39510
rect 42120 39480 42150 50610
rect 42770 50610 42780 50630
rect 42840 50610 42850 50670
rect 43610 50670 43690 50680
rect 43610 50610 43620 50670
rect 43680 50660 43690 50670
rect 44470 50660 44480 50680
rect 43680 50630 44480 50660
rect 43680 50610 43690 50630
rect 42770 50600 42850 50610
rect 43190 50600 43270 50610
rect 43610 50600 43690 50610
rect 44470 50620 44480 50630
rect 44540 50620 44550 50680
rect 44470 50610 44550 50620
rect 43190 50540 43200 50600
rect 43260 50560 43270 50600
rect 43260 50550 43960 50560
rect 43260 50540 43900 50550
rect 43190 50530 43900 50540
rect 43900 50480 43960 50490
rect 43840 49370 43900 49380
rect 43190 49340 43840 49350
rect 42210 49280 42270 49290
rect 43190 49280 43200 49340
rect 43260 49320 43840 49340
rect 43260 49280 43270 49320
rect 43840 49300 43900 49310
rect 44350 49280 44410 49290
rect 42770 49270 42850 49280
rect 43190 49270 43270 49280
rect 43610 49270 43690 49280
rect 42770 49260 42780 49270
rect 42270 49230 42780 49260
rect 42210 49210 42270 49220
rect 42770 49210 42780 49230
rect 42840 49210 42850 49270
rect 42770 49200 42850 49210
rect 43610 49210 43620 49270
rect 43680 49260 43690 49270
rect 43680 49230 44350 49260
rect 43680 49210 43690 49230
rect 44350 49210 44410 49220
rect 43610 49200 43690 49210
rect 43180 49180 43280 49190
rect 43180 49110 43200 49180
rect 43270 49110 43280 49180
rect 43180 49070 43280 49110
rect 43180 49000 43200 49070
rect 43270 49000 43280 49070
rect 43180 48980 43280 49000
rect 42190 48970 42270 48980
rect 44350 48970 44430 48980
rect 42190 48910 42200 48970
rect 42260 48950 42270 48970
rect 42770 48960 42850 48970
rect 42770 48950 42780 48960
rect 42260 48920 42780 48950
rect 42260 48910 42270 48920
rect 42190 48900 42270 48910
rect 41650 39470 41710 39480
rect 41650 39400 41710 39410
rect 41740 39450 42150 39480
rect 41530 38270 41610 38280
rect 41530 38210 41540 38270
rect 41600 38210 41610 38270
rect 41530 38200 41610 38210
rect 41440 38130 41520 38140
rect 41440 38070 41450 38130
rect 41510 38070 41520 38130
rect 41440 38060 41520 38070
rect 41350 37990 41430 38000
rect 41350 37930 41360 37990
rect 41420 37930 41430 37990
rect 41350 37920 41430 37930
rect 41290 37850 41370 37860
rect 41290 37790 41300 37850
rect 41360 37790 41370 37850
rect 41290 37780 41370 37790
rect 39900 37240 39910 37300
rect 39970 37240 39980 37300
rect 41650 37300 41680 39400
rect 41740 37440 41770 39450
rect 42240 39420 42270 48900
rect 42770 48900 42780 48920
rect 42840 48900 42850 48960
rect 43610 48960 43690 48970
rect 43610 48900 43620 48960
rect 43680 48950 43690 48960
rect 44350 48950 44360 48970
rect 43680 48920 44360 48950
rect 43680 48900 43690 48920
rect 42770 48890 42850 48900
rect 43190 48890 43270 48900
rect 43610 48890 43690 48900
rect 44350 48910 44360 48920
rect 44420 48910 44430 48970
rect 44350 48900 44430 48910
rect 43190 48830 43200 48890
rect 43260 48850 43270 48890
rect 43260 48840 43960 48850
rect 43260 48830 43900 48840
rect 43190 48820 43900 48830
rect 43900 48770 43960 48780
rect 43840 47660 43900 47670
rect 43190 47630 43840 47640
rect 42330 47570 42390 47580
rect 43190 47570 43200 47630
rect 43260 47610 43840 47630
rect 43260 47570 43270 47610
rect 43840 47590 43900 47600
rect 44230 47570 44290 47580
rect 42770 47560 42850 47570
rect 43190 47560 43270 47570
rect 43610 47560 43690 47570
rect 42770 47550 42780 47560
rect 42390 47520 42780 47550
rect 42330 47500 42390 47510
rect 42770 47500 42780 47520
rect 42840 47500 42850 47560
rect 42770 47490 42850 47500
rect 43610 47500 43620 47560
rect 43680 47550 43690 47560
rect 43680 47520 44230 47550
rect 43680 47500 43690 47520
rect 44230 47500 44290 47510
rect 43610 47490 43690 47500
rect 43180 47470 43280 47480
rect 43180 47400 43200 47470
rect 43270 47400 43280 47470
rect 43180 47360 43280 47400
rect 43180 47290 43200 47360
rect 43270 47290 43280 47360
rect 43180 47270 43280 47290
rect 42310 47260 42390 47270
rect 44230 47260 44310 47270
rect 42310 47200 42320 47260
rect 42380 47240 42390 47260
rect 42770 47250 42850 47260
rect 42770 47240 42780 47250
rect 42380 47210 42780 47240
rect 42380 47200 42390 47210
rect 42310 47190 42390 47200
rect 41830 39410 41890 39420
rect 41830 39340 41890 39350
rect 41920 39390 42270 39420
rect 41710 37430 41790 37440
rect 41710 37370 41720 37430
rect 41780 37370 41790 37430
rect 41710 37360 41790 37370
rect 41650 37290 41730 37300
rect 41650 37230 41660 37290
rect 41720 37230 41730 37290
rect 41650 37220 41730 37230
rect 39720 36960 39730 37020
rect 39790 36960 39800 37020
rect 41830 37020 41860 39340
rect 41920 37160 41950 39390
rect 42360 39360 42390 47190
rect 42770 47190 42780 47210
rect 42840 47190 42850 47250
rect 43610 47250 43690 47260
rect 43610 47190 43620 47250
rect 43680 47240 43690 47250
rect 44230 47240 44240 47260
rect 43680 47210 44240 47240
rect 43680 47190 43690 47210
rect 42770 47180 42850 47190
rect 43190 47180 43270 47190
rect 43610 47180 43690 47190
rect 44230 47200 44240 47210
rect 44300 47200 44310 47260
rect 44230 47190 44310 47200
rect 43190 47120 43200 47180
rect 43260 47140 43270 47180
rect 43260 47130 43960 47140
rect 43260 47120 43900 47130
rect 43190 47110 43900 47120
rect 43900 47060 43960 47070
rect 43840 45950 43900 45960
rect 43190 45920 43840 45930
rect 42450 45860 42510 45870
rect 43190 45860 43200 45920
rect 43260 45900 43840 45920
rect 43260 45860 43270 45900
rect 43840 45880 43900 45890
rect 44110 45860 44170 45870
rect 42770 45850 42850 45860
rect 43190 45850 43270 45860
rect 43610 45850 43690 45860
rect 42770 45840 42780 45850
rect 42510 45810 42780 45840
rect 42450 45790 42510 45800
rect 42770 45790 42780 45810
rect 42840 45790 42850 45850
rect 42770 45780 42850 45790
rect 43610 45790 43620 45850
rect 43680 45840 43690 45850
rect 43680 45810 44110 45840
rect 43680 45790 43690 45810
rect 44110 45790 44170 45800
rect 43610 45780 43690 45790
rect 43180 45760 43280 45770
rect 43180 45690 43200 45760
rect 43270 45690 43280 45760
rect 43180 45650 43280 45690
rect 43180 45580 43200 45650
rect 43270 45580 43280 45650
rect 43180 45560 43280 45580
rect 42430 45550 42510 45560
rect 44110 45550 44190 45560
rect 42430 45490 42440 45550
rect 42500 45530 42510 45550
rect 42770 45540 42850 45550
rect 42770 45530 42780 45540
rect 42500 45500 42780 45530
rect 42500 45490 42510 45500
rect 42430 45480 42510 45490
rect 42770 45480 42780 45500
rect 42840 45480 42850 45540
rect 43610 45540 43690 45550
rect 43610 45480 43620 45540
rect 43680 45530 43690 45540
rect 44110 45530 44120 45550
rect 43680 45500 44120 45530
rect 43680 45480 43690 45500
rect 44110 45490 44120 45500
rect 44180 45490 44190 45550
rect 44110 45480 44190 45490
rect 42770 45470 42850 45480
rect 43190 45470 43270 45480
rect 43610 45470 43690 45480
rect 43190 45410 43200 45470
rect 43260 45430 43270 45470
rect 43260 45420 43960 45430
rect 43260 45410 43900 45420
rect 43190 45400 43900 45410
rect 43900 45350 43960 45360
rect 43840 44240 43900 44250
rect 43190 44210 43840 44220
rect 42450 44150 42510 44160
rect 43190 44150 43200 44210
rect 43260 44190 43840 44210
rect 43260 44150 43270 44190
rect 43840 44170 43900 44180
rect 42770 44140 42850 44150
rect 43190 44140 43270 44150
rect 43610 44140 43690 44150
rect 42770 44130 42780 44140
rect 42510 44100 42780 44130
rect 42450 44080 42510 44090
rect 42770 44080 42780 44100
rect 42840 44080 42850 44140
rect 42770 44070 42850 44080
rect 43610 44080 43620 44140
rect 43680 44130 43690 44140
rect 44110 44140 44170 44150
rect 43680 44100 44110 44130
rect 43680 44080 43690 44100
rect 43610 44070 43690 44080
rect 44110 44070 44170 44080
rect 43180 44050 43280 44060
rect 43180 43980 43200 44050
rect 43270 43980 43280 44050
rect 43180 43940 43280 43980
rect 43180 43870 43200 43940
rect 43270 43870 43280 43940
rect 43180 43850 43280 43870
rect 42430 43840 42510 43850
rect 42430 43780 42440 43840
rect 42500 43820 42510 43840
rect 42770 43830 42850 43840
rect 42770 43820 42780 43830
rect 42500 43790 42780 43820
rect 42500 43780 42510 43790
rect 42430 43770 42510 43780
rect 42010 39350 42070 39360
rect 42010 39280 42070 39290
rect 42100 39330 42390 39360
rect 41890 37150 41970 37160
rect 41890 37090 41900 37150
rect 41960 37090 41970 37150
rect 41890 37080 41970 37090
rect 41830 37010 41910 37020
rect 41830 36950 41840 37010
rect 41900 36950 41910 37010
rect 41830 36940 41910 36950
rect 39540 36680 39550 36740
rect 39610 36680 39620 36740
rect 42010 36740 42040 39280
rect 42100 36880 42130 39330
rect 42480 39300 42510 43770
rect 42770 43770 42780 43790
rect 42840 43770 42850 43830
rect 43610 43830 43690 43840
rect 43610 43770 43620 43830
rect 43680 43820 43690 43830
rect 44110 43830 44190 43840
rect 44110 43820 44120 43830
rect 43680 43790 44120 43820
rect 43680 43770 43690 43790
rect 42770 43760 42850 43770
rect 43190 43760 43270 43770
rect 43610 43760 43690 43770
rect 44110 43770 44120 43790
rect 44180 43770 44190 43830
rect 44110 43760 44190 43770
rect 43190 43700 43200 43760
rect 43260 43720 43270 43760
rect 43260 43710 43960 43720
rect 43260 43700 43900 43710
rect 43190 43690 43900 43700
rect 43900 43640 43960 43650
rect 43840 42530 43900 42540
rect 43190 42500 43840 42510
rect 42570 42440 42630 42450
rect 43190 42440 43200 42500
rect 43260 42480 43840 42500
rect 43260 42440 43270 42480
rect 43840 42460 43900 42470
rect 42770 42430 42850 42440
rect 43190 42430 43270 42440
rect 43610 42430 43690 42440
rect 42770 42420 42780 42430
rect 42630 42390 42780 42420
rect 42570 42370 42630 42380
rect 42770 42370 42780 42390
rect 42840 42370 42850 42430
rect 42770 42360 42850 42370
rect 43610 42370 43620 42430
rect 43680 42420 43690 42430
rect 43990 42430 44050 42440
rect 43680 42390 43990 42420
rect 43680 42370 43690 42390
rect 43610 42360 43690 42370
rect 43990 42360 44050 42370
rect 43180 42340 43280 42350
rect 43180 42270 43200 42340
rect 43270 42270 43280 42340
rect 43180 42230 43280 42270
rect 43180 42160 43200 42230
rect 43270 42160 43280 42230
rect 43180 42140 43280 42160
rect 42550 42130 42630 42140
rect 42550 42070 42560 42130
rect 42620 42110 42630 42130
rect 42770 42120 42850 42130
rect 42770 42110 42780 42120
rect 42620 42080 42780 42110
rect 42620 42070 42630 42080
rect 42550 42060 42630 42070
rect 42770 42060 42780 42080
rect 42840 42060 42850 42120
rect 43610 42120 43690 42130
rect 43610 42060 43620 42120
rect 43680 42110 43690 42120
rect 43990 42120 44070 42130
rect 43990 42110 44000 42120
rect 43680 42080 44000 42110
rect 43680 42060 43690 42080
rect 42770 42050 42850 42060
rect 43190 42050 43270 42060
rect 43610 42050 43690 42060
rect 43990 42060 44000 42080
rect 44060 42060 44070 42120
rect 43990 42050 44070 42060
rect 43190 41990 43200 42050
rect 43260 42010 43270 42050
rect 43260 42000 43960 42010
rect 43260 41990 43900 42000
rect 43190 41980 43900 41990
rect 43900 41930 43960 41940
rect 43840 40820 43900 40830
rect 43190 40790 43840 40800
rect 42570 40730 42630 40740
rect 43190 40730 43200 40790
rect 43260 40770 43840 40790
rect 43260 40730 43270 40770
rect 43840 40750 43900 40760
rect 43990 40730 44050 40740
rect 42770 40720 42850 40730
rect 43190 40720 43270 40730
rect 43610 40720 43690 40730
rect 42770 40710 42780 40720
rect 42630 40680 42780 40710
rect 42570 40660 42630 40670
rect 42770 40660 42780 40680
rect 42840 40660 42850 40720
rect 42770 40650 42850 40660
rect 43610 40660 43620 40720
rect 43680 40710 43690 40720
rect 43680 40680 43990 40710
rect 43680 40660 43690 40680
rect 43990 40660 44050 40670
rect 43610 40650 43690 40660
rect 43180 40630 43280 40640
rect 43180 40560 43200 40630
rect 43270 40560 43280 40630
rect 43180 40520 43280 40560
rect 43180 40450 43200 40520
rect 43270 40450 43280 40520
rect 43180 40430 43280 40450
rect 42550 40420 42630 40430
rect 43990 40420 44070 40430
rect 42550 40360 42560 40420
rect 42620 40400 42630 40420
rect 42770 40410 42850 40420
rect 42770 40400 42780 40410
rect 42620 40370 42780 40400
rect 42620 40360 42630 40370
rect 42550 40350 42630 40360
rect 42190 39290 42250 39300
rect 42190 39220 42250 39230
rect 42280 39270 42510 39300
rect 42070 36870 42150 36880
rect 42070 36810 42080 36870
rect 42140 36810 42150 36870
rect 42070 36800 42150 36810
rect 42010 36730 42090 36740
rect 42010 36670 42020 36730
rect 42080 36670 42090 36730
rect 42010 36660 42090 36670
rect 39360 36400 39370 36460
rect 39430 36400 39440 36460
rect 42190 36460 42220 39220
rect 42280 36600 42310 39270
rect 42600 39240 42630 40350
rect 42770 40350 42780 40370
rect 42840 40350 42850 40410
rect 43610 40410 43690 40420
rect 43610 40350 43620 40410
rect 43680 40400 43690 40410
rect 43990 40400 44000 40420
rect 43680 40370 44000 40400
rect 43680 40350 43690 40370
rect 43990 40360 44000 40370
rect 44060 40360 44070 40420
rect 43990 40350 44070 40360
rect 42770 40340 42850 40350
rect 43190 40340 43270 40350
rect 43610 40340 43690 40350
rect 43190 40280 43200 40340
rect 43260 40300 43270 40340
rect 43260 40290 43960 40300
rect 43260 40280 43900 40290
rect 43190 40270 43900 40280
rect 43900 40220 43960 40230
rect 43990 40210 44070 40220
rect 43990 40150 44000 40210
rect 44060 40150 44070 40210
rect 43990 40140 44070 40150
rect 42370 39230 42430 39240
rect 42370 39160 42430 39170
rect 42460 39210 42630 39240
rect 42660 39680 42740 39690
rect 42660 39620 42670 39680
rect 42730 39620 42740 39680
rect 43730 39680 43810 39690
rect 43730 39620 43740 39680
rect 43800 39620 43810 39680
rect 42250 36590 42330 36600
rect 42250 36530 42260 36590
rect 42320 36530 42330 36590
rect 42250 36520 42330 36530
rect 42190 36450 42270 36460
rect 42190 36390 42200 36450
rect 42260 36390 42270 36450
rect 42190 36380 42270 36390
rect 37380 36170 37460 36180
rect 32390 36100 32470 36110
rect 37380 36110 37390 36170
rect 37450 36110 37460 36170
rect 39180 36120 39190 36180
rect 39250 36120 39260 36180
rect 42370 36180 42400 39160
rect 42460 36320 42490 39210
rect 42660 38840 42730 39620
rect 43730 39610 43810 39620
rect 43900 39680 43960 39690
rect 43900 39610 43960 39620
rect 42660 38830 42740 38840
rect 42660 38770 42670 38830
rect 42730 38770 42740 38830
rect 42660 38760 42740 38770
rect 43740 38700 43810 39610
rect 43930 38700 43960 39610
rect 43990 39240 44020 40140
rect 44110 39300 44140 43760
rect 44230 39360 44260 47190
rect 44350 39420 44380 48900
rect 44470 39480 44500 50610
rect 44590 39540 44620 52320
rect 44710 39600 44740 54050
rect 46940 54090 47020 54100
rect 46940 54030 46950 54090
rect 47010 54080 47020 54090
rect 47760 54090 47840 54100
rect 47760 54080 47770 54090
rect 47010 54050 47770 54080
rect 47010 54030 47020 54050
rect 46940 54020 47020 54030
rect 47760 54030 47770 54050
rect 47830 54030 47840 54090
rect 48600 54090 48680 54100
rect 48600 54030 48610 54090
rect 48670 54080 48680 54090
rect 49580 54090 49660 54100
rect 49580 54080 49590 54090
rect 48670 54050 49590 54080
rect 48670 54030 48680 54050
rect 47760 54020 47840 54030
rect 48180 54020 48260 54030
rect 48600 54020 48680 54030
rect 49580 54030 49590 54050
rect 49650 54030 49660 54090
rect 49580 54020 49660 54030
rect 52170 54090 52250 54100
rect 52170 54030 52180 54090
rect 52240 54080 52250 54090
rect 52750 54090 52830 54100
rect 52750 54080 52760 54090
rect 52240 54050 52760 54080
rect 52240 54030 52250 54050
rect 52170 54020 52250 54030
rect 52750 54030 52760 54050
rect 52820 54030 52830 54090
rect 53590 54090 53670 54100
rect 53590 54030 53600 54090
rect 53660 54080 53670 54090
rect 54330 54090 54410 54100
rect 54330 54080 54340 54090
rect 53660 54050 54340 54080
rect 53660 54030 53670 54050
rect 52750 54020 52830 54030
rect 53170 54020 53250 54030
rect 53590 54020 53670 54030
rect 54330 54030 54340 54050
rect 54400 54030 54410 54090
rect 54330 54020 54410 54030
rect 57160 54090 57240 54100
rect 57160 54030 57170 54090
rect 57230 54080 57240 54090
rect 57740 54090 57820 54100
rect 57740 54080 57750 54090
rect 57230 54050 57750 54080
rect 57230 54030 57240 54050
rect 57160 54020 57240 54030
rect 57740 54030 57750 54050
rect 57810 54030 57820 54090
rect 58580 54090 58660 54100
rect 58580 54030 58590 54090
rect 58650 54080 58660 54090
rect 59320 54090 59400 54100
rect 59320 54080 59330 54090
rect 58650 54050 59330 54080
rect 58650 54030 58660 54050
rect 57740 54020 57820 54030
rect 58160 54020 58240 54030
rect 58580 54020 58660 54030
rect 59320 54030 59330 54050
rect 59390 54030 59400 54090
rect 59320 54020 59400 54030
rect 62390 54090 62470 54100
rect 62390 54030 62400 54090
rect 62460 54080 62470 54090
rect 62730 54090 62810 54100
rect 62730 54080 62740 54090
rect 62460 54050 62740 54080
rect 62460 54030 62470 54050
rect 62390 54020 62470 54030
rect 62730 54030 62740 54050
rect 62800 54030 62810 54090
rect 63570 54090 63650 54100
rect 63570 54030 63580 54090
rect 63640 54080 63650 54090
rect 64070 54090 64150 54100
rect 64070 54080 64080 54090
rect 63640 54050 64080 54080
rect 63640 54030 63650 54050
rect 62730 54020 62810 54030
rect 63150 54020 63230 54030
rect 63570 54020 63650 54030
rect 64070 54030 64080 54050
rect 64140 54030 64150 54090
rect 64070 54020 64150 54030
rect 67380 54090 67460 54100
rect 67380 54030 67390 54090
rect 67450 54080 67460 54090
rect 67720 54090 67800 54100
rect 67720 54080 67730 54090
rect 67450 54050 67730 54080
rect 67450 54030 67460 54050
rect 67380 54020 67460 54030
rect 67720 54030 67730 54050
rect 67790 54030 67800 54090
rect 68560 54090 68640 54100
rect 68560 54030 68570 54090
rect 68630 54080 68640 54090
rect 69060 54090 69140 54100
rect 69060 54080 69070 54090
rect 68630 54050 69070 54080
rect 68630 54030 68640 54050
rect 67720 54020 67800 54030
rect 68140 54020 68220 54030
rect 68560 54020 68640 54030
rect 69060 54030 69070 54050
rect 69130 54030 69140 54090
rect 69060 54020 69140 54030
rect 72490 54090 72570 54100
rect 72490 54030 72500 54090
rect 72560 54080 72570 54090
rect 72710 54090 72790 54100
rect 72710 54080 72720 54090
rect 72560 54050 72720 54080
rect 72560 54030 72570 54050
rect 72490 54020 72570 54030
rect 72710 54030 72720 54050
rect 72780 54030 72790 54090
rect 73550 54090 73630 54100
rect 73550 54030 73560 54090
rect 73620 54080 73630 54090
rect 73930 54090 74010 54100
rect 73930 54080 73940 54090
rect 73620 54050 73940 54080
rect 73620 54030 73630 54050
rect 72710 54020 72790 54030
rect 73130 54020 73210 54030
rect 73550 54020 73630 54030
rect 73930 54030 73940 54050
rect 74000 54030 74010 54090
rect 73930 54020 74010 54030
rect 77480 54090 77560 54100
rect 77480 54030 77490 54090
rect 77550 54080 77560 54090
rect 77700 54090 77780 54100
rect 77700 54080 77710 54090
rect 77550 54050 77710 54080
rect 77550 54030 77560 54050
rect 77480 54020 77560 54030
rect 77700 54030 77710 54050
rect 77770 54030 77780 54090
rect 78540 54090 78620 54100
rect 78540 54030 78550 54090
rect 78610 54080 78620 54090
rect 78920 54090 79000 54100
rect 78920 54080 78930 54090
rect 78610 54050 78930 54080
rect 78610 54030 78620 54050
rect 77700 54020 77780 54030
rect 78120 54020 78200 54030
rect 78540 54020 78620 54030
rect 78920 54030 78930 54050
rect 78990 54030 79000 54090
rect 78920 54020 79000 54030
rect 48180 53960 48190 54020
rect 48250 53980 48260 54020
rect 48250 53970 48950 53980
rect 48250 53960 48890 53970
rect 48180 53950 48890 53960
rect 53170 53960 53180 54020
rect 53240 53980 53250 54020
rect 53240 53970 53940 53980
rect 53240 53960 53880 53970
rect 53170 53950 53880 53960
rect 48890 53900 48950 53910
rect 58160 53960 58170 54020
rect 58230 53980 58240 54020
rect 58230 53970 58930 53980
rect 58230 53960 58870 53970
rect 58160 53950 58870 53960
rect 53880 53900 53940 53910
rect 63150 53960 63160 54020
rect 63220 53980 63230 54020
rect 63220 53970 63920 53980
rect 63220 53960 63860 53970
rect 63150 53950 63860 53960
rect 58870 53900 58930 53910
rect 68140 53960 68150 54020
rect 68210 53980 68220 54020
rect 68210 53970 68910 53980
rect 68210 53960 68850 53970
rect 68140 53950 68850 53960
rect 63860 53900 63920 53910
rect 73130 53960 73140 54020
rect 73200 53980 73210 54020
rect 73200 53970 73900 53980
rect 73200 53960 73840 53970
rect 73130 53950 73840 53960
rect 68850 53900 68910 53910
rect 78120 53960 78130 54020
rect 78190 53980 78200 54020
rect 78190 53970 78890 53980
rect 78190 53960 78830 53970
rect 78120 53950 78830 53960
rect 73840 53900 73900 53910
rect 78830 53900 78890 53910
rect 48830 52790 48890 52800
rect 48180 52760 48830 52770
rect 46960 52700 47020 52710
rect 48180 52700 48190 52760
rect 48250 52740 48830 52760
rect 48250 52700 48260 52740
rect 53820 52790 53880 52800
rect 48830 52720 48890 52730
rect 53170 52760 53820 52770
rect 49580 52700 49640 52710
rect 47760 52690 47840 52700
rect 48180 52690 48260 52700
rect 48600 52690 48680 52700
rect 47760 52680 47770 52690
rect 47020 52650 47770 52680
rect 46960 52630 47020 52640
rect 47760 52630 47770 52650
rect 47830 52630 47840 52690
rect 47760 52620 47840 52630
rect 48600 52630 48610 52690
rect 48670 52680 48680 52690
rect 48670 52650 49580 52680
rect 48670 52630 48680 52650
rect 49580 52630 49640 52640
rect 52190 52700 52250 52710
rect 53170 52700 53180 52760
rect 53240 52740 53820 52760
rect 53240 52700 53250 52740
rect 58810 52790 58870 52800
rect 53820 52720 53880 52730
rect 58160 52760 58810 52770
rect 54330 52700 54390 52710
rect 52750 52690 52830 52700
rect 53170 52690 53250 52700
rect 53590 52690 53670 52700
rect 52750 52680 52760 52690
rect 52250 52650 52760 52680
rect 52190 52630 52250 52640
rect 52750 52630 52760 52650
rect 52820 52630 52830 52690
rect 48600 52620 48680 52630
rect 52750 52620 52830 52630
rect 53590 52630 53600 52690
rect 53660 52680 53670 52690
rect 53660 52650 54330 52680
rect 53660 52630 53670 52650
rect 54330 52630 54390 52640
rect 57180 52700 57240 52710
rect 58160 52700 58170 52760
rect 58230 52740 58810 52760
rect 58230 52700 58240 52740
rect 63800 52790 63860 52800
rect 58810 52720 58870 52730
rect 63150 52760 63800 52770
rect 59320 52700 59380 52710
rect 57740 52690 57820 52700
rect 58160 52690 58240 52700
rect 58580 52690 58660 52700
rect 57740 52680 57750 52690
rect 57240 52650 57750 52680
rect 57180 52630 57240 52640
rect 57740 52630 57750 52650
rect 57810 52630 57820 52690
rect 53590 52620 53670 52630
rect 57740 52620 57820 52630
rect 58580 52630 58590 52690
rect 58650 52680 58660 52690
rect 58650 52650 59320 52680
rect 58650 52630 58660 52650
rect 59320 52630 59380 52640
rect 62410 52700 62470 52710
rect 63150 52700 63160 52760
rect 63220 52740 63800 52760
rect 63220 52700 63230 52740
rect 68790 52790 68850 52800
rect 63800 52720 63860 52730
rect 68140 52760 68790 52770
rect 64070 52700 64130 52710
rect 62730 52690 62810 52700
rect 63150 52690 63230 52700
rect 63570 52690 63650 52700
rect 62730 52680 62740 52690
rect 62470 52650 62740 52680
rect 62410 52630 62470 52640
rect 62730 52630 62740 52650
rect 62800 52630 62810 52690
rect 58580 52620 58660 52630
rect 62730 52620 62810 52630
rect 63570 52630 63580 52690
rect 63640 52680 63650 52690
rect 63640 52650 64070 52680
rect 63640 52630 63650 52650
rect 64070 52630 64130 52640
rect 67400 52700 67460 52710
rect 68140 52700 68150 52760
rect 68210 52740 68790 52760
rect 68210 52700 68220 52740
rect 73780 52790 73840 52800
rect 68790 52720 68850 52730
rect 73130 52760 73780 52770
rect 69060 52700 69120 52710
rect 67720 52690 67800 52700
rect 68140 52690 68220 52700
rect 68560 52690 68640 52700
rect 67720 52680 67730 52690
rect 67460 52650 67730 52680
rect 67400 52630 67460 52640
rect 67720 52630 67730 52650
rect 67790 52630 67800 52690
rect 63570 52620 63650 52630
rect 67720 52620 67800 52630
rect 68560 52630 68570 52690
rect 68630 52680 68640 52690
rect 68630 52650 69060 52680
rect 68630 52630 68640 52650
rect 69060 52630 69120 52640
rect 72510 52700 72570 52710
rect 73130 52700 73140 52760
rect 73200 52740 73780 52760
rect 73200 52700 73210 52740
rect 78770 52790 78830 52800
rect 73780 52720 73840 52730
rect 78120 52760 78770 52770
rect 73930 52700 73990 52710
rect 72710 52690 72790 52700
rect 73130 52690 73210 52700
rect 73550 52690 73630 52700
rect 72710 52680 72720 52690
rect 72570 52650 72720 52680
rect 72510 52630 72570 52640
rect 72710 52630 72720 52650
rect 72780 52630 72790 52690
rect 68560 52620 68640 52630
rect 72710 52620 72790 52630
rect 73550 52630 73560 52690
rect 73620 52680 73630 52690
rect 73620 52650 73930 52680
rect 73620 52630 73630 52650
rect 73930 52630 73990 52640
rect 77500 52700 77560 52710
rect 78120 52700 78130 52760
rect 78190 52740 78770 52760
rect 78190 52700 78200 52740
rect 78770 52720 78830 52730
rect 78920 52700 78980 52710
rect 77700 52690 77780 52700
rect 78120 52690 78200 52700
rect 78540 52690 78620 52700
rect 77700 52680 77710 52690
rect 77560 52650 77710 52680
rect 77500 52630 77560 52640
rect 77700 52630 77710 52650
rect 77770 52630 77780 52690
rect 73550 52620 73630 52630
rect 77700 52620 77780 52630
rect 78540 52630 78550 52690
rect 78610 52680 78620 52690
rect 78610 52650 78920 52680
rect 78610 52630 78620 52650
rect 78920 52630 78980 52640
rect 78540 52620 78620 52630
rect 48170 52600 48270 52610
rect 48170 52530 48190 52600
rect 48260 52530 48270 52600
rect 48170 52490 48270 52530
rect 48170 52420 48190 52490
rect 48260 52420 48270 52490
rect 48170 52400 48270 52420
rect 53160 52600 53260 52610
rect 53160 52530 53180 52600
rect 53250 52530 53260 52600
rect 53160 52490 53260 52530
rect 53160 52420 53180 52490
rect 53250 52420 53260 52490
rect 53160 52400 53260 52420
rect 58150 52600 58250 52610
rect 58150 52530 58170 52600
rect 58240 52530 58250 52600
rect 58150 52490 58250 52530
rect 58150 52420 58170 52490
rect 58240 52420 58250 52490
rect 58150 52400 58250 52420
rect 63140 52600 63240 52610
rect 63140 52530 63160 52600
rect 63230 52530 63240 52600
rect 63140 52490 63240 52530
rect 63140 52420 63160 52490
rect 63230 52420 63240 52490
rect 63140 52400 63240 52420
rect 68130 52600 68230 52610
rect 68130 52530 68150 52600
rect 68220 52530 68230 52600
rect 68130 52490 68230 52530
rect 68130 52420 68150 52490
rect 68220 52420 68230 52490
rect 68130 52400 68230 52420
rect 73120 52600 73220 52610
rect 73120 52530 73140 52600
rect 73210 52530 73220 52600
rect 73120 52490 73220 52530
rect 73120 52420 73140 52490
rect 73210 52420 73220 52490
rect 73120 52400 73220 52420
rect 78110 52600 78210 52610
rect 78110 52530 78130 52600
rect 78200 52530 78210 52600
rect 78110 52490 78210 52530
rect 78110 52420 78130 52490
rect 78200 52420 78210 52490
rect 78110 52400 78210 52420
rect 46940 52380 47020 52390
rect 46940 52320 46950 52380
rect 47010 52370 47020 52380
rect 47760 52380 47840 52390
rect 47760 52370 47770 52380
rect 47010 52340 47770 52370
rect 47010 52320 47020 52340
rect 46940 52310 47020 52320
rect 47760 52320 47770 52340
rect 47830 52320 47840 52380
rect 48600 52380 48680 52390
rect 48600 52320 48610 52380
rect 48670 52370 48680 52380
rect 49580 52380 49660 52390
rect 49580 52370 49590 52380
rect 48670 52340 49590 52370
rect 48670 52320 48680 52340
rect 47760 52310 47840 52320
rect 48180 52310 48260 52320
rect 48600 52310 48680 52320
rect 49580 52320 49590 52340
rect 49650 52320 49660 52380
rect 49580 52310 49660 52320
rect 52170 52380 52250 52390
rect 52170 52320 52180 52380
rect 52240 52370 52250 52380
rect 52750 52380 52830 52390
rect 52750 52370 52760 52380
rect 52240 52340 52760 52370
rect 52240 52320 52250 52340
rect 52170 52310 52250 52320
rect 52750 52320 52760 52340
rect 52820 52320 52830 52380
rect 53590 52380 53670 52390
rect 53590 52320 53600 52380
rect 53660 52370 53670 52380
rect 54330 52380 54410 52390
rect 54330 52370 54340 52380
rect 53660 52340 54340 52370
rect 53660 52320 53670 52340
rect 52750 52310 52830 52320
rect 53170 52310 53250 52320
rect 53590 52310 53670 52320
rect 54330 52320 54340 52340
rect 54400 52320 54410 52380
rect 54330 52310 54410 52320
rect 57160 52380 57240 52390
rect 57160 52320 57170 52380
rect 57230 52370 57240 52380
rect 57740 52380 57820 52390
rect 57740 52370 57750 52380
rect 57230 52340 57750 52370
rect 57230 52320 57240 52340
rect 57160 52310 57240 52320
rect 57740 52320 57750 52340
rect 57810 52320 57820 52380
rect 58580 52380 58660 52390
rect 58580 52320 58590 52380
rect 58650 52370 58660 52380
rect 59320 52380 59400 52390
rect 59320 52370 59330 52380
rect 58650 52340 59330 52370
rect 58650 52320 58660 52340
rect 57740 52310 57820 52320
rect 58160 52310 58240 52320
rect 58580 52310 58660 52320
rect 59320 52320 59330 52340
rect 59390 52320 59400 52380
rect 59320 52310 59400 52320
rect 62390 52380 62470 52390
rect 62390 52320 62400 52380
rect 62460 52370 62470 52380
rect 62730 52380 62810 52390
rect 62730 52370 62740 52380
rect 62460 52340 62740 52370
rect 62460 52320 62470 52340
rect 62390 52310 62470 52320
rect 62730 52320 62740 52340
rect 62800 52320 62810 52380
rect 63570 52380 63650 52390
rect 63570 52320 63580 52380
rect 63640 52370 63650 52380
rect 64070 52380 64150 52390
rect 64070 52370 64080 52380
rect 63640 52340 64080 52370
rect 63640 52320 63650 52340
rect 62730 52310 62810 52320
rect 63150 52310 63230 52320
rect 63570 52310 63650 52320
rect 64070 52320 64080 52340
rect 64140 52320 64150 52380
rect 64070 52310 64150 52320
rect 67380 52380 67460 52390
rect 67380 52320 67390 52380
rect 67450 52370 67460 52380
rect 67720 52380 67800 52390
rect 67720 52370 67730 52380
rect 67450 52340 67730 52370
rect 67450 52320 67460 52340
rect 67380 52310 67460 52320
rect 67720 52320 67730 52340
rect 67790 52320 67800 52380
rect 68560 52380 68640 52390
rect 68560 52320 68570 52380
rect 68630 52370 68640 52380
rect 69060 52380 69140 52390
rect 69060 52370 69070 52380
rect 68630 52340 69070 52370
rect 68630 52320 68640 52340
rect 67720 52310 67800 52320
rect 68140 52310 68220 52320
rect 68560 52310 68640 52320
rect 69060 52320 69070 52340
rect 69130 52320 69140 52380
rect 69060 52310 69140 52320
rect 72490 52380 72570 52390
rect 72490 52320 72500 52380
rect 72560 52370 72570 52380
rect 72710 52380 72790 52390
rect 72710 52370 72720 52380
rect 72560 52340 72720 52370
rect 72560 52320 72570 52340
rect 72490 52310 72570 52320
rect 72710 52320 72720 52340
rect 72780 52320 72790 52380
rect 73550 52380 73630 52390
rect 73550 52320 73560 52380
rect 73620 52370 73630 52380
rect 73930 52380 74010 52390
rect 73930 52370 73940 52380
rect 73620 52340 73940 52370
rect 73620 52320 73630 52340
rect 72710 52310 72790 52320
rect 73130 52310 73210 52320
rect 73550 52310 73630 52320
rect 73930 52320 73940 52340
rect 74000 52320 74010 52380
rect 73930 52310 74010 52320
rect 77480 52380 77560 52390
rect 77480 52320 77490 52380
rect 77550 52370 77560 52380
rect 77700 52380 77780 52390
rect 77700 52370 77710 52380
rect 77550 52340 77710 52370
rect 77550 52320 77560 52340
rect 77480 52310 77560 52320
rect 77700 52320 77710 52340
rect 77770 52320 77780 52380
rect 78540 52380 78620 52390
rect 78540 52320 78550 52380
rect 78610 52370 78620 52380
rect 78920 52380 79000 52390
rect 78920 52370 78930 52380
rect 78610 52340 78930 52370
rect 78610 52320 78620 52340
rect 77700 52310 77780 52320
rect 78120 52310 78200 52320
rect 78540 52310 78620 52320
rect 78920 52320 78930 52340
rect 78990 52320 79000 52380
rect 78920 52310 79000 52320
rect 44710 39570 45240 39600
rect 44590 39510 45060 39540
rect 44470 39450 44880 39480
rect 44350 39390 44700 39420
rect 44230 39330 44520 39360
rect 44110 39270 44340 39300
rect 43990 39210 44160 39240
rect 43730 38690 43810 38700
rect 43730 38630 43740 38690
rect 43800 38630 43810 38690
rect 43880 38640 43890 38700
rect 43950 38640 43960 38700
rect 43730 38620 43810 38630
rect 44130 36320 44160 39210
rect 44190 39230 44250 39240
rect 44190 39160 44250 39170
rect 42430 36310 42510 36320
rect 42430 36250 42440 36310
rect 42500 36250 42510 36310
rect 44110 36260 44120 36320
rect 44180 36260 44190 36320
rect 42430 36240 42510 36250
rect 44220 36180 44250 39160
rect 44310 36600 44340 39270
rect 44370 39290 44430 39300
rect 44370 39220 44430 39230
rect 44290 36540 44300 36600
rect 44360 36540 44370 36600
rect 44400 36460 44430 39220
rect 44490 36880 44520 39330
rect 44550 39350 44610 39360
rect 44550 39280 44610 39290
rect 44470 36820 44480 36880
rect 44540 36820 44550 36880
rect 44580 36740 44610 39280
rect 44670 37160 44700 39390
rect 44730 39410 44790 39420
rect 44730 39340 44790 39350
rect 44650 37100 44660 37160
rect 44720 37100 44730 37160
rect 44760 37020 44790 39340
rect 44850 37440 44880 39450
rect 44910 39470 44970 39480
rect 44910 39400 44970 39410
rect 44830 37380 44840 37440
rect 44900 37380 44910 37440
rect 44940 37300 44970 39400
rect 45030 38280 45060 39510
rect 45090 39530 45150 39540
rect 45090 39460 45150 39470
rect 45010 38220 45020 38280
rect 45080 38220 45090 38280
rect 45120 38140 45150 39460
rect 45100 38080 45110 38140
rect 45170 38080 45180 38140
rect 45210 38000 45240 39570
rect 45270 39590 45330 39600
rect 46990 39540 47020 52310
rect 48180 52250 48190 52310
rect 48250 52270 48260 52310
rect 48250 52260 48950 52270
rect 48250 52250 48890 52260
rect 48180 52240 48890 52250
rect 48890 52190 48950 52200
rect 48830 51080 48890 51090
rect 48180 51050 48830 51060
rect 47080 50990 47140 51000
rect 48180 50990 48190 51050
rect 48250 51030 48830 51050
rect 48250 50990 48260 51030
rect 48830 51010 48890 51020
rect 49460 50990 49520 51000
rect 47760 50980 47840 50990
rect 48180 50980 48260 50990
rect 48600 50980 48680 50990
rect 47760 50970 47770 50980
rect 47140 50940 47770 50970
rect 47080 50920 47140 50930
rect 47760 50920 47770 50940
rect 47830 50920 47840 50980
rect 47760 50910 47840 50920
rect 48600 50920 48610 50980
rect 48670 50970 48680 50980
rect 48670 50940 49460 50970
rect 48670 50920 48680 50940
rect 49460 50920 49520 50930
rect 48600 50910 48680 50920
rect 48170 50890 48270 50900
rect 48170 50820 48190 50890
rect 48260 50820 48270 50890
rect 48170 50780 48270 50820
rect 48170 50710 48190 50780
rect 48260 50710 48270 50780
rect 48170 50690 48270 50710
rect 47060 50670 47140 50680
rect 47060 50610 47070 50670
rect 47130 50660 47140 50670
rect 47760 50670 47840 50680
rect 47760 50660 47770 50670
rect 47130 50630 47770 50660
rect 47130 50610 47140 50630
rect 47060 50600 47140 50610
rect 47760 50610 47770 50630
rect 47830 50610 47840 50670
rect 48600 50670 48680 50680
rect 48600 50610 48610 50670
rect 48670 50660 48680 50670
rect 49460 50670 49540 50680
rect 49460 50660 49470 50670
rect 48670 50630 49470 50660
rect 48670 50610 48680 50630
rect 47760 50600 47840 50610
rect 48180 50600 48260 50610
rect 48600 50600 48680 50610
rect 49460 50610 49470 50630
rect 49530 50610 49540 50670
rect 49460 50600 49540 50610
rect 45270 39520 45330 39530
rect 45190 37940 45200 38000
rect 45260 37940 45270 38000
rect 45300 37860 45330 39520
rect 45250 37800 45260 37860
rect 45320 37800 45330 37860
rect 46460 39530 46520 39540
rect 46460 39460 46520 39470
rect 46550 39510 47020 39540
rect 44890 37240 44900 37300
rect 44960 37240 44970 37300
rect 46460 37300 46490 39460
rect 46550 37440 46580 39510
rect 47110 39480 47140 50600
rect 48180 50540 48190 50600
rect 48250 50560 48260 50600
rect 48250 50550 48950 50560
rect 48250 50540 48890 50550
rect 48180 50530 48890 50540
rect 48890 50480 48950 50490
rect 48830 49370 48890 49380
rect 48180 49340 48830 49350
rect 47200 49280 47260 49290
rect 48180 49280 48190 49340
rect 48250 49320 48830 49340
rect 48250 49280 48260 49320
rect 48830 49300 48890 49310
rect 49340 49280 49400 49290
rect 47760 49270 47840 49280
rect 48180 49270 48260 49280
rect 48600 49270 48680 49280
rect 47760 49260 47770 49270
rect 47260 49230 47770 49260
rect 47200 49210 47260 49220
rect 47760 49210 47770 49230
rect 47830 49210 47840 49270
rect 47760 49200 47840 49210
rect 48600 49210 48610 49270
rect 48670 49260 48680 49270
rect 48670 49230 49340 49260
rect 48670 49210 48680 49230
rect 49340 49210 49400 49220
rect 48600 49200 48680 49210
rect 48170 49180 48270 49190
rect 48170 49110 48190 49180
rect 48260 49110 48270 49180
rect 48170 49070 48270 49110
rect 48170 49000 48190 49070
rect 48260 49000 48270 49070
rect 48170 48980 48270 49000
rect 47180 48960 47260 48970
rect 47180 48900 47190 48960
rect 47250 48950 47260 48960
rect 47760 48960 47840 48970
rect 47760 48950 47770 48960
rect 47250 48920 47770 48950
rect 47250 48900 47260 48920
rect 47180 48890 47260 48900
rect 47760 48900 47770 48920
rect 47830 48900 47840 48960
rect 48600 48960 48680 48970
rect 48600 48900 48610 48960
rect 48670 48950 48680 48960
rect 49340 48960 49420 48970
rect 49340 48950 49350 48960
rect 48670 48920 49350 48950
rect 48670 48900 48680 48920
rect 47760 48890 47840 48900
rect 48180 48890 48260 48900
rect 48600 48890 48680 48900
rect 49340 48900 49350 48920
rect 49410 48900 49420 48960
rect 49340 48890 49420 48900
rect 46640 39470 46700 39480
rect 46640 39400 46700 39410
rect 46730 39450 47140 39480
rect 46640 37580 46670 39400
rect 46730 37720 46760 39450
rect 47230 39420 47260 48890
rect 48180 48830 48190 48890
rect 48250 48850 48260 48890
rect 48250 48840 48950 48850
rect 48250 48830 48890 48840
rect 48180 48820 48890 48830
rect 48890 48770 48950 48780
rect 48830 47660 48890 47670
rect 48180 47630 48830 47640
rect 47320 47570 47380 47580
rect 48180 47570 48190 47630
rect 48250 47610 48830 47630
rect 48250 47570 48260 47610
rect 48830 47590 48890 47600
rect 49220 47570 49280 47580
rect 47760 47560 47840 47570
rect 48180 47560 48260 47570
rect 48600 47560 48680 47570
rect 47760 47550 47770 47560
rect 47380 47520 47770 47550
rect 47320 47500 47380 47510
rect 47760 47500 47770 47520
rect 47830 47500 47840 47560
rect 47760 47490 47840 47500
rect 48600 47500 48610 47560
rect 48670 47550 48680 47560
rect 48670 47520 49220 47550
rect 48670 47500 48680 47520
rect 49220 47500 49280 47510
rect 48600 47490 48680 47500
rect 48170 47470 48270 47480
rect 48170 47400 48190 47470
rect 48260 47400 48270 47470
rect 48170 47360 48270 47400
rect 48170 47290 48190 47360
rect 48260 47290 48270 47360
rect 48170 47270 48270 47290
rect 47300 47250 47380 47260
rect 47300 47190 47310 47250
rect 47370 47240 47380 47250
rect 47760 47250 47840 47260
rect 47760 47240 47770 47250
rect 47370 47210 47770 47240
rect 47370 47190 47380 47210
rect 47300 47180 47380 47190
rect 47760 47190 47770 47210
rect 47830 47190 47840 47250
rect 48600 47250 48680 47260
rect 48600 47190 48610 47250
rect 48670 47240 48680 47250
rect 49220 47250 49300 47260
rect 49220 47240 49230 47250
rect 48670 47210 49230 47240
rect 48670 47190 48680 47210
rect 47760 47180 47840 47190
rect 48180 47180 48260 47190
rect 48600 47180 48680 47190
rect 49220 47190 49230 47210
rect 49290 47190 49300 47250
rect 49220 47180 49300 47190
rect 46820 39410 46880 39420
rect 46820 39340 46880 39350
rect 46910 39390 47260 39420
rect 46700 37710 46780 37720
rect 46700 37650 46710 37710
rect 46770 37650 46780 37710
rect 46700 37640 46780 37650
rect 46640 37570 46720 37580
rect 46640 37510 46650 37570
rect 46710 37510 46720 37570
rect 46640 37500 46720 37510
rect 46520 37430 46600 37440
rect 46520 37370 46530 37430
rect 46590 37370 46600 37430
rect 46520 37360 46600 37370
rect 46460 37290 46540 37300
rect 46460 37230 46470 37290
rect 46530 37230 46540 37290
rect 46460 37220 46540 37230
rect 44710 36960 44720 37020
rect 44780 36960 44790 37020
rect 46820 37020 46850 39340
rect 46910 37160 46940 39390
rect 47350 39360 47380 47180
rect 48180 47120 48190 47180
rect 48250 47140 48260 47180
rect 48250 47130 48950 47140
rect 48250 47120 48890 47130
rect 48180 47110 48890 47120
rect 48890 47060 48950 47070
rect 48830 45950 48890 45960
rect 48180 45920 48830 45930
rect 47440 45860 47500 45870
rect 48180 45860 48190 45920
rect 48250 45900 48830 45920
rect 48250 45860 48260 45900
rect 48830 45880 48890 45890
rect 49100 45860 49160 45870
rect 47760 45850 47840 45860
rect 48180 45850 48260 45860
rect 48600 45850 48680 45860
rect 47760 45840 47770 45850
rect 47500 45810 47770 45840
rect 47440 45790 47500 45800
rect 47760 45790 47770 45810
rect 47830 45790 47840 45850
rect 47760 45780 47840 45790
rect 48600 45790 48610 45850
rect 48670 45840 48680 45850
rect 48670 45810 49100 45840
rect 48670 45790 48680 45810
rect 49100 45790 49160 45800
rect 48600 45780 48680 45790
rect 48170 45760 48270 45770
rect 48170 45690 48190 45760
rect 48260 45690 48270 45760
rect 48170 45650 48270 45690
rect 48170 45580 48190 45650
rect 48260 45580 48270 45650
rect 48170 45560 48270 45580
rect 47420 45540 47500 45550
rect 47420 45480 47430 45540
rect 47490 45530 47500 45540
rect 47760 45540 47840 45550
rect 47760 45530 47770 45540
rect 47490 45500 47770 45530
rect 47490 45480 47500 45500
rect 47420 45470 47500 45480
rect 47760 45480 47770 45500
rect 47830 45480 47840 45540
rect 48600 45540 48680 45550
rect 48600 45480 48610 45540
rect 48670 45530 48680 45540
rect 49100 45540 49180 45550
rect 49100 45530 49110 45540
rect 48670 45500 49110 45530
rect 48670 45480 48680 45500
rect 47760 45470 47840 45480
rect 48180 45470 48260 45480
rect 48600 45470 48680 45480
rect 49100 45480 49110 45500
rect 49170 45480 49180 45540
rect 49100 45470 49180 45480
rect 48180 45410 48190 45470
rect 48250 45430 48260 45470
rect 48250 45420 48950 45430
rect 48250 45410 48890 45420
rect 48180 45400 48890 45410
rect 48890 45350 48950 45360
rect 48830 44240 48890 44250
rect 48180 44210 48830 44220
rect 47440 44150 47500 44160
rect 48180 44150 48190 44210
rect 48250 44190 48830 44210
rect 48250 44150 48260 44190
rect 48830 44170 48890 44180
rect 49100 44150 49160 44160
rect 47760 44140 47840 44150
rect 48180 44140 48260 44150
rect 48600 44140 48680 44150
rect 47760 44130 47770 44140
rect 47500 44100 47770 44130
rect 47440 44080 47500 44090
rect 47760 44080 47770 44100
rect 47830 44080 47840 44140
rect 47760 44070 47840 44080
rect 48600 44080 48610 44140
rect 48670 44130 48680 44140
rect 48670 44100 49100 44130
rect 48670 44080 48680 44100
rect 49100 44080 49160 44090
rect 48600 44070 48680 44080
rect 48170 44050 48270 44060
rect 48170 43980 48190 44050
rect 48260 43980 48270 44050
rect 48170 43940 48270 43980
rect 48170 43870 48190 43940
rect 48260 43870 48270 43940
rect 48170 43850 48270 43870
rect 47420 43830 47500 43840
rect 47420 43770 47430 43830
rect 47490 43820 47500 43830
rect 47760 43830 47840 43840
rect 47760 43820 47770 43830
rect 47490 43790 47770 43820
rect 47490 43770 47500 43790
rect 47420 43760 47500 43770
rect 47760 43770 47770 43790
rect 47830 43770 47840 43830
rect 48600 43830 48680 43840
rect 48600 43770 48610 43830
rect 48670 43820 48680 43830
rect 49100 43830 49180 43840
rect 49100 43820 49110 43830
rect 48670 43790 49110 43820
rect 48670 43770 48680 43790
rect 47760 43760 47840 43770
rect 48180 43760 48260 43770
rect 48600 43760 48680 43770
rect 49100 43770 49110 43790
rect 49170 43770 49180 43830
rect 49100 43760 49180 43770
rect 47000 39350 47060 39360
rect 47000 39280 47060 39290
rect 47090 39330 47380 39360
rect 46880 37150 46960 37160
rect 46880 37090 46890 37150
rect 46950 37090 46960 37150
rect 46880 37080 46960 37090
rect 46820 37010 46900 37020
rect 46820 36950 46830 37010
rect 46890 36950 46900 37010
rect 46820 36940 46900 36950
rect 44530 36680 44540 36740
rect 44600 36680 44610 36740
rect 47000 36740 47030 39280
rect 47090 36880 47120 39330
rect 47470 39300 47500 43760
rect 48180 43700 48190 43760
rect 48250 43720 48260 43760
rect 48250 43710 48950 43720
rect 48250 43700 48890 43710
rect 48180 43690 48890 43700
rect 48890 43640 48950 43650
rect 48830 42530 48890 42540
rect 48180 42500 48830 42510
rect 47560 42440 47620 42450
rect 48180 42440 48190 42500
rect 48250 42480 48830 42500
rect 48250 42440 48260 42480
rect 48830 42460 48890 42470
rect 48980 42440 49040 42450
rect 47760 42430 47840 42440
rect 48180 42430 48260 42440
rect 48600 42430 48680 42440
rect 47760 42420 47770 42430
rect 47620 42390 47770 42420
rect 47560 42370 47620 42380
rect 47760 42370 47770 42390
rect 47830 42370 47840 42430
rect 47760 42360 47840 42370
rect 48600 42370 48610 42430
rect 48670 42420 48680 42430
rect 48670 42390 48980 42420
rect 48670 42370 48680 42390
rect 48980 42370 49040 42380
rect 48600 42360 48680 42370
rect 48170 42340 48270 42350
rect 48170 42270 48190 42340
rect 48260 42270 48270 42340
rect 48170 42230 48270 42270
rect 48170 42160 48190 42230
rect 48260 42160 48270 42230
rect 48170 42140 48270 42160
rect 47540 42120 47620 42130
rect 47540 42060 47550 42120
rect 47610 42110 47620 42120
rect 47760 42120 47840 42130
rect 47760 42110 47770 42120
rect 47610 42080 47770 42110
rect 47610 42060 47620 42080
rect 47540 42050 47620 42060
rect 47760 42060 47770 42080
rect 47830 42060 47840 42120
rect 48600 42120 48680 42130
rect 48600 42060 48610 42120
rect 48670 42110 48680 42120
rect 48980 42120 49060 42130
rect 48980 42110 48990 42120
rect 48670 42080 48990 42110
rect 48670 42060 48680 42080
rect 47760 42050 47840 42060
rect 48180 42050 48260 42060
rect 48600 42050 48680 42060
rect 48980 42060 48990 42080
rect 49050 42060 49060 42120
rect 48980 42050 49060 42060
rect 48180 41990 48190 42050
rect 48250 42010 48260 42050
rect 48250 42000 48950 42010
rect 48250 41990 48890 42000
rect 48180 41980 48890 41990
rect 48890 41930 48950 41940
rect 48830 40820 48890 40830
rect 48180 40790 48830 40800
rect 47560 40730 47620 40740
rect 48180 40730 48190 40790
rect 48250 40770 48830 40790
rect 48250 40730 48260 40770
rect 48830 40750 48890 40760
rect 48980 40730 49040 40740
rect 47760 40720 47840 40730
rect 48180 40720 48260 40730
rect 48600 40720 48680 40730
rect 47760 40710 47770 40720
rect 47620 40680 47770 40710
rect 47560 40660 47620 40670
rect 47760 40660 47770 40680
rect 47830 40660 47840 40720
rect 47760 40650 47840 40660
rect 48600 40660 48610 40720
rect 48670 40710 48680 40720
rect 48670 40680 48980 40710
rect 48670 40660 48680 40680
rect 48980 40660 49040 40670
rect 48600 40650 48680 40660
rect 48170 40630 48270 40640
rect 48170 40560 48190 40630
rect 48260 40560 48270 40630
rect 48170 40520 48270 40560
rect 48170 40450 48190 40520
rect 48260 40450 48270 40520
rect 48170 40430 48270 40450
rect 47540 40410 47620 40420
rect 47540 40350 47550 40410
rect 47610 40400 47620 40410
rect 47760 40410 47840 40420
rect 47760 40400 47770 40410
rect 47610 40370 47770 40400
rect 47610 40350 47620 40370
rect 47540 40340 47620 40350
rect 47760 40350 47770 40370
rect 47830 40350 47840 40410
rect 48600 40410 48680 40420
rect 48600 40350 48610 40410
rect 48670 40400 48680 40410
rect 48980 40410 49060 40420
rect 48980 40400 48990 40410
rect 48670 40370 48990 40400
rect 48670 40350 48680 40370
rect 47760 40340 47840 40350
rect 48180 40340 48260 40350
rect 48600 40340 48680 40350
rect 48980 40350 48990 40370
rect 49050 40350 49060 40410
rect 48980 40340 49060 40350
rect 47180 39290 47240 39300
rect 47180 39220 47240 39230
rect 47270 39270 47500 39300
rect 47060 36870 47140 36880
rect 47060 36810 47070 36870
rect 47130 36810 47140 36870
rect 47060 36800 47140 36810
rect 47000 36730 47080 36740
rect 47000 36670 47010 36730
rect 47070 36670 47080 36730
rect 47000 36660 47080 36670
rect 44350 36400 44360 36460
rect 44420 36400 44430 36460
rect 47180 36460 47210 39220
rect 47270 36600 47300 39270
rect 47590 39240 47620 40340
rect 48180 40280 48190 40340
rect 48250 40300 48260 40340
rect 48250 40290 48950 40300
rect 48250 40280 48890 40290
rect 48180 40270 48890 40280
rect 48890 40220 48950 40230
rect 47360 39230 47420 39240
rect 47360 39160 47420 39170
rect 47450 39210 47620 39240
rect 47650 39680 47730 39690
rect 47650 39620 47660 39680
rect 47720 39620 47730 39680
rect 48720 39680 48800 39690
rect 48720 39620 48730 39680
rect 48790 39620 48800 39680
rect 47240 36590 47320 36600
rect 47240 36530 47250 36590
rect 47310 36530 47320 36590
rect 47240 36520 47320 36530
rect 47180 36450 47260 36460
rect 47180 36390 47190 36450
rect 47250 36390 47260 36450
rect 47180 36380 47260 36390
rect 42370 36170 42450 36180
rect 37380 36100 37460 36110
rect 42370 36110 42380 36170
rect 42440 36110 42450 36170
rect 44170 36120 44180 36180
rect 44240 36120 44250 36180
rect 47360 36180 47390 39160
rect 47450 36320 47480 39210
rect 47650 38840 47720 39620
rect 48720 39610 48800 39620
rect 48890 39680 48950 39690
rect 48890 39610 48950 39620
rect 47650 38830 47730 38840
rect 47650 38770 47660 38830
rect 47720 38770 47730 38830
rect 47650 38760 47730 38770
rect 48730 38700 48800 39610
rect 48920 38700 48950 39610
rect 48980 39240 49010 40340
rect 49100 39300 49130 43760
rect 49220 39360 49250 47180
rect 49340 39420 49370 48890
rect 49460 39480 49490 50600
rect 49580 39540 49610 52310
rect 53170 52250 53180 52310
rect 53240 52270 53250 52310
rect 53240 52260 53940 52270
rect 53240 52250 53880 52260
rect 53170 52240 53880 52250
rect 58160 52250 58170 52310
rect 58230 52270 58240 52310
rect 58230 52260 58930 52270
rect 58230 52250 58870 52260
rect 58160 52240 58870 52250
rect 53880 52190 53940 52200
rect 63150 52250 63160 52310
rect 63220 52270 63230 52310
rect 63220 52260 63920 52270
rect 63220 52250 63860 52260
rect 63150 52240 63860 52250
rect 58870 52190 58930 52200
rect 68140 52250 68150 52310
rect 68210 52270 68220 52310
rect 68210 52260 68910 52270
rect 68210 52250 68850 52260
rect 68140 52240 68850 52250
rect 63860 52190 63920 52200
rect 73130 52250 73140 52310
rect 73200 52270 73210 52310
rect 73200 52260 73900 52270
rect 73200 52250 73840 52260
rect 73130 52240 73840 52250
rect 68850 52190 68910 52200
rect 78120 52250 78130 52310
rect 78190 52270 78200 52310
rect 78190 52260 78890 52270
rect 78190 52250 78830 52260
rect 78120 52240 78830 52250
rect 73840 52190 73900 52200
rect 78830 52190 78890 52200
rect 53820 51080 53880 51090
rect 53170 51050 53820 51060
rect 52190 50990 52250 51000
rect 53170 50990 53180 51050
rect 53240 51030 53820 51050
rect 53240 50990 53250 51030
rect 58810 51080 58870 51090
rect 53820 51010 53880 51020
rect 58160 51050 58810 51060
rect 54330 50990 54390 51000
rect 52750 50980 52830 50990
rect 53170 50980 53250 50990
rect 53590 50980 53670 50990
rect 52750 50970 52760 50980
rect 52250 50940 52760 50970
rect 52190 50920 52250 50930
rect 52750 50920 52760 50940
rect 52820 50920 52830 50980
rect 52750 50910 52830 50920
rect 53590 50920 53600 50980
rect 53660 50970 53670 50980
rect 53660 50940 54330 50970
rect 53660 50920 53670 50940
rect 54330 50920 54390 50930
rect 57180 50990 57240 51000
rect 58160 50990 58170 51050
rect 58230 51030 58810 51050
rect 58230 50990 58240 51030
rect 63800 51080 63860 51090
rect 58810 51010 58870 51020
rect 63150 51050 63800 51060
rect 59320 50990 59380 51000
rect 57740 50980 57820 50990
rect 58160 50980 58240 50990
rect 58580 50980 58660 50990
rect 57740 50970 57750 50980
rect 57240 50940 57750 50970
rect 57180 50920 57240 50930
rect 57740 50920 57750 50940
rect 57810 50920 57820 50980
rect 53590 50910 53670 50920
rect 57740 50910 57820 50920
rect 58580 50920 58590 50980
rect 58650 50970 58660 50980
rect 58650 50940 59320 50970
rect 58650 50920 58660 50940
rect 59320 50920 59380 50930
rect 62410 50990 62470 51000
rect 63150 50990 63160 51050
rect 63220 51030 63800 51050
rect 63220 50990 63230 51030
rect 68790 51080 68850 51090
rect 63800 51010 63860 51020
rect 68140 51050 68790 51060
rect 64070 50990 64130 51000
rect 62730 50980 62810 50990
rect 63150 50980 63230 50990
rect 63570 50980 63650 50990
rect 62730 50970 62740 50980
rect 62470 50940 62740 50970
rect 62410 50920 62470 50930
rect 62730 50920 62740 50940
rect 62800 50920 62810 50980
rect 58580 50910 58660 50920
rect 62730 50910 62810 50920
rect 63570 50920 63580 50980
rect 63640 50970 63650 50980
rect 63640 50940 64070 50970
rect 63640 50920 63650 50940
rect 64070 50920 64130 50930
rect 67400 50990 67460 51000
rect 68140 50990 68150 51050
rect 68210 51030 68790 51050
rect 68210 50990 68220 51030
rect 73780 51080 73840 51090
rect 68790 51010 68850 51020
rect 73130 51050 73780 51060
rect 69060 50990 69120 51000
rect 67720 50980 67800 50990
rect 68140 50980 68220 50990
rect 68560 50980 68640 50990
rect 67720 50970 67730 50980
rect 67460 50940 67730 50970
rect 67400 50920 67460 50930
rect 67720 50920 67730 50940
rect 67790 50920 67800 50980
rect 63570 50910 63650 50920
rect 67720 50910 67800 50920
rect 68560 50920 68570 50980
rect 68630 50970 68640 50980
rect 68630 50940 69060 50970
rect 68630 50920 68640 50940
rect 69060 50920 69120 50930
rect 72510 50990 72570 51000
rect 73130 50990 73140 51050
rect 73200 51030 73780 51050
rect 73200 50990 73210 51030
rect 78770 51080 78830 51090
rect 73780 51010 73840 51020
rect 78120 51050 78770 51060
rect 73930 50990 73990 51000
rect 72710 50980 72790 50990
rect 73130 50980 73210 50990
rect 73550 50980 73630 50990
rect 72710 50970 72720 50980
rect 72570 50940 72720 50970
rect 72510 50920 72570 50930
rect 72710 50920 72720 50940
rect 72780 50920 72790 50980
rect 68560 50910 68640 50920
rect 72710 50910 72790 50920
rect 73550 50920 73560 50980
rect 73620 50970 73630 50980
rect 73620 50940 73930 50970
rect 73620 50920 73630 50940
rect 73930 50920 73990 50930
rect 77500 50990 77560 51000
rect 78120 50990 78130 51050
rect 78190 51030 78770 51050
rect 78190 50990 78200 51030
rect 78770 51010 78830 51020
rect 78920 50990 78980 51000
rect 77700 50980 77780 50990
rect 78120 50980 78200 50990
rect 78540 50980 78620 50990
rect 77700 50970 77710 50980
rect 77560 50940 77710 50970
rect 77500 50920 77560 50930
rect 77700 50920 77710 50940
rect 77770 50920 77780 50980
rect 73550 50910 73630 50920
rect 77700 50910 77780 50920
rect 78540 50920 78550 50980
rect 78610 50970 78620 50980
rect 78610 50940 78920 50970
rect 78610 50920 78620 50940
rect 78920 50920 78980 50930
rect 78540 50910 78620 50920
rect 53160 50890 53260 50900
rect 53160 50820 53180 50890
rect 53250 50820 53260 50890
rect 53160 50780 53260 50820
rect 53160 50710 53180 50780
rect 53250 50710 53260 50780
rect 53160 50690 53260 50710
rect 58150 50890 58250 50900
rect 58150 50820 58170 50890
rect 58240 50820 58250 50890
rect 58150 50780 58250 50820
rect 58150 50710 58170 50780
rect 58240 50710 58250 50780
rect 58150 50690 58250 50710
rect 63140 50890 63240 50900
rect 63140 50820 63160 50890
rect 63230 50820 63240 50890
rect 63140 50780 63240 50820
rect 63140 50710 63160 50780
rect 63230 50710 63240 50780
rect 63140 50690 63240 50710
rect 68130 50890 68230 50900
rect 68130 50820 68150 50890
rect 68220 50820 68230 50890
rect 68130 50780 68230 50820
rect 68130 50710 68150 50780
rect 68220 50710 68230 50780
rect 68130 50690 68230 50710
rect 73120 50890 73220 50900
rect 73120 50820 73140 50890
rect 73210 50820 73220 50890
rect 73120 50780 73220 50820
rect 73120 50710 73140 50780
rect 73210 50710 73220 50780
rect 73120 50690 73220 50710
rect 78110 50890 78210 50900
rect 78110 50820 78130 50890
rect 78200 50820 78210 50890
rect 78110 50780 78210 50820
rect 78110 50710 78130 50780
rect 78200 50710 78210 50780
rect 78110 50690 78210 50710
rect 52170 50670 52250 50680
rect 52170 50610 52180 50670
rect 52240 50660 52250 50670
rect 52750 50670 52830 50680
rect 52750 50660 52760 50670
rect 52240 50630 52760 50660
rect 52240 50610 52250 50630
rect 52170 50600 52250 50610
rect 52750 50610 52760 50630
rect 52820 50610 52830 50670
rect 53590 50670 53670 50680
rect 53590 50610 53600 50670
rect 53660 50660 53670 50670
rect 54330 50670 54410 50680
rect 54330 50660 54340 50670
rect 53660 50630 54340 50660
rect 53660 50610 53670 50630
rect 52750 50600 52830 50610
rect 53170 50600 53250 50610
rect 53590 50600 53670 50610
rect 54330 50610 54340 50630
rect 54400 50610 54410 50670
rect 54330 50600 54410 50610
rect 57160 50670 57240 50680
rect 57160 50610 57170 50670
rect 57230 50660 57240 50670
rect 57740 50670 57820 50680
rect 57740 50660 57750 50670
rect 57230 50630 57750 50660
rect 57230 50610 57240 50630
rect 57160 50600 57240 50610
rect 57740 50610 57750 50630
rect 57810 50610 57820 50670
rect 58580 50670 58660 50680
rect 58580 50610 58590 50670
rect 58650 50660 58660 50670
rect 59320 50670 59400 50680
rect 59320 50660 59330 50670
rect 58650 50630 59330 50660
rect 58650 50610 58660 50630
rect 57740 50600 57820 50610
rect 58160 50600 58240 50610
rect 58580 50600 58660 50610
rect 59320 50610 59330 50630
rect 59390 50610 59400 50670
rect 59320 50600 59400 50610
rect 62390 50670 62470 50680
rect 62390 50610 62400 50670
rect 62460 50660 62470 50670
rect 62730 50670 62810 50680
rect 62730 50660 62740 50670
rect 62460 50630 62740 50660
rect 62460 50610 62470 50630
rect 62390 50600 62470 50610
rect 62730 50610 62740 50630
rect 62800 50610 62810 50670
rect 63570 50670 63650 50680
rect 63570 50610 63580 50670
rect 63640 50660 63650 50670
rect 64070 50670 64150 50680
rect 64070 50660 64080 50670
rect 63640 50630 64080 50660
rect 63640 50610 63650 50630
rect 62730 50600 62810 50610
rect 63150 50600 63230 50610
rect 63570 50600 63650 50610
rect 64070 50610 64080 50630
rect 64140 50610 64150 50670
rect 64070 50600 64150 50610
rect 67380 50670 67460 50680
rect 67380 50610 67390 50670
rect 67450 50660 67460 50670
rect 67720 50670 67800 50680
rect 67720 50660 67730 50670
rect 67450 50630 67730 50660
rect 67450 50610 67460 50630
rect 67380 50600 67460 50610
rect 67720 50610 67730 50630
rect 67790 50610 67800 50670
rect 68560 50670 68640 50680
rect 68560 50610 68570 50670
rect 68630 50660 68640 50670
rect 69060 50670 69140 50680
rect 69060 50660 69070 50670
rect 68630 50630 69070 50660
rect 68630 50610 68640 50630
rect 67720 50600 67800 50610
rect 68140 50600 68220 50610
rect 68560 50600 68640 50610
rect 69060 50610 69070 50630
rect 69130 50610 69140 50670
rect 69060 50600 69140 50610
rect 72490 50670 72570 50680
rect 72490 50610 72500 50670
rect 72560 50660 72570 50670
rect 72710 50670 72790 50680
rect 72710 50660 72720 50670
rect 72560 50630 72720 50660
rect 72560 50610 72570 50630
rect 72490 50600 72570 50610
rect 72710 50610 72720 50630
rect 72780 50610 72790 50670
rect 73550 50670 73630 50680
rect 73550 50610 73560 50670
rect 73620 50660 73630 50670
rect 73930 50670 74010 50680
rect 73930 50660 73940 50670
rect 73620 50630 73940 50660
rect 73620 50610 73630 50630
rect 72710 50600 72790 50610
rect 73130 50600 73210 50610
rect 73550 50600 73630 50610
rect 73930 50610 73940 50630
rect 74000 50610 74010 50670
rect 73930 50600 74010 50610
rect 77480 50670 77560 50680
rect 77480 50610 77490 50670
rect 77550 50660 77560 50670
rect 77700 50670 77780 50680
rect 77700 50660 77710 50670
rect 77550 50630 77710 50660
rect 77550 50610 77560 50630
rect 77480 50600 77560 50610
rect 77700 50610 77710 50630
rect 77770 50610 77780 50670
rect 78540 50670 78620 50680
rect 78540 50610 78550 50670
rect 78610 50660 78620 50670
rect 78920 50670 79000 50680
rect 78920 50660 78930 50670
rect 78610 50630 78930 50660
rect 78610 50610 78620 50630
rect 77700 50600 77780 50610
rect 78120 50600 78200 50610
rect 78540 50600 78620 50610
rect 78920 50610 78930 50630
rect 78990 50610 79000 50670
rect 78920 50600 79000 50610
rect 53170 50540 53180 50600
rect 53240 50560 53250 50600
rect 53240 50550 53940 50560
rect 53240 50540 53880 50550
rect 53170 50530 53880 50540
rect 58160 50540 58170 50600
rect 58230 50560 58240 50600
rect 58230 50550 58930 50560
rect 58230 50540 58870 50550
rect 58160 50530 58870 50540
rect 53880 50480 53940 50490
rect 63150 50540 63160 50600
rect 63220 50560 63230 50600
rect 63220 50550 63920 50560
rect 63220 50540 63860 50550
rect 63150 50530 63860 50540
rect 58870 50480 58930 50490
rect 68140 50540 68150 50600
rect 68210 50560 68220 50600
rect 68210 50550 68910 50560
rect 68210 50540 68850 50550
rect 68140 50530 68850 50540
rect 63860 50480 63920 50490
rect 73130 50540 73140 50600
rect 73200 50560 73210 50600
rect 73200 50550 73900 50560
rect 73200 50540 73840 50550
rect 73130 50530 73840 50540
rect 68850 50480 68910 50490
rect 78120 50540 78130 50600
rect 78190 50560 78200 50600
rect 78190 50550 78890 50560
rect 78190 50540 78830 50550
rect 78120 50530 78830 50540
rect 73840 50480 73900 50490
rect 78830 50480 78890 50490
rect 53820 49370 53880 49380
rect 53170 49340 53820 49350
rect 52190 49280 52250 49290
rect 53170 49280 53180 49340
rect 53240 49320 53820 49340
rect 53240 49280 53250 49320
rect 58810 49370 58870 49380
rect 53820 49300 53880 49310
rect 58160 49340 58810 49350
rect 54330 49280 54390 49290
rect 52750 49270 52830 49280
rect 53170 49270 53250 49280
rect 53590 49270 53670 49280
rect 52750 49260 52760 49270
rect 52250 49230 52760 49260
rect 52190 49210 52250 49220
rect 52750 49210 52760 49230
rect 52820 49210 52830 49270
rect 52750 49200 52830 49210
rect 53590 49210 53600 49270
rect 53660 49260 53670 49270
rect 53660 49230 54330 49260
rect 53660 49210 53670 49230
rect 54330 49210 54390 49220
rect 57180 49280 57240 49290
rect 58160 49280 58170 49340
rect 58230 49320 58810 49340
rect 58230 49280 58240 49320
rect 63800 49370 63860 49380
rect 58810 49300 58870 49310
rect 63150 49340 63800 49350
rect 59320 49280 59380 49290
rect 57740 49270 57820 49280
rect 58160 49270 58240 49280
rect 58580 49270 58660 49280
rect 57740 49260 57750 49270
rect 57240 49230 57750 49260
rect 57180 49210 57240 49220
rect 57740 49210 57750 49230
rect 57810 49210 57820 49270
rect 53590 49200 53670 49210
rect 57740 49200 57820 49210
rect 58580 49210 58590 49270
rect 58650 49260 58660 49270
rect 58650 49230 59320 49260
rect 58650 49210 58660 49230
rect 59320 49210 59380 49220
rect 62410 49280 62470 49290
rect 63150 49280 63160 49340
rect 63220 49320 63800 49340
rect 63220 49280 63230 49320
rect 68790 49370 68850 49380
rect 63800 49300 63860 49310
rect 68140 49340 68790 49350
rect 64070 49280 64130 49290
rect 62730 49270 62810 49280
rect 63150 49270 63230 49280
rect 63570 49270 63650 49280
rect 62730 49260 62740 49270
rect 62470 49230 62740 49260
rect 62410 49210 62470 49220
rect 62730 49210 62740 49230
rect 62800 49210 62810 49270
rect 58580 49200 58660 49210
rect 62730 49200 62810 49210
rect 63570 49210 63580 49270
rect 63640 49260 63650 49270
rect 63640 49230 64070 49260
rect 63640 49210 63650 49230
rect 64070 49210 64130 49220
rect 67400 49280 67460 49290
rect 68140 49280 68150 49340
rect 68210 49320 68790 49340
rect 68210 49280 68220 49320
rect 73780 49370 73840 49380
rect 68790 49300 68850 49310
rect 73130 49340 73780 49350
rect 69060 49280 69120 49290
rect 67720 49270 67800 49280
rect 68140 49270 68220 49280
rect 68560 49270 68640 49280
rect 67720 49260 67730 49270
rect 67460 49230 67730 49260
rect 67400 49210 67460 49220
rect 67720 49210 67730 49230
rect 67790 49210 67800 49270
rect 63570 49200 63650 49210
rect 67720 49200 67800 49210
rect 68560 49210 68570 49270
rect 68630 49260 68640 49270
rect 68630 49230 69060 49260
rect 68630 49210 68640 49230
rect 69060 49210 69120 49220
rect 72510 49280 72570 49290
rect 73130 49280 73140 49340
rect 73200 49320 73780 49340
rect 73200 49280 73210 49320
rect 78770 49370 78830 49380
rect 73780 49300 73840 49310
rect 78120 49340 78770 49350
rect 73930 49280 73990 49290
rect 72710 49270 72790 49280
rect 73130 49270 73210 49280
rect 73550 49270 73630 49280
rect 72710 49260 72720 49270
rect 72570 49230 72720 49260
rect 72510 49210 72570 49220
rect 72710 49210 72720 49230
rect 72780 49210 72790 49270
rect 68560 49200 68640 49210
rect 72710 49200 72790 49210
rect 73550 49210 73560 49270
rect 73620 49260 73630 49270
rect 73620 49230 73930 49260
rect 73620 49210 73630 49230
rect 73930 49210 73990 49220
rect 77500 49280 77560 49290
rect 78120 49280 78130 49340
rect 78190 49320 78770 49340
rect 78190 49280 78200 49320
rect 78770 49300 78830 49310
rect 78920 49280 78980 49290
rect 77700 49270 77780 49280
rect 78120 49270 78200 49280
rect 78540 49270 78620 49280
rect 77700 49260 77710 49270
rect 77560 49230 77710 49260
rect 77500 49210 77560 49220
rect 77700 49210 77710 49230
rect 77770 49210 77780 49270
rect 73550 49200 73630 49210
rect 77700 49200 77780 49210
rect 78540 49210 78550 49270
rect 78610 49260 78620 49270
rect 78610 49230 78920 49260
rect 78610 49210 78620 49230
rect 78920 49210 78980 49220
rect 78540 49200 78620 49210
rect 53160 49180 53260 49190
rect 53160 49110 53180 49180
rect 53250 49110 53260 49180
rect 53160 49070 53260 49110
rect 53160 49000 53180 49070
rect 53250 49000 53260 49070
rect 53160 48980 53260 49000
rect 58150 49180 58250 49190
rect 58150 49110 58170 49180
rect 58240 49110 58250 49180
rect 58150 49070 58250 49110
rect 58150 49000 58170 49070
rect 58240 49000 58250 49070
rect 58150 48980 58250 49000
rect 63140 49180 63240 49190
rect 63140 49110 63160 49180
rect 63230 49110 63240 49180
rect 63140 49070 63240 49110
rect 63140 49000 63160 49070
rect 63230 49000 63240 49070
rect 63140 48980 63240 49000
rect 68130 49180 68230 49190
rect 68130 49110 68150 49180
rect 68220 49110 68230 49180
rect 68130 49070 68230 49110
rect 68130 49000 68150 49070
rect 68220 49000 68230 49070
rect 68130 48980 68230 49000
rect 73120 49180 73220 49190
rect 73120 49110 73140 49180
rect 73210 49110 73220 49180
rect 73120 49070 73220 49110
rect 73120 49000 73140 49070
rect 73210 49000 73220 49070
rect 73120 48980 73220 49000
rect 78110 49180 78210 49190
rect 78110 49110 78130 49180
rect 78200 49110 78210 49180
rect 78110 49070 78210 49110
rect 78110 49000 78130 49070
rect 78200 49000 78210 49070
rect 78110 48980 78210 49000
rect 52170 48960 52250 48970
rect 52170 48900 52180 48960
rect 52240 48950 52250 48960
rect 52750 48960 52830 48970
rect 52750 48950 52760 48960
rect 52240 48920 52760 48950
rect 52240 48900 52250 48920
rect 52170 48890 52250 48900
rect 52750 48900 52760 48920
rect 52820 48900 52830 48960
rect 53590 48960 53670 48970
rect 53590 48900 53600 48960
rect 53660 48950 53670 48960
rect 54330 48960 54410 48970
rect 54330 48950 54340 48960
rect 53660 48920 54340 48950
rect 53660 48900 53670 48920
rect 52750 48890 52830 48900
rect 53170 48890 53250 48900
rect 53590 48890 53670 48900
rect 54330 48900 54340 48920
rect 54400 48900 54410 48960
rect 54330 48890 54410 48900
rect 57160 48960 57240 48970
rect 57160 48900 57170 48960
rect 57230 48950 57240 48960
rect 57740 48960 57820 48970
rect 57740 48950 57750 48960
rect 57230 48920 57750 48950
rect 57230 48900 57240 48920
rect 57160 48890 57240 48900
rect 57740 48900 57750 48920
rect 57810 48900 57820 48960
rect 58580 48960 58660 48970
rect 58580 48900 58590 48960
rect 58650 48950 58660 48960
rect 59320 48960 59400 48970
rect 59320 48950 59330 48960
rect 58650 48920 59330 48950
rect 58650 48900 58660 48920
rect 57740 48890 57820 48900
rect 58160 48890 58240 48900
rect 58580 48890 58660 48900
rect 59320 48900 59330 48920
rect 59390 48900 59400 48960
rect 59320 48890 59400 48900
rect 62390 48960 62470 48970
rect 62390 48900 62400 48960
rect 62460 48950 62470 48960
rect 62730 48960 62810 48970
rect 62730 48950 62740 48960
rect 62460 48920 62740 48950
rect 62460 48900 62470 48920
rect 62390 48890 62470 48900
rect 62730 48900 62740 48920
rect 62800 48900 62810 48960
rect 63570 48960 63650 48970
rect 63570 48900 63580 48960
rect 63640 48950 63650 48960
rect 64070 48960 64150 48970
rect 64070 48950 64080 48960
rect 63640 48920 64080 48950
rect 63640 48900 63650 48920
rect 62730 48890 62810 48900
rect 63150 48890 63230 48900
rect 63570 48890 63650 48900
rect 64070 48900 64080 48920
rect 64140 48900 64150 48960
rect 64070 48890 64150 48900
rect 67380 48960 67460 48970
rect 67380 48900 67390 48960
rect 67450 48950 67460 48960
rect 67720 48960 67800 48970
rect 67720 48950 67730 48960
rect 67450 48920 67730 48950
rect 67450 48900 67460 48920
rect 67380 48890 67460 48900
rect 67720 48900 67730 48920
rect 67790 48900 67800 48960
rect 68560 48960 68640 48970
rect 68560 48900 68570 48960
rect 68630 48950 68640 48960
rect 69060 48960 69140 48970
rect 69060 48950 69070 48960
rect 68630 48920 69070 48950
rect 68630 48900 68640 48920
rect 67720 48890 67800 48900
rect 68140 48890 68220 48900
rect 68560 48890 68640 48900
rect 69060 48900 69070 48920
rect 69130 48900 69140 48960
rect 69060 48890 69140 48900
rect 72490 48960 72570 48970
rect 72490 48900 72500 48960
rect 72560 48950 72570 48960
rect 72710 48960 72790 48970
rect 72710 48950 72720 48960
rect 72560 48920 72720 48950
rect 72560 48900 72570 48920
rect 72490 48890 72570 48900
rect 72710 48900 72720 48920
rect 72780 48900 72790 48960
rect 73550 48960 73630 48970
rect 73550 48900 73560 48960
rect 73620 48950 73630 48960
rect 73930 48960 74010 48970
rect 73930 48950 73940 48960
rect 73620 48920 73940 48950
rect 73620 48900 73630 48920
rect 72710 48890 72790 48900
rect 73130 48890 73210 48900
rect 73550 48890 73630 48900
rect 73930 48900 73940 48920
rect 74000 48900 74010 48960
rect 73930 48890 74010 48900
rect 77480 48960 77560 48970
rect 77480 48900 77490 48960
rect 77550 48950 77560 48960
rect 77700 48960 77780 48970
rect 77700 48950 77710 48960
rect 77550 48920 77710 48950
rect 77550 48900 77560 48920
rect 77480 48890 77560 48900
rect 77700 48900 77710 48920
rect 77770 48900 77780 48960
rect 78540 48960 78620 48970
rect 78540 48900 78550 48960
rect 78610 48950 78620 48960
rect 78920 48960 79000 48970
rect 78920 48950 78930 48960
rect 78610 48920 78930 48950
rect 78610 48900 78620 48920
rect 77700 48890 77780 48900
rect 78120 48890 78200 48900
rect 78540 48890 78620 48900
rect 78920 48900 78930 48920
rect 78990 48900 79000 48960
rect 78920 48890 79000 48900
rect 49580 39510 50050 39540
rect 49460 39450 49870 39480
rect 49340 39390 49690 39420
rect 49220 39330 49510 39360
rect 49100 39270 49330 39300
rect 48980 39210 49150 39240
rect 48720 38690 48800 38700
rect 48720 38630 48730 38690
rect 48790 38630 48800 38690
rect 48870 38640 48880 38700
rect 48940 38640 48950 38700
rect 48720 38620 48800 38630
rect 49120 36320 49150 39210
rect 49180 39230 49240 39240
rect 49180 39160 49240 39170
rect 47420 36310 47500 36320
rect 47420 36250 47430 36310
rect 47490 36250 47500 36310
rect 49100 36260 49110 36320
rect 49170 36260 49180 36320
rect 47420 36240 47500 36250
rect 49210 36180 49240 39160
rect 49300 36600 49330 39270
rect 49360 39290 49420 39300
rect 49360 39220 49420 39230
rect 49280 36540 49290 36600
rect 49350 36540 49360 36600
rect 49390 36460 49420 39220
rect 49480 36880 49510 39330
rect 49540 39350 49600 39360
rect 49540 39280 49600 39290
rect 49460 36820 49470 36880
rect 49530 36820 49540 36880
rect 49570 36740 49600 39280
rect 49660 37160 49690 39390
rect 49720 39410 49780 39420
rect 49720 39340 49780 39350
rect 49640 37100 49650 37160
rect 49710 37100 49720 37160
rect 49750 37020 49780 39340
rect 49840 37720 49870 39450
rect 49900 39470 49960 39480
rect 49900 39400 49960 39410
rect 49820 37660 49830 37720
rect 49890 37660 49900 37720
rect 49930 37580 49960 39400
rect 49880 37520 49890 37580
rect 49950 37520 49960 37580
rect 50020 37440 50050 39510
rect 50080 39530 50140 39540
rect 50080 39460 50140 39470
rect 50000 37380 50010 37440
rect 50070 37380 50080 37440
rect 50110 37300 50140 39460
rect 52220 39420 52250 48890
rect 53170 48830 53180 48890
rect 53240 48850 53250 48890
rect 53240 48840 53940 48850
rect 53240 48830 53880 48840
rect 53170 48820 53880 48830
rect 53880 48770 53940 48780
rect 53820 47660 53880 47670
rect 53170 47630 53820 47640
rect 52310 47570 52370 47580
rect 53170 47570 53180 47630
rect 53240 47610 53820 47630
rect 53240 47570 53250 47610
rect 53820 47590 53880 47600
rect 54210 47570 54270 47580
rect 52750 47560 52830 47570
rect 53170 47560 53250 47570
rect 53590 47560 53670 47570
rect 52750 47550 52760 47560
rect 52370 47520 52760 47550
rect 52310 47500 52370 47510
rect 52750 47500 52760 47520
rect 52820 47500 52830 47560
rect 52750 47490 52830 47500
rect 53590 47500 53600 47560
rect 53660 47550 53670 47560
rect 53660 47520 54210 47550
rect 53660 47500 53670 47520
rect 54210 47500 54270 47510
rect 53590 47490 53670 47500
rect 53160 47470 53260 47480
rect 53160 47400 53180 47470
rect 53250 47400 53260 47470
rect 53160 47360 53260 47400
rect 53160 47290 53180 47360
rect 53250 47290 53260 47360
rect 53160 47270 53260 47290
rect 52290 47250 52370 47260
rect 52290 47190 52300 47250
rect 52360 47240 52370 47250
rect 52750 47250 52830 47260
rect 52750 47240 52760 47250
rect 52360 47210 52760 47240
rect 52360 47190 52370 47210
rect 52290 47180 52370 47190
rect 52750 47190 52760 47210
rect 52820 47190 52830 47250
rect 53590 47250 53670 47260
rect 53590 47190 53600 47250
rect 53660 47240 53670 47250
rect 54210 47250 54290 47260
rect 54210 47240 54220 47250
rect 53660 47210 54220 47240
rect 53660 47190 53670 47210
rect 52750 47180 52830 47190
rect 53170 47180 53250 47190
rect 53590 47180 53670 47190
rect 54210 47190 54220 47210
rect 54280 47190 54290 47250
rect 54210 47180 54290 47190
rect 50060 37240 50070 37300
rect 50130 37240 50140 37300
rect 51810 39410 51870 39420
rect 51810 39340 51870 39350
rect 51900 39390 52250 39420
rect 49700 36960 49710 37020
rect 49770 36960 49780 37020
rect 49520 36680 49530 36740
rect 49590 36680 49600 36740
rect 51810 36740 51840 39340
rect 51900 36880 51930 39390
rect 52340 39360 52370 47180
rect 53170 47120 53180 47180
rect 53240 47140 53250 47180
rect 53240 47130 53940 47140
rect 53240 47120 53880 47130
rect 53170 47110 53880 47120
rect 53880 47060 53940 47070
rect 53820 45950 53880 45960
rect 53170 45920 53820 45930
rect 52430 45860 52490 45870
rect 53170 45860 53180 45920
rect 53240 45900 53820 45920
rect 53240 45860 53250 45900
rect 53820 45880 53880 45890
rect 54090 45860 54150 45870
rect 52750 45850 52830 45860
rect 53170 45850 53250 45860
rect 53590 45850 53670 45860
rect 52750 45840 52760 45850
rect 52490 45810 52760 45840
rect 52430 45790 52490 45800
rect 52750 45790 52760 45810
rect 52820 45790 52830 45850
rect 52750 45780 52830 45790
rect 53590 45790 53600 45850
rect 53660 45840 53670 45850
rect 53660 45810 54090 45840
rect 53660 45790 53670 45810
rect 54090 45790 54150 45800
rect 53590 45780 53670 45790
rect 53160 45760 53260 45770
rect 53160 45690 53180 45760
rect 53250 45690 53260 45760
rect 53160 45650 53260 45690
rect 53160 45580 53180 45650
rect 53250 45580 53260 45650
rect 53160 45560 53260 45580
rect 52410 45540 52490 45550
rect 52410 45480 52420 45540
rect 52480 45530 52490 45540
rect 52750 45540 52830 45550
rect 52750 45530 52760 45540
rect 52480 45500 52760 45530
rect 52480 45480 52490 45500
rect 52410 45470 52490 45480
rect 52750 45480 52760 45500
rect 52820 45480 52830 45540
rect 53590 45540 53670 45550
rect 53590 45480 53600 45540
rect 53660 45530 53670 45540
rect 54090 45540 54170 45550
rect 54090 45530 54100 45540
rect 53660 45500 54100 45530
rect 53660 45480 53670 45500
rect 52750 45470 52830 45480
rect 53170 45470 53250 45480
rect 53590 45470 53670 45480
rect 54090 45480 54100 45500
rect 54160 45480 54170 45540
rect 54090 45470 54170 45480
rect 53170 45410 53180 45470
rect 53240 45430 53250 45470
rect 53240 45420 53940 45430
rect 53240 45410 53880 45420
rect 53170 45400 53880 45410
rect 53880 45350 53940 45360
rect 53820 44240 53880 44250
rect 53170 44210 53820 44220
rect 52430 44150 52490 44160
rect 53170 44150 53180 44210
rect 53240 44190 53820 44210
rect 53240 44150 53250 44190
rect 53820 44170 53880 44180
rect 54090 44150 54150 44160
rect 52750 44140 52830 44150
rect 53170 44140 53250 44150
rect 53590 44140 53670 44150
rect 52750 44130 52760 44140
rect 52490 44100 52760 44130
rect 52430 44080 52490 44090
rect 52750 44080 52760 44100
rect 52820 44080 52830 44140
rect 52750 44070 52830 44080
rect 53590 44080 53600 44140
rect 53660 44130 53670 44140
rect 53660 44100 54090 44130
rect 53660 44080 53670 44100
rect 54090 44080 54150 44090
rect 53590 44070 53670 44080
rect 53160 44050 53260 44060
rect 53160 43980 53180 44050
rect 53250 43980 53260 44050
rect 53160 43940 53260 43980
rect 53160 43870 53180 43940
rect 53250 43870 53260 43940
rect 53160 43850 53260 43870
rect 52410 43830 52490 43840
rect 52410 43770 52420 43830
rect 52480 43820 52490 43830
rect 52750 43830 52830 43840
rect 52750 43820 52760 43830
rect 52480 43790 52760 43820
rect 52480 43770 52490 43790
rect 52410 43760 52490 43770
rect 52750 43770 52760 43790
rect 52820 43770 52830 43830
rect 53590 43830 53670 43840
rect 53590 43770 53600 43830
rect 53660 43820 53670 43830
rect 54090 43830 54170 43840
rect 54090 43820 54100 43830
rect 53660 43790 54100 43820
rect 53660 43770 53670 43790
rect 52750 43760 52830 43770
rect 53170 43760 53250 43770
rect 53590 43760 53670 43770
rect 54090 43770 54100 43790
rect 54160 43770 54170 43830
rect 54090 43760 54170 43770
rect 51990 39350 52050 39360
rect 51990 39280 52050 39290
rect 52080 39330 52370 39360
rect 51990 37020 52020 39280
rect 52080 37160 52110 39330
rect 52460 39300 52490 43760
rect 53170 43700 53180 43760
rect 53240 43720 53250 43760
rect 53240 43710 53940 43720
rect 53240 43700 53880 43710
rect 53170 43690 53880 43700
rect 53880 43640 53940 43650
rect 53820 42530 53880 42540
rect 53170 42500 53820 42510
rect 52550 42440 52610 42450
rect 53170 42440 53180 42500
rect 53240 42480 53820 42500
rect 53240 42440 53250 42480
rect 53820 42460 53880 42470
rect 53970 42440 54030 42450
rect 52750 42430 52830 42440
rect 53170 42430 53250 42440
rect 53590 42430 53670 42440
rect 52750 42420 52760 42430
rect 52610 42390 52760 42420
rect 52550 42370 52610 42380
rect 52750 42370 52760 42390
rect 52820 42370 52830 42430
rect 52750 42360 52830 42370
rect 53590 42370 53600 42430
rect 53660 42420 53670 42430
rect 53660 42390 53970 42420
rect 53660 42370 53670 42390
rect 53970 42370 54030 42380
rect 53590 42360 53670 42370
rect 53160 42340 53260 42350
rect 53160 42270 53180 42340
rect 53250 42270 53260 42340
rect 53160 42230 53260 42270
rect 53160 42160 53180 42230
rect 53250 42160 53260 42230
rect 53160 42140 53260 42160
rect 52530 42120 52610 42130
rect 52530 42060 52540 42120
rect 52600 42110 52610 42120
rect 52750 42120 52830 42130
rect 52750 42110 52760 42120
rect 52600 42080 52760 42110
rect 52600 42060 52610 42080
rect 52530 42050 52610 42060
rect 52750 42060 52760 42080
rect 52820 42060 52830 42120
rect 53590 42120 53670 42130
rect 53590 42060 53600 42120
rect 53660 42110 53670 42120
rect 53970 42120 54050 42130
rect 53970 42110 53980 42120
rect 53660 42080 53980 42110
rect 53660 42060 53670 42080
rect 52750 42050 52830 42060
rect 53170 42050 53250 42060
rect 53590 42050 53670 42060
rect 53970 42060 53980 42080
rect 54040 42060 54050 42120
rect 53970 42050 54050 42060
rect 53170 41990 53180 42050
rect 53240 42010 53250 42050
rect 53240 42000 53940 42010
rect 53240 41990 53880 42000
rect 53170 41980 53880 41990
rect 53880 41930 53940 41940
rect 53820 40820 53880 40830
rect 53170 40790 53820 40800
rect 52550 40730 52610 40740
rect 53170 40730 53180 40790
rect 53240 40770 53820 40790
rect 53240 40730 53250 40770
rect 53820 40750 53880 40760
rect 53970 40730 54030 40740
rect 52750 40720 52830 40730
rect 53170 40720 53250 40730
rect 53590 40720 53670 40730
rect 52750 40710 52760 40720
rect 52610 40680 52760 40710
rect 52550 40660 52610 40670
rect 52750 40660 52760 40680
rect 52820 40660 52830 40720
rect 52750 40650 52830 40660
rect 53590 40660 53600 40720
rect 53660 40710 53670 40720
rect 53660 40680 53970 40710
rect 53660 40660 53670 40680
rect 53970 40660 54030 40670
rect 53590 40650 53670 40660
rect 53160 40630 53260 40640
rect 53160 40560 53180 40630
rect 53250 40560 53260 40630
rect 53160 40520 53260 40560
rect 53160 40450 53180 40520
rect 53250 40450 53260 40520
rect 53160 40430 53260 40450
rect 52530 40410 52610 40420
rect 52530 40350 52540 40410
rect 52600 40400 52610 40410
rect 52750 40410 52830 40420
rect 52750 40400 52760 40410
rect 52600 40370 52760 40400
rect 52600 40350 52610 40370
rect 52530 40340 52610 40350
rect 52750 40350 52760 40370
rect 52820 40350 52830 40410
rect 53590 40410 53670 40420
rect 53590 40350 53600 40410
rect 53660 40400 53670 40410
rect 53970 40410 54050 40420
rect 53970 40400 53980 40410
rect 53660 40370 53980 40400
rect 53660 40350 53670 40370
rect 52750 40340 52830 40350
rect 53170 40340 53250 40350
rect 53590 40340 53670 40350
rect 53970 40350 53980 40370
rect 54040 40350 54050 40410
rect 53970 40340 54050 40350
rect 52170 39290 52230 39300
rect 52170 39220 52230 39230
rect 52260 39270 52490 39300
rect 52050 37150 52130 37160
rect 52050 37090 52060 37150
rect 52120 37090 52130 37150
rect 52050 37080 52130 37090
rect 51990 37010 52070 37020
rect 51990 36950 52000 37010
rect 52060 36950 52070 37010
rect 51990 36940 52070 36950
rect 51870 36870 51950 36880
rect 51870 36810 51880 36870
rect 51940 36810 51950 36870
rect 51870 36800 51950 36810
rect 51810 36730 51890 36740
rect 51810 36670 51820 36730
rect 51880 36670 51890 36730
rect 51810 36660 51890 36670
rect 49340 36400 49350 36460
rect 49410 36400 49420 36460
rect 52170 36460 52200 39220
rect 52260 36600 52290 39270
rect 52580 39240 52610 40340
rect 53170 40280 53180 40340
rect 53240 40300 53250 40340
rect 53240 40290 53940 40300
rect 53240 40280 53880 40290
rect 53170 40270 53880 40280
rect 53880 40220 53940 40230
rect 52350 39230 52410 39240
rect 52350 39160 52410 39170
rect 52440 39210 52610 39240
rect 52640 39680 52720 39690
rect 52640 39620 52650 39680
rect 52710 39620 52720 39680
rect 53710 39680 53790 39690
rect 53710 39620 53720 39680
rect 53780 39620 53790 39680
rect 52230 36590 52310 36600
rect 52230 36530 52240 36590
rect 52300 36530 52310 36590
rect 52230 36520 52310 36530
rect 52170 36450 52250 36460
rect 52170 36390 52180 36450
rect 52240 36390 52250 36450
rect 52170 36380 52250 36390
rect 47360 36170 47440 36180
rect 42370 36100 42450 36110
rect 47360 36110 47370 36170
rect 47430 36110 47440 36170
rect 49160 36120 49170 36180
rect 49230 36120 49240 36180
rect 52350 36180 52380 39160
rect 52440 36320 52470 39210
rect 52640 38840 52710 39620
rect 53710 39610 53790 39620
rect 53880 39680 53940 39690
rect 53880 39610 53940 39620
rect 52640 38830 52720 38840
rect 52640 38770 52650 38830
rect 52710 38770 52720 38830
rect 52640 38760 52720 38770
rect 53720 38700 53790 39610
rect 53910 38700 53940 39610
rect 53970 39240 54000 40340
rect 54090 39300 54120 43760
rect 54210 39360 54240 47180
rect 54330 39420 54360 48890
rect 57210 39420 57240 48890
rect 58160 48830 58170 48890
rect 58230 48850 58240 48890
rect 58230 48840 58930 48850
rect 58230 48830 58870 48840
rect 58160 48820 58870 48830
rect 58870 48770 58930 48780
rect 58810 47660 58870 47670
rect 58160 47630 58810 47640
rect 57300 47570 57360 47580
rect 58160 47570 58170 47630
rect 58230 47610 58810 47630
rect 58230 47570 58240 47610
rect 58810 47590 58870 47600
rect 59200 47570 59260 47580
rect 57740 47560 57820 47570
rect 58160 47560 58240 47570
rect 58580 47560 58660 47570
rect 57740 47550 57750 47560
rect 57360 47520 57750 47550
rect 57300 47500 57360 47510
rect 57740 47500 57750 47520
rect 57810 47500 57820 47560
rect 57740 47490 57820 47500
rect 58580 47500 58590 47560
rect 58650 47550 58660 47560
rect 58650 47520 59200 47550
rect 58650 47500 58660 47520
rect 59200 47500 59260 47510
rect 58580 47490 58660 47500
rect 58150 47470 58250 47480
rect 58150 47400 58170 47470
rect 58240 47400 58250 47470
rect 58150 47360 58250 47400
rect 58150 47290 58170 47360
rect 58240 47290 58250 47360
rect 58150 47270 58250 47290
rect 57280 47250 57360 47260
rect 57280 47190 57290 47250
rect 57350 47240 57360 47250
rect 57740 47250 57820 47260
rect 57740 47240 57750 47250
rect 57350 47210 57750 47240
rect 57350 47190 57360 47210
rect 57280 47180 57360 47190
rect 57740 47190 57750 47210
rect 57810 47190 57820 47250
rect 58580 47250 58660 47260
rect 58580 47190 58590 47250
rect 58650 47240 58660 47250
rect 59200 47250 59280 47260
rect 59200 47240 59210 47250
rect 58650 47210 59210 47240
rect 58650 47190 58660 47210
rect 57740 47180 57820 47190
rect 58160 47180 58240 47190
rect 58580 47180 58660 47190
rect 59200 47190 59210 47210
rect 59270 47190 59280 47250
rect 59200 47180 59280 47190
rect 54330 39390 54680 39420
rect 54210 39330 54500 39360
rect 54090 39270 54320 39300
rect 53970 39210 54140 39240
rect 53710 38690 53790 38700
rect 53710 38630 53720 38690
rect 53780 38630 53790 38690
rect 53860 38640 53870 38700
rect 53930 38640 53940 38700
rect 53710 38620 53790 38630
rect 54110 36320 54140 39210
rect 54170 39230 54230 39240
rect 54170 39160 54230 39170
rect 52410 36310 52490 36320
rect 52410 36250 52420 36310
rect 52480 36250 52490 36310
rect 54090 36260 54100 36320
rect 54160 36260 54170 36320
rect 52410 36240 52490 36250
rect 54200 36180 54230 39160
rect 54290 36600 54320 39270
rect 54350 39290 54410 39300
rect 54350 39220 54410 39230
rect 54270 36540 54280 36600
rect 54340 36540 54350 36600
rect 54380 36460 54410 39220
rect 54470 37160 54500 39330
rect 54530 39350 54590 39360
rect 54530 39280 54590 39290
rect 54450 37100 54460 37160
rect 54520 37100 54530 37160
rect 54560 37020 54590 39280
rect 54510 36960 54520 37020
rect 54580 36960 54590 37020
rect 54650 36880 54680 39390
rect 54710 39410 54770 39420
rect 54710 39340 54770 39350
rect 54630 36820 54640 36880
rect 54700 36820 54710 36880
rect 54740 36740 54770 39340
rect 54690 36680 54700 36740
rect 54760 36680 54770 36740
rect 56800 39410 56860 39420
rect 56800 39340 56860 39350
rect 56890 39390 57240 39420
rect 56800 36740 56830 39340
rect 56890 36880 56920 39390
rect 57330 39360 57360 47180
rect 58160 47120 58170 47180
rect 58230 47140 58240 47180
rect 58230 47130 58930 47140
rect 58230 47120 58870 47130
rect 58160 47110 58870 47120
rect 58870 47060 58930 47070
rect 58810 45950 58870 45960
rect 58160 45920 58810 45930
rect 57420 45860 57480 45870
rect 58160 45860 58170 45920
rect 58230 45900 58810 45920
rect 58230 45860 58240 45900
rect 58810 45880 58870 45890
rect 59080 45860 59140 45870
rect 57740 45850 57820 45860
rect 58160 45850 58240 45860
rect 58580 45850 58660 45860
rect 57740 45840 57750 45850
rect 57480 45810 57750 45840
rect 57420 45790 57480 45800
rect 57740 45790 57750 45810
rect 57810 45790 57820 45850
rect 57740 45780 57820 45790
rect 58580 45790 58590 45850
rect 58650 45840 58660 45850
rect 58650 45810 59080 45840
rect 58650 45790 58660 45810
rect 59080 45790 59140 45800
rect 58580 45780 58660 45790
rect 58150 45760 58250 45770
rect 58150 45690 58170 45760
rect 58240 45690 58250 45760
rect 58150 45650 58250 45690
rect 58150 45580 58170 45650
rect 58240 45580 58250 45650
rect 58150 45560 58250 45580
rect 57400 45540 57480 45550
rect 57400 45480 57410 45540
rect 57470 45530 57480 45540
rect 57740 45540 57820 45550
rect 57740 45530 57750 45540
rect 57470 45500 57750 45530
rect 57470 45480 57480 45500
rect 57400 45470 57480 45480
rect 57740 45480 57750 45500
rect 57810 45480 57820 45540
rect 58580 45540 58660 45550
rect 58580 45480 58590 45540
rect 58650 45530 58660 45540
rect 59080 45540 59160 45550
rect 59080 45530 59090 45540
rect 58650 45500 59090 45530
rect 58650 45480 58660 45500
rect 57740 45470 57820 45480
rect 58160 45470 58240 45480
rect 58580 45470 58660 45480
rect 59080 45480 59090 45500
rect 59150 45480 59160 45540
rect 59080 45470 59160 45480
rect 58160 45410 58170 45470
rect 58230 45430 58240 45470
rect 58230 45420 58930 45430
rect 58230 45410 58870 45420
rect 58160 45400 58870 45410
rect 58870 45350 58930 45360
rect 58810 44240 58870 44250
rect 58160 44210 58810 44220
rect 57420 44150 57480 44160
rect 58160 44150 58170 44210
rect 58230 44190 58810 44210
rect 58230 44150 58240 44190
rect 58810 44170 58870 44180
rect 59080 44150 59140 44160
rect 57740 44140 57820 44150
rect 58160 44140 58240 44150
rect 58580 44140 58660 44150
rect 57740 44130 57750 44140
rect 57480 44100 57750 44130
rect 57420 44080 57480 44090
rect 57740 44080 57750 44100
rect 57810 44080 57820 44140
rect 57740 44070 57820 44080
rect 58580 44080 58590 44140
rect 58650 44130 58660 44140
rect 58650 44100 59080 44130
rect 58650 44080 58660 44100
rect 59080 44080 59140 44090
rect 58580 44070 58660 44080
rect 58150 44050 58250 44060
rect 58150 43980 58170 44050
rect 58240 43980 58250 44050
rect 58150 43940 58250 43980
rect 58150 43870 58170 43940
rect 58240 43870 58250 43940
rect 58150 43850 58250 43870
rect 57400 43830 57480 43840
rect 57400 43770 57410 43830
rect 57470 43820 57480 43830
rect 57740 43830 57820 43840
rect 57740 43820 57750 43830
rect 57470 43790 57750 43820
rect 57470 43770 57480 43790
rect 57400 43760 57480 43770
rect 57740 43770 57750 43790
rect 57810 43770 57820 43830
rect 58580 43830 58660 43840
rect 58580 43770 58590 43830
rect 58650 43820 58660 43830
rect 59080 43830 59160 43840
rect 59080 43820 59090 43830
rect 58650 43790 59090 43820
rect 58650 43770 58660 43790
rect 57740 43760 57820 43770
rect 58160 43760 58240 43770
rect 58580 43760 58660 43770
rect 59080 43770 59090 43790
rect 59150 43770 59160 43830
rect 59080 43760 59160 43770
rect 56980 39350 57040 39360
rect 56980 39280 57040 39290
rect 57070 39330 57360 39360
rect 56980 37020 57010 39280
rect 57070 37160 57100 39330
rect 57450 39300 57480 43760
rect 58160 43700 58170 43760
rect 58230 43720 58240 43760
rect 58230 43710 58930 43720
rect 58230 43700 58870 43710
rect 58160 43690 58870 43700
rect 58870 43640 58930 43650
rect 58810 42530 58870 42540
rect 58160 42500 58810 42510
rect 57540 42440 57600 42450
rect 58160 42440 58170 42500
rect 58230 42480 58810 42500
rect 58230 42440 58240 42480
rect 58810 42460 58870 42470
rect 58960 42440 59020 42450
rect 57740 42430 57820 42440
rect 58160 42430 58240 42440
rect 58580 42430 58660 42440
rect 57740 42420 57750 42430
rect 57600 42390 57750 42420
rect 57540 42370 57600 42380
rect 57740 42370 57750 42390
rect 57810 42370 57820 42430
rect 57740 42360 57820 42370
rect 58580 42370 58590 42430
rect 58650 42420 58660 42430
rect 58650 42390 58960 42420
rect 58650 42370 58660 42390
rect 58960 42370 59020 42380
rect 58580 42360 58660 42370
rect 58150 42340 58250 42350
rect 58150 42270 58170 42340
rect 58240 42270 58250 42340
rect 58150 42230 58250 42270
rect 58150 42160 58170 42230
rect 58240 42160 58250 42230
rect 58150 42140 58250 42160
rect 57520 42120 57600 42130
rect 57520 42060 57530 42120
rect 57590 42110 57600 42120
rect 57740 42120 57820 42130
rect 57740 42110 57750 42120
rect 57590 42080 57750 42110
rect 57590 42060 57600 42080
rect 57520 42050 57600 42060
rect 57740 42060 57750 42080
rect 57810 42060 57820 42120
rect 58580 42120 58660 42130
rect 58580 42060 58590 42120
rect 58650 42110 58660 42120
rect 58960 42120 59040 42130
rect 58960 42110 58970 42120
rect 58650 42080 58970 42110
rect 58650 42060 58660 42080
rect 57740 42050 57820 42060
rect 58160 42050 58240 42060
rect 58580 42050 58660 42060
rect 58960 42060 58970 42080
rect 59030 42060 59040 42120
rect 58960 42050 59040 42060
rect 58160 41990 58170 42050
rect 58230 42010 58240 42050
rect 58230 42000 58930 42010
rect 58230 41990 58870 42000
rect 58160 41980 58870 41990
rect 58870 41930 58930 41940
rect 58810 40820 58870 40830
rect 58160 40790 58810 40800
rect 57540 40730 57600 40740
rect 58160 40730 58170 40790
rect 58230 40770 58810 40790
rect 58230 40730 58240 40770
rect 58810 40750 58870 40760
rect 58960 40730 59020 40740
rect 57740 40720 57820 40730
rect 58160 40720 58240 40730
rect 58580 40720 58660 40730
rect 57740 40710 57750 40720
rect 57600 40680 57750 40710
rect 57540 40660 57600 40670
rect 57740 40660 57750 40680
rect 57810 40660 57820 40720
rect 57740 40650 57820 40660
rect 58580 40660 58590 40720
rect 58650 40710 58660 40720
rect 58650 40680 58960 40710
rect 58650 40660 58660 40680
rect 58960 40660 59020 40670
rect 58580 40650 58660 40660
rect 58150 40630 58250 40640
rect 58150 40560 58170 40630
rect 58240 40560 58250 40630
rect 58150 40520 58250 40560
rect 58150 40450 58170 40520
rect 58240 40450 58250 40520
rect 58150 40430 58250 40450
rect 57520 40410 57600 40420
rect 57520 40350 57530 40410
rect 57590 40400 57600 40410
rect 57740 40410 57820 40420
rect 57740 40400 57750 40410
rect 57590 40370 57750 40400
rect 57590 40350 57600 40370
rect 57520 40340 57600 40350
rect 57740 40350 57750 40370
rect 57810 40350 57820 40410
rect 58580 40410 58660 40420
rect 58580 40350 58590 40410
rect 58650 40400 58660 40410
rect 58960 40410 59040 40420
rect 58960 40400 58970 40410
rect 58650 40370 58970 40400
rect 58650 40350 58660 40370
rect 57740 40340 57820 40350
rect 58160 40340 58240 40350
rect 58580 40340 58660 40350
rect 58960 40350 58970 40370
rect 59030 40350 59040 40410
rect 58960 40340 59040 40350
rect 57160 39290 57220 39300
rect 57160 39220 57220 39230
rect 57250 39270 57480 39300
rect 57040 37150 57120 37160
rect 57040 37090 57050 37150
rect 57110 37090 57120 37150
rect 57040 37080 57120 37090
rect 56980 37010 57060 37020
rect 56980 36950 56990 37010
rect 57050 36950 57060 37010
rect 56980 36940 57060 36950
rect 56860 36870 56940 36880
rect 56860 36810 56870 36870
rect 56930 36810 56940 36870
rect 56860 36800 56940 36810
rect 56800 36730 56880 36740
rect 56800 36670 56810 36730
rect 56870 36670 56880 36730
rect 56800 36660 56880 36670
rect 54330 36400 54340 36460
rect 54400 36400 54410 36460
rect 57160 36460 57190 39220
rect 57250 36600 57280 39270
rect 57570 39240 57600 40340
rect 58160 40280 58170 40340
rect 58230 40300 58240 40340
rect 58230 40290 58930 40300
rect 58230 40280 58870 40290
rect 58160 40270 58870 40280
rect 58870 40220 58930 40230
rect 57340 39230 57400 39240
rect 57340 39160 57400 39170
rect 57430 39210 57600 39240
rect 57630 39680 57710 39690
rect 57630 39620 57640 39680
rect 57700 39620 57710 39680
rect 58700 39680 58780 39690
rect 58700 39620 58710 39680
rect 58770 39620 58780 39680
rect 57220 36590 57300 36600
rect 57220 36530 57230 36590
rect 57290 36530 57300 36590
rect 57220 36520 57300 36530
rect 57160 36450 57240 36460
rect 57160 36390 57170 36450
rect 57230 36390 57240 36450
rect 57160 36380 57240 36390
rect 52350 36170 52430 36180
rect 47360 36100 47440 36110
rect 52350 36110 52360 36170
rect 52420 36110 52430 36170
rect 54150 36120 54160 36180
rect 54220 36120 54230 36180
rect 57340 36180 57370 39160
rect 57430 36320 57460 39210
rect 57630 38840 57700 39620
rect 58700 39610 58780 39620
rect 58870 39680 58930 39690
rect 58870 39610 58930 39620
rect 57630 38830 57710 38840
rect 57630 38770 57640 38830
rect 57700 38770 57710 38830
rect 57630 38760 57710 38770
rect 58710 38700 58780 39610
rect 58900 38700 58930 39610
rect 58960 39240 58990 40340
rect 59080 39300 59110 43760
rect 59200 39360 59230 47180
rect 59320 39420 59350 48890
rect 63150 48830 63160 48890
rect 63220 48850 63230 48890
rect 63220 48840 63920 48850
rect 63220 48830 63860 48840
rect 63150 48820 63860 48830
rect 68140 48830 68150 48890
rect 68210 48850 68220 48890
rect 68210 48840 68910 48850
rect 68210 48830 68850 48840
rect 68140 48820 68850 48830
rect 63860 48770 63920 48780
rect 73130 48830 73140 48890
rect 73200 48850 73210 48890
rect 73200 48840 73900 48850
rect 73200 48830 73840 48840
rect 73130 48820 73840 48830
rect 68850 48770 68910 48780
rect 78120 48830 78130 48890
rect 78190 48850 78200 48890
rect 78190 48840 78890 48850
rect 78190 48830 78830 48840
rect 78120 48820 78830 48830
rect 73840 48770 73900 48780
rect 78830 48770 78890 48780
rect 63800 47660 63860 47670
rect 63150 47630 63800 47640
rect 62410 47570 62470 47580
rect 63150 47570 63160 47630
rect 63220 47610 63800 47630
rect 63220 47570 63230 47610
rect 68790 47660 68850 47670
rect 63800 47590 63860 47600
rect 68140 47630 68790 47640
rect 64070 47570 64130 47580
rect 62730 47560 62810 47570
rect 63150 47560 63230 47570
rect 63570 47560 63650 47570
rect 62730 47550 62740 47560
rect 62470 47520 62740 47550
rect 62410 47500 62470 47510
rect 62730 47500 62740 47520
rect 62800 47500 62810 47560
rect 62730 47490 62810 47500
rect 63570 47500 63580 47560
rect 63640 47550 63650 47560
rect 63640 47520 64070 47550
rect 63640 47500 63650 47520
rect 64070 47500 64130 47510
rect 67400 47570 67460 47580
rect 68140 47570 68150 47630
rect 68210 47610 68790 47630
rect 68210 47570 68220 47610
rect 73780 47660 73840 47670
rect 68790 47590 68850 47600
rect 73130 47630 73780 47640
rect 69060 47570 69120 47580
rect 67720 47560 67800 47570
rect 68140 47560 68220 47570
rect 68560 47560 68640 47570
rect 67720 47550 67730 47560
rect 67460 47520 67730 47550
rect 67400 47500 67460 47510
rect 67720 47500 67730 47520
rect 67790 47500 67800 47560
rect 63570 47490 63650 47500
rect 67720 47490 67800 47500
rect 68560 47500 68570 47560
rect 68630 47550 68640 47560
rect 68630 47520 69060 47550
rect 68630 47500 68640 47520
rect 69060 47500 69120 47510
rect 72510 47570 72570 47580
rect 73130 47570 73140 47630
rect 73200 47610 73780 47630
rect 73200 47570 73210 47610
rect 78770 47660 78830 47670
rect 73780 47590 73840 47600
rect 78120 47630 78770 47640
rect 73930 47570 73990 47580
rect 72710 47560 72790 47570
rect 73130 47560 73210 47570
rect 73550 47560 73630 47570
rect 72710 47550 72720 47560
rect 72570 47520 72720 47550
rect 72510 47500 72570 47510
rect 72710 47500 72720 47520
rect 72780 47500 72790 47560
rect 68560 47490 68640 47500
rect 72710 47490 72790 47500
rect 73550 47500 73560 47560
rect 73620 47550 73630 47560
rect 73620 47520 73930 47550
rect 73620 47500 73630 47520
rect 73930 47500 73990 47510
rect 77500 47570 77560 47580
rect 78120 47570 78130 47630
rect 78190 47610 78770 47630
rect 78190 47570 78200 47610
rect 78770 47590 78830 47600
rect 78920 47570 78980 47580
rect 77700 47560 77780 47570
rect 78120 47560 78200 47570
rect 78540 47560 78620 47570
rect 77700 47550 77710 47560
rect 77560 47520 77710 47550
rect 77500 47500 77560 47510
rect 77700 47500 77710 47520
rect 77770 47500 77780 47560
rect 73550 47490 73630 47500
rect 77700 47490 77780 47500
rect 78540 47500 78550 47560
rect 78610 47550 78620 47560
rect 78610 47520 78920 47550
rect 78610 47500 78620 47520
rect 78920 47500 78980 47510
rect 78540 47490 78620 47500
rect 63140 47470 63240 47480
rect 63140 47400 63160 47470
rect 63230 47400 63240 47470
rect 63140 47360 63240 47400
rect 63140 47290 63160 47360
rect 63230 47290 63240 47360
rect 63140 47270 63240 47290
rect 68130 47470 68230 47480
rect 68130 47400 68150 47470
rect 68220 47400 68230 47470
rect 68130 47360 68230 47400
rect 68130 47290 68150 47360
rect 68220 47290 68230 47360
rect 68130 47270 68230 47290
rect 73120 47470 73220 47480
rect 73120 47400 73140 47470
rect 73210 47400 73220 47470
rect 73120 47360 73220 47400
rect 73120 47290 73140 47360
rect 73210 47290 73220 47360
rect 73120 47270 73220 47290
rect 78110 47470 78210 47480
rect 78110 47400 78130 47470
rect 78200 47400 78210 47470
rect 78110 47360 78210 47400
rect 78110 47290 78130 47360
rect 78200 47290 78210 47360
rect 78110 47270 78210 47290
rect 62390 47250 62470 47260
rect 62390 47190 62400 47250
rect 62460 47240 62470 47250
rect 62730 47250 62810 47260
rect 62730 47240 62740 47250
rect 62460 47210 62740 47240
rect 62460 47190 62470 47210
rect 62390 47180 62470 47190
rect 62730 47190 62740 47210
rect 62800 47190 62810 47250
rect 63570 47250 63650 47260
rect 63570 47190 63580 47250
rect 63640 47240 63650 47250
rect 64070 47250 64150 47260
rect 64070 47240 64080 47250
rect 63640 47210 64080 47240
rect 63640 47190 63650 47210
rect 62730 47180 62810 47190
rect 63150 47180 63230 47190
rect 63570 47180 63650 47190
rect 64070 47190 64080 47210
rect 64140 47190 64150 47250
rect 64070 47180 64150 47190
rect 67380 47250 67460 47260
rect 67380 47190 67390 47250
rect 67450 47240 67460 47250
rect 67720 47250 67800 47260
rect 67720 47240 67730 47250
rect 67450 47210 67730 47240
rect 67450 47190 67460 47210
rect 67380 47180 67460 47190
rect 67720 47190 67730 47210
rect 67790 47190 67800 47250
rect 68560 47250 68640 47260
rect 68560 47190 68570 47250
rect 68630 47240 68640 47250
rect 69060 47250 69140 47260
rect 69060 47240 69070 47250
rect 68630 47210 69070 47240
rect 68630 47190 68640 47210
rect 67720 47180 67800 47190
rect 68140 47180 68220 47190
rect 68560 47180 68640 47190
rect 69060 47190 69070 47210
rect 69130 47190 69140 47250
rect 69060 47180 69140 47190
rect 72490 47250 72570 47260
rect 72490 47190 72500 47250
rect 72560 47240 72570 47250
rect 72710 47250 72790 47260
rect 72710 47240 72720 47250
rect 72560 47210 72720 47240
rect 72560 47190 72570 47210
rect 72490 47180 72570 47190
rect 72710 47190 72720 47210
rect 72780 47190 72790 47250
rect 73550 47250 73630 47260
rect 73550 47190 73560 47250
rect 73620 47240 73630 47250
rect 73930 47250 74010 47260
rect 73930 47240 73940 47250
rect 73620 47210 73940 47240
rect 73620 47190 73630 47210
rect 72710 47180 72790 47190
rect 73130 47180 73210 47190
rect 73550 47180 73630 47190
rect 73930 47190 73940 47210
rect 74000 47190 74010 47250
rect 73930 47180 74010 47190
rect 77480 47250 77560 47260
rect 77480 47190 77490 47250
rect 77550 47240 77560 47250
rect 77700 47250 77780 47260
rect 77700 47240 77710 47250
rect 77550 47210 77710 47240
rect 77550 47190 77560 47210
rect 77480 47180 77560 47190
rect 77700 47190 77710 47210
rect 77770 47190 77780 47250
rect 78540 47250 78620 47260
rect 78540 47190 78550 47250
rect 78610 47240 78620 47250
rect 78920 47250 79000 47260
rect 78920 47240 78930 47250
rect 78610 47210 78930 47240
rect 78610 47190 78620 47210
rect 77700 47180 77780 47190
rect 78120 47180 78200 47190
rect 78540 47180 78620 47190
rect 78920 47190 78930 47210
rect 78990 47190 79000 47250
rect 78920 47180 79000 47190
rect 59320 39390 59670 39420
rect 59200 39330 59490 39360
rect 59080 39270 59310 39300
rect 58960 39210 59130 39240
rect 58700 38690 58780 38700
rect 58700 38630 58710 38690
rect 58770 38630 58780 38690
rect 58850 38640 58860 38700
rect 58920 38640 58930 38700
rect 58700 38620 58780 38630
rect 59100 36320 59130 39210
rect 59160 39230 59220 39240
rect 59160 39160 59220 39170
rect 57400 36310 57480 36320
rect 57400 36250 57410 36310
rect 57470 36250 57480 36310
rect 59080 36260 59090 36320
rect 59150 36260 59160 36320
rect 57400 36240 57480 36250
rect 59190 36180 59220 39160
rect 59280 36600 59310 39270
rect 59340 39290 59400 39300
rect 59340 39220 59400 39230
rect 59260 36540 59270 36600
rect 59330 36540 59340 36600
rect 59370 36460 59400 39220
rect 59460 37160 59490 39330
rect 59520 39350 59580 39360
rect 59520 39280 59580 39290
rect 59440 37100 59450 37160
rect 59510 37100 59520 37160
rect 59550 37020 59580 39280
rect 59500 36960 59510 37020
rect 59570 36960 59580 37020
rect 59640 36880 59670 39390
rect 59700 39410 59760 39420
rect 59700 39340 59760 39350
rect 59620 36820 59630 36880
rect 59690 36820 59700 36880
rect 59730 36740 59760 39340
rect 62440 39300 62470 47180
rect 63150 47120 63160 47180
rect 63220 47140 63230 47180
rect 63220 47130 63920 47140
rect 63220 47120 63860 47130
rect 63150 47110 63860 47120
rect 63860 47060 63920 47070
rect 63800 45950 63860 45960
rect 63150 45920 63800 45930
rect 62530 45860 62590 45870
rect 63150 45860 63160 45920
rect 63220 45900 63800 45920
rect 63220 45860 63230 45900
rect 63800 45880 63860 45890
rect 63950 45860 64010 45870
rect 62730 45850 62810 45860
rect 63150 45850 63230 45860
rect 63570 45850 63650 45860
rect 62730 45840 62740 45850
rect 62590 45810 62740 45840
rect 62530 45790 62590 45800
rect 62730 45790 62740 45810
rect 62800 45790 62810 45850
rect 62730 45780 62810 45790
rect 63570 45790 63580 45850
rect 63640 45840 63650 45850
rect 63640 45810 63950 45840
rect 63640 45790 63650 45810
rect 63950 45790 64010 45800
rect 63570 45780 63650 45790
rect 63140 45760 63240 45770
rect 63140 45690 63160 45760
rect 63230 45690 63240 45760
rect 63140 45650 63240 45690
rect 63140 45580 63160 45650
rect 63230 45580 63240 45650
rect 63140 45560 63240 45580
rect 62510 45540 62590 45550
rect 62510 45480 62520 45540
rect 62580 45530 62590 45540
rect 62730 45540 62810 45550
rect 62730 45530 62740 45540
rect 62580 45500 62740 45530
rect 62580 45480 62590 45500
rect 62510 45470 62590 45480
rect 62730 45480 62740 45500
rect 62800 45480 62810 45540
rect 63570 45540 63650 45550
rect 63570 45480 63580 45540
rect 63640 45530 63650 45540
rect 63950 45540 64030 45550
rect 63950 45530 63960 45540
rect 63640 45500 63960 45530
rect 63640 45480 63650 45500
rect 62730 45470 62810 45480
rect 63150 45470 63230 45480
rect 63570 45470 63650 45480
rect 63950 45480 63960 45500
rect 64020 45480 64030 45540
rect 63950 45470 64030 45480
rect 63150 45410 63160 45470
rect 63220 45430 63230 45470
rect 63220 45420 63920 45430
rect 63220 45410 63860 45420
rect 63150 45400 63860 45410
rect 63860 45350 63920 45360
rect 63800 44240 63860 44250
rect 63150 44210 63800 44220
rect 62530 44150 62590 44160
rect 63150 44150 63160 44210
rect 63220 44190 63800 44210
rect 63220 44150 63230 44190
rect 63800 44170 63860 44180
rect 63950 44150 64010 44160
rect 62730 44140 62810 44150
rect 63150 44140 63230 44150
rect 63570 44140 63650 44150
rect 62730 44130 62740 44140
rect 62590 44100 62740 44130
rect 62530 44080 62590 44090
rect 62730 44080 62740 44100
rect 62800 44080 62810 44140
rect 62730 44070 62810 44080
rect 63570 44080 63580 44140
rect 63640 44130 63650 44140
rect 63640 44100 63950 44130
rect 63640 44080 63650 44100
rect 63950 44080 64010 44090
rect 63570 44070 63650 44080
rect 63140 44050 63240 44060
rect 63140 43980 63160 44050
rect 63230 43980 63240 44050
rect 63140 43940 63240 43980
rect 63140 43870 63160 43940
rect 63230 43870 63240 43940
rect 63140 43850 63240 43870
rect 62510 43830 62590 43840
rect 62510 43770 62520 43830
rect 62580 43820 62590 43830
rect 62730 43830 62810 43840
rect 62730 43820 62740 43830
rect 62580 43790 62740 43820
rect 62580 43770 62590 43790
rect 62510 43760 62590 43770
rect 62730 43770 62740 43790
rect 62800 43770 62810 43830
rect 63570 43830 63650 43840
rect 63570 43770 63580 43830
rect 63640 43820 63650 43830
rect 63950 43830 64030 43840
rect 63950 43820 63960 43830
rect 63640 43790 63960 43820
rect 63640 43770 63650 43790
rect 62730 43760 62810 43770
rect 63150 43760 63230 43770
rect 63570 43760 63650 43770
rect 63950 43770 63960 43790
rect 64020 43770 64030 43830
rect 63950 43760 64030 43770
rect 63150 43700 63160 43760
rect 63220 43720 63230 43760
rect 63220 43710 63920 43720
rect 63220 43700 63860 43710
rect 63150 43690 63860 43700
rect 63860 43640 63920 43650
rect 63800 42530 63860 42540
rect 63150 42500 63800 42510
rect 62530 42440 62590 42450
rect 63150 42440 63160 42500
rect 63220 42480 63800 42500
rect 63220 42440 63230 42480
rect 63800 42460 63860 42470
rect 63950 42440 64010 42450
rect 62730 42430 62810 42440
rect 63150 42430 63230 42440
rect 63570 42430 63650 42440
rect 62730 42420 62740 42430
rect 62590 42390 62740 42420
rect 62530 42370 62590 42380
rect 62730 42370 62740 42390
rect 62800 42370 62810 42430
rect 62730 42360 62810 42370
rect 63570 42370 63580 42430
rect 63640 42420 63650 42430
rect 63640 42390 63950 42420
rect 63640 42370 63650 42390
rect 63950 42370 64010 42380
rect 63570 42360 63650 42370
rect 63140 42340 63240 42350
rect 63140 42270 63160 42340
rect 63230 42270 63240 42340
rect 63140 42230 63240 42270
rect 63140 42160 63160 42230
rect 63230 42160 63240 42230
rect 63140 42140 63240 42160
rect 62510 42120 62590 42130
rect 62510 42060 62520 42120
rect 62580 42110 62590 42120
rect 62730 42120 62810 42130
rect 62730 42110 62740 42120
rect 62580 42080 62740 42110
rect 62580 42060 62590 42080
rect 62510 42050 62590 42060
rect 62730 42060 62740 42080
rect 62800 42060 62810 42120
rect 63570 42120 63650 42130
rect 63570 42060 63580 42120
rect 63640 42110 63650 42120
rect 63950 42120 64030 42130
rect 63950 42110 63960 42120
rect 63640 42080 63960 42110
rect 63640 42060 63650 42080
rect 62730 42050 62810 42060
rect 63150 42050 63230 42060
rect 63570 42050 63650 42060
rect 63950 42060 63960 42080
rect 64020 42060 64030 42120
rect 63950 42050 64030 42060
rect 63150 41990 63160 42050
rect 63220 42010 63230 42050
rect 63220 42000 63920 42010
rect 63220 41990 63860 42000
rect 63150 41980 63860 41990
rect 63860 41930 63920 41940
rect 63800 40820 63860 40830
rect 63150 40790 63800 40800
rect 62530 40730 62590 40740
rect 63150 40730 63160 40790
rect 63220 40770 63800 40790
rect 63220 40730 63230 40770
rect 63800 40750 63860 40760
rect 63950 40730 64010 40740
rect 62730 40720 62810 40730
rect 63150 40720 63230 40730
rect 63570 40720 63650 40730
rect 62730 40710 62740 40720
rect 62590 40680 62740 40710
rect 62530 40660 62590 40670
rect 62730 40660 62740 40680
rect 62800 40660 62810 40720
rect 62730 40650 62810 40660
rect 63570 40660 63580 40720
rect 63640 40710 63650 40720
rect 63640 40680 63950 40710
rect 63640 40660 63650 40680
rect 63950 40660 64010 40670
rect 63570 40650 63650 40660
rect 63140 40630 63240 40640
rect 63140 40560 63160 40630
rect 63230 40560 63240 40630
rect 63140 40520 63240 40560
rect 63140 40450 63160 40520
rect 63230 40450 63240 40520
rect 63140 40430 63240 40450
rect 62510 40410 62590 40420
rect 62510 40350 62520 40410
rect 62580 40400 62590 40410
rect 62730 40410 62810 40420
rect 62730 40400 62740 40410
rect 62580 40370 62740 40400
rect 62580 40350 62590 40370
rect 62510 40340 62590 40350
rect 62730 40350 62740 40370
rect 62800 40350 62810 40410
rect 63570 40410 63650 40420
rect 63570 40350 63580 40410
rect 63640 40400 63650 40410
rect 63950 40410 64030 40420
rect 63950 40400 63960 40410
rect 63640 40370 63960 40400
rect 63640 40350 63650 40370
rect 62730 40340 62810 40350
rect 63150 40340 63230 40350
rect 63570 40340 63650 40350
rect 63950 40350 63960 40370
rect 64020 40350 64030 40410
rect 63950 40340 64030 40350
rect 59680 36680 59690 36740
rect 59750 36680 59760 36740
rect 62150 39290 62210 39300
rect 62150 39220 62210 39230
rect 62240 39270 62470 39300
rect 59320 36400 59330 36460
rect 59390 36400 59400 36460
rect 62150 36460 62180 39220
rect 62240 36600 62270 39270
rect 62560 39240 62590 40340
rect 63150 40280 63160 40340
rect 63220 40300 63230 40340
rect 63220 40290 63920 40300
rect 63220 40280 63860 40290
rect 63150 40270 63860 40280
rect 63860 40220 63920 40230
rect 62330 39230 62390 39240
rect 62330 39160 62390 39170
rect 62420 39210 62590 39240
rect 62620 39680 62700 39690
rect 62620 39620 62630 39680
rect 62690 39620 62700 39680
rect 63690 39680 63770 39690
rect 63690 39620 63700 39680
rect 63760 39620 63770 39680
rect 62210 36590 62290 36600
rect 62210 36530 62220 36590
rect 62280 36530 62290 36590
rect 62210 36520 62290 36530
rect 62150 36450 62230 36460
rect 62150 36390 62160 36450
rect 62220 36390 62230 36450
rect 62150 36380 62230 36390
rect 57340 36170 57420 36180
rect 52350 36100 52430 36110
rect 57340 36110 57350 36170
rect 57410 36110 57420 36170
rect 59140 36120 59150 36180
rect 59210 36120 59220 36180
rect 62330 36180 62360 39160
rect 62420 36320 62450 39210
rect 62620 38840 62690 39620
rect 63690 39610 63770 39620
rect 63860 39680 63920 39690
rect 63860 39610 63920 39620
rect 62620 38830 62700 38840
rect 62620 38770 62630 38830
rect 62690 38770 62700 38830
rect 62620 38760 62700 38770
rect 63700 38700 63770 39610
rect 63890 38700 63920 39610
rect 63950 39240 63980 40340
rect 64070 39300 64100 47180
rect 67430 39300 67460 47180
rect 68140 47120 68150 47180
rect 68210 47140 68220 47180
rect 68210 47130 68910 47140
rect 68210 47120 68850 47130
rect 68140 47110 68850 47120
rect 68850 47060 68910 47070
rect 68790 45950 68850 45960
rect 68140 45920 68790 45930
rect 67520 45860 67580 45870
rect 68140 45860 68150 45920
rect 68210 45900 68790 45920
rect 68210 45860 68220 45900
rect 68790 45880 68850 45890
rect 68940 45860 69000 45870
rect 67720 45850 67800 45860
rect 68140 45850 68220 45860
rect 68560 45850 68640 45860
rect 67720 45840 67730 45850
rect 67580 45810 67730 45840
rect 67520 45790 67580 45800
rect 67720 45790 67730 45810
rect 67790 45790 67800 45850
rect 67720 45780 67800 45790
rect 68560 45790 68570 45850
rect 68630 45840 68640 45850
rect 68630 45810 68940 45840
rect 68630 45790 68640 45810
rect 68940 45790 69000 45800
rect 68560 45780 68640 45790
rect 68130 45760 68230 45770
rect 68130 45690 68150 45760
rect 68220 45690 68230 45760
rect 68130 45650 68230 45690
rect 68130 45580 68150 45650
rect 68220 45580 68230 45650
rect 68130 45560 68230 45580
rect 67500 45540 67580 45550
rect 67500 45480 67510 45540
rect 67570 45530 67580 45540
rect 67720 45540 67800 45550
rect 67720 45530 67730 45540
rect 67570 45500 67730 45530
rect 67570 45480 67580 45500
rect 67500 45470 67580 45480
rect 67720 45480 67730 45500
rect 67790 45480 67800 45540
rect 68560 45540 68640 45550
rect 68560 45480 68570 45540
rect 68630 45530 68640 45540
rect 68940 45540 69020 45550
rect 68940 45530 68950 45540
rect 68630 45500 68950 45530
rect 68630 45480 68640 45500
rect 67720 45470 67800 45480
rect 68140 45470 68220 45480
rect 68560 45470 68640 45480
rect 68940 45480 68950 45500
rect 69010 45480 69020 45540
rect 68940 45470 69020 45480
rect 68140 45410 68150 45470
rect 68210 45430 68220 45470
rect 68210 45420 68910 45430
rect 68210 45410 68850 45420
rect 68140 45400 68850 45410
rect 68850 45350 68910 45360
rect 68790 44240 68850 44250
rect 68140 44210 68790 44220
rect 67520 44150 67580 44160
rect 68140 44150 68150 44210
rect 68210 44190 68790 44210
rect 68210 44150 68220 44190
rect 68790 44170 68850 44180
rect 68940 44150 69000 44160
rect 67720 44140 67800 44150
rect 68140 44140 68220 44150
rect 68560 44140 68640 44150
rect 67720 44130 67730 44140
rect 67580 44100 67730 44130
rect 67520 44080 67580 44090
rect 67720 44080 67730 44100
rect 67790 44080 67800 44140
rect 67720 44070 67800 44080
rect 68560 44080 68570 44140
rect 68630 44130 68640 44140
rect 68630 44100 68940 44130
rect 68630 44080 68640 44100
rect 68940 44080 69000 44090
rect 68560 44070 68640 44080
rect 68130 44050 68230 44060
rect 68130 43980 68150 44050
rect 68220 43980 68230 44050
rect 68130 43940 68230 43980
rect 68130 43870 68150 43940
rect 68220 43870 68230 43940
rect 68130 43850 68230 43870
rect 67500 43830 67580 43840
rect 67500 43770 67510 43830
rect 67570 43820 67580 43830
rect 67720 43830 67800 43840
rect 67720 43820 67730 43830
rect 67570 43790 67730 43820
rect 67570 43770 67580 43790
rect 67500 43760 67580 43770
rect 67720 43770 67730 43790
rect 67790 43770 67800 43830
rect 68560 43830 68640 43840
rect 68560 43770 68570 43830
rect 68630 43820 68640 43830
rect 68940 43830 69020 43840
rect 68940 43820 68950 43830
rect 68630 43790 68950 43820
rect 68630 43770 68640 43790
rect 67720 43760 67800 43770
rect 68140 43760 68220 43770
rect 68560 43760 68640 43770
rect 68940 43770 68950 43790
rect 69010 43770 69020 43830
rect 68940 43760 69020 43770
rect 68140 43700 68150 43760
rect 68210 43720 68220 43760
rect 68210 43710 68910 43720
rect 68210 43700 68850 43710
rect 68140 43690 68850 43700
rect 68850 43640 68910 43650
rect 68790 42530 68850 42540
rect 68140 42500 68790 42510
rect 67520 42440 67580 42450
rect 68140 42440 68150 42500
rect 68210 42480 68790 42500
rect 68210 42440 68220 42480
rect 68790 42460 68850 42470
rect 68940 42440 69000 42450
rect 67720 42430 67800 42440
rect 68140 42430 68220 42440
rect 68560 42430 68640 42440
rect 67720 42420 67730 42430
rect 67580 42390 67730 42420
rect 67520 42370 67580 42380
rect 67720 42370 67730 42390
rect 67790 42370 67800 42430
rect 67720 42360 67800 42370
rect 68560 42370 68570 42430
rect 68630 42420 68640 42430
rect 68630 42390 68940 42420
rect 68630 42370 68640 42390
rect 68940 42370 69000 42380
rect 68560 42360 68640 42370
rect 68130 42340 68230 42350
rect 68130 42270 68150 42340
rect 68220 42270 68230 42340
rect 68130 42230 68230 42270
rect 68130 42160 68150 42230
rect 68220 42160 68230 42230
rect 68130 42140 68230 42160
rect 67500 42120 67580 42130
rect 67500 42060 67510 42120
rect 67570 42110 67580 42120
rect 67720 42120 67800 42130
rect 67720 42110 67730 42120
rect 67570 42080 67730 42110
rect 67570 42060 67580 42080
rect 67500 42050 67580 42060
rect 67720 42060 67730 42080
rect 67790 42060 67800 42120
rect 68560 42120 68640 42130
rect 68560 42060 68570 42120
rect 68630 42110 68640 42120
rect 68940 42120 69020 42130
rect 68940 42110 68950 42120
rect 68630 42080 68950 42110
rect 68630 42060 68640 42080
rect 67720 42050 67800 42060
rect 68140 42050 68220 42060
rect 68560 42050 68640 42060
rect 68940 42060 68950 42080
rect 69010 42060 69020 42120
rect 68940 42050 69020 42060
rect 68140 41990 68150 42050
rect 68210 42010 68220 42050
rect 68210 42000 68910 42010
rect 68210 41990 68850 42000
rect 68140 41980 68850 41990
rect 68850 41930 68910 41940
rect 68790 40820 68850 40830
rect 68140 40790 68790 40800
rect 67520 40730 67580 40740
rect 68140 40730 68150 40790
rect 68210 40770 68790 40790
rect 68210 40730 68220 40770
rect 68790 40750 68850 40760
rect 68940 40730 69000 40740
rect 67720 40720 67800 40730
rect 68140 40720 68220 40730
rect 68560 40720 68640 40730
rect 67720 40710 67730 40720
rect 67580 40680 67730 40710
rect 67520 40660 67580 40670
rect 67720 40660 67730 40680
rect 67790 40660 67800 40720
rect 67720 40650 67800 40660
rect 68560 40660 68570 40720
rect 68630 40710 68640 40720
rect 68630 40680 68940 40710
rect 68630 40660 68640 40680
rect 68940 40660 69000 40670
rect 68560 40650 68640 40660
rect 68130 40630 68230 40640
rect 68130 40560 68150 40630
rect 68220 40560 68230 40630
rect 68130 40520 68230 40560
rect 68130 40450 68150 40520
rect 68220 40450 68230 40520
rect 68130 40430 68230 40450
rect 67500 40410 67580 40420
rect 67500 40350 67510 40410
rect 67570 40400 67580 40410
rect 67720 40410 67800 40420
rect 67720 40400 67730 40410
rect 67570 40370 67730 40400
rect 67570 40350 67580 40370
rect 67500 40340 67580 40350
rect 67720 40350 67730 40370
rect 67790 40350 67800 40410
rect 68560 40410 68640 40420
rect 68560 40350 68570 40410
rect 68630 40400 68640 40410
rect 68940 40410 69020 40420
rect 68940 40400 68950 40410
rect 68630 40370 68950 40400
rect 68630 40350 68640 40370
rect 67720 40340 67800 40350
rect 68140 40340 68220 40350
rect 68560 40340 68640 40350
rect 68940 40350 68950 40370
rect 69010 40350 69020 40410
rect 68940 40340 69020 40350
rect 64070 39270 64300 39300
rect 63950 39210 64120 39240
rect 63690 38690 63770 38700
rect 63690 38630 63700 38690
rect 63760 38630 63770 38690
rect 63840 38640 63850 38700
rect 63910 38640 63920 38700
rect 63690 38620 63770 38630
rect 64090 36320 64120 39210
rect 64150 39230 64210 39240
rect 64150 39160 64210 39170
rect 62390 36310 62470 36320
rect 62390 36250 62400 36310
rect 62460 36250 62470 36310
rect 64070 36260 64080 36320
rect 64140 36260 64150 36320
rect 62390 36240 62470 36250
rect 64180 36180 64210 39160
rect 64270 36600 64300 39270
rect 64330 39290 64390 39300
rect 64330 39220 64390 39230
rect 64250 36540 64260 36600
rect 64320 36540 64330 36600
rect 64360 36460 64390 39220
rect 64310 36400 64320 36460
rect 64380 36400 64390 36460
rect 67140 39290 67200 39300
rect 67140 39220 67200 39230
rect 67230 39270 67460 39300
rect 67140 36460 67170 39220
rect 67230 36600 67260 39270
rect 67550 39240 67580 40340
rect 68140 40280 68150 40340
rect 68210 40300 68220 40340
rect 68210 40290 68910 40300
rect 68210 40280 68850 40290
rect 68140 40270 68850 40280
rect 68850 40220 68910 40230
rect 67320 39230 67380 39240
rect 67320 39160 67380 39170
rect 67410 39210 67580 39240
rect 67610 39680 67690 39690
rect 67610 39620 67620 39680
rect 67680 39620 67690 39680
rect 68680 39680 68760 39690
rect 68680 39620 68690 39680
rect 68750 39620 68760 39680
rect 67200 36590 67280 36600
rect 67200 36530 67210 36590
rect 67270 36530 67280 36590
rect 67200 36520 67280 36530
rect 67140 36450 67220 36460
rect 67140 36390 67150 36450
rect 67210 36390 67220 36450
rect 67140 36380 67220 36390
rect 62330 36170 62410 36180
rect 57340 36100 57420 36110
rect 62330 36110 62340 36170
rect 62400 36110 62410 36170
rect 64130 36120 64140 36180
rect 64200 36120 64210 36180
rect 67320 36180 67350 39160
rect 67410 36320 67440 39210
rect 67610 38840 67680 39620
rect 68680 39610 68760 39620
rect 68850 39680 68910 39690
rect 68850 39610 68910 39620
rect 67610 38830 67690 38840
rect 67610 38770 67620 38830
rect 67680 38770 67690 38830
rect 67610 38760 67690 38770
rect 68690 38700 68760 39610
rect 68880 38700 68910 39610
rect 68940 39240 68970 40340
rect 69060 39300 69090 47180
rect 73130 47120 73140 47180
rect 73200 47140 73210 47180
rect 73200 47130 73900 47140
rect 73200 47120 73840 47130
rect 73130 47110 73840 47120
rect 78120 47120 78130 47180
rect 78190 47140 78200 47180
rect 78190 47130 78890 47140
rect 78190 47120 78830 47130
rect 78120 47110 78830 47120
rect 73840 47060 73900 47070
rect 78830 47060 78890 47070
rect 73780 45950 73840 45960
rect 73130 45920 73780 45930
rect 72510 45860 72570 45870
rect 73130 45860 73140 45920
rect 73200 45900 73780 45920
rect 73200 45860 73210 45900
rect 78770 45950 78830 45960
rect 73780 45880 73840 45890
rect 78120 45920 78770 45930
rect 73930 45860 73990 45870
rect 72710 45850 72790 45860
rect 73130 45850 73210 45860
rect 73550 45850 73630 45860
rect 72710 45840 72720 45850
rect 72570 45810 72720 45840
rect 72510 45790 72570 45800
rect 72710 45790 72720 45810
rect 72780 45790 72790 45850
rect 72710 45780 72790 45790
rect 73550 45790 73560 45850
rect 73620 45840 73630 45850
rect 73620 45810 73930 45840
rect 73620 45790 73630 45810
rect 73930 45790 73990 45800
rect 77500 45860 77560 45870
rect 78120 45860 78130 45920
rect 78190 45900 78770 45920
rect 78190 45860 78200 45900
rect 78770 45880 78830 45890
rect 78920 45860 78980 45870
rect 77700 45850 77780 45860
rect 78120 45850 78200 45860
rect 78540 45850 78620 45860
rect 77700 45840 77710 45850
rect 77560 45810 77710 45840
rect 77500 45790 77560 45800
rect 77700 45790 77710 45810
rect 77770 45790 77780 45850
rect 73550 45780 73630 45790
rect 77700 45780 77780 45790
rect 78540 45790 78550 45850
rect 78610 45840 78620 45850
rect 78610 45810 78920 45840
rect 78610 45790 78620 45810
rect 78920 45790 78980 45800
rect 78540 45780 78620 45790
rect 73120 45760 73220 45770
rect 73120 45690 73140 45760
rect 73210 45690 73220 45760
rect 73120 45650 73220 45690
rect 73120 45580 73140 45650
rect 73210 45580 73220 45650
rect 73120 45560 73220 45580
rect 78110 45760 78210 45770
rect 78110 45690 78130 45760
rect 78200 45690 78210 45760
rect 78110 45650 78210 45690
rect 78110 45580 78130 45650
rect 78200 45580 78210 45650
rect 78110 45560 78210 45580
rect 72490 45540 72570 45550
rect 72490 45480 72500 45540
rect 72560 45530 72570 45540
rect 72710 45540 72790 45550
rect 72710 45530 72720 45540
rect 72560 45500 72720 45530
rect 72560 45480 72570 45500
rect 72490 45470 72570 45480
rect 72710 45480 72720 45500
rect 72780 45480 72790 45540
rect 73550 45540 73630 45550
rect 73550 45480 73560 45540
rect 73620 45530 73630 45540
rect 73930 45540 74010 45550
rect 73930 45530 73940 45540
rect 73620 45500 73940 45530
rect 73620 45480 73630 45500
rect 72710 45470 72790 45480
rect 73130 45470 73210 45480
rect 73550 45470 73630 45480
rect 73930 45480 73940 45500
rect 74000 45480 74010 45540
rect 73930 45470 74010 45480
rect 77480 45540 77560 45550
rect 77480 45480 77490 45540
rect 77550 45530 77560 45540
rect 77700 45540 77780 45550
rect 77700 45530 77710 45540
rect 77550 45500 77710 45530
rect 77550 45480 77560 45500
rect 77480 45470 77560 45480
rect 77700 45480 77710 45500
rect 77770 45480 77780 45540
rect 78540 45540 78620 45550
rect 78540 45480 78550 45540
rect 78610 45530 78620 45540
rect 78920 45540 79000 45550
rect 78920 45530 78930 45540
rect 78610 45500 78930 45530
rect 78610 45480 78620 45500
rect 77700 45470 77780 45480
rect 78120 45470 78200 45480
rect 78540 45470 78620 45480
rect 78920 45480 78930 45500
rect 78990 45480 79000 45540
rect 78920 45470 79000 45480
rect 73130 45410 73140 45470
rect 73200 45430 73210 45470
rect 73200 45420 73900 45430
rect 73200 45410 73840 45420
rect 73130 45400 73840 45410
rect 78120 45410 78130 45470
rect 78190 45430 78200 45470
rect 78190 45420 78890 45430
rect 78190 45410 78830 45420
rect 78120 45400 78830 45410
rect 73840 45350 73900 45360
rect 78830 45350 78890 45360
rect 73780 44240 73840 44250
rect 73130 44210 73780 44220
rect 72510 44150 72570 44160
rect 73130 44150 73140 44210
rect 73200 44190 73780 44210
rect 73200 44150 73210 44190
rect 78770 44240 78830 44250
rect 73780 44170 73840 44180
rect 78120 44210 78770 44220
rect 73930 44150 73990 44160
rect 72710 44140 72790 44150
rect 73130 44140 73210 44150
rect 73550 44140 73630 44150
rect 72710 44130 72720 44140
rect 72570 44100 72720 44130
rect 72510 44080 72570 44090
rect 72710 44080 72720 44100
rect 72780 44080 72790 44140
rect 72710 44070 72790 44080
rect 73550 44080 73560 44140
rect 73620 44130 73630 44140
rect 73620 44100 73930 44130
rect 73620 44080 73630 44100
rect 73930 44080 73990 44090
rect 77500 44150 77560 44160
rect 78120 44150 78130 44210
rect 78190 44190 78770 44210
rect 78190 44150 78200 44190
rect 78770 44170 78830 44180
rect 78920 44150 78980 44160
rect 77700 44140 77780 44150
rect 78120 44140 78200 44150
rect 78540 44140 78620 44150
rect 77700 44130 77710 44140
rect 77560 44100 77710 44130
rect 77500 44080 77560 44090
rect 77700 44080 77710 44100
rect 77770 44080 77780 44140
rect 73550 44070 73630 44080
rect 77700 44070 77780 44080
rect 78540 44080 78550 44140
rect 78610 44130 78620 44140
rect 78610 44100 78920 44130
rect 78610 44080 78620 44100
rect 78920 44080 78980 44090
rect 78540 44070 78620 44080
rect 73120 44050 73220 44060
rect 73120 43980 73140 44050
rect 73210 43980 73220 44050
rect 73120 43940 73220 43980
rect 73120 43870 73140 43940
rect 73210 43870 73220 43940
rect 73120 43850 73220 43870
rect 78110 44050 78210 44060
rect 78110 43980 78130 44050
rect 78200 43980 78210 44050
rect 78110 43940 78210 43980
rect 78110 43870 78130 43940
rect 78200 43870 78210 43940
rect 78110 43850 78210 43870
rect 72490 43830 72570 43840
rect 72490 43770 72500 43830
rect 72560 43820 72570 43830
rect 72710 43830 72790 43840
rect 72710 43820 72720 43830
rect 72560 43790 72720 43820
rect 72560 43770 72570 43790
rect 72490 43760 72570 43770
rect 72710 43770 72720 43790
rect 72780 43770 72790 43830
rect 73550 43830 73630 43840
rect 73550 43770 73560 43830
rect 73620 43820 73630 43830
rect 73930 43830 74010 43840
rect 73930 43820 73940 43830
rect 73620 43790 73940 43820
rect 73620 43770 73630 43790
rect 72710 43760 72790 43770
rect 73130 43760 73210 43770
rect 73550 43760 73630 43770
rect 73930 43770 73940 43790
rect 74000 43770 74010 43830
rect 73930 43760 74010 43770
rect 77480 43830 77560 43840
rect 77480 43770 77490 43830
rect 77550 43820 77560 43830
rect 77700 43830 77780 43840
rect 77700 43820 77710 43830
rect 77550 43790 77710 43820
rect 77550 43770 77560 43790
rect 77480 43760 77560 43770
rect 77700 43770 77710 43790
rect 77770 43770 77780 43830
rect 78540 43830 78620 43840
rect 78540 43770 78550 43830
rect 78610 43820 78620 43830
rect 78920 43830 79000 43840
rect 78920 43820 78930 43830
rect 78610 43790 78930 43820
rect 78610 43770 78620 43790
rect 77700 43760 77780 43770
rect 78120 43760 78200 43770
rect 78540 43760 78620 43770
rect 78920 43770 78930 43790
rect 78990 43770 79000 43830
rect 78920 43760 79000 43770
rect 73130 43700 73140 43760
rect 73200 43720 73210 43760
rect 73200 43710 73900 43720
rect 73200 43700 73840 43710
rect 73130 43690 73840 43700
rect 78120 43700 78130 43760
rect 78190 43720 78200 43760
rect 78190 43710 78890 43720
rect 78190 43700 78830 43710
rect 78120 43690 78830 43700
rect 73840 43640 73900 43650
rect 78830 43640 78890 43650
rect 73780 42530 73840 42540
rect 73130 42500 73780 42510
rect 72510 42440 72570 42450
rect 73130 42440 73140 42500
rect 73200 42480 73780 42500
rect 73200 42440 73210 42480
rect 78770 42530 78830 42540
rect 73780 42460 73840 42470
rect 78120 42500 78770 42510
rect 73930 42440 73990 42450
rect 72710 42430 72790 42440
rect 73130 42430 73210 42440
rect 73550 42430 73630 42440
rect 72710 42420 72720 42430
rect 72570 42390 72720 42420
rect 72510 42370 72570 42380
rect 72710 42370 72720 42390
rect 72780 42370 72790 42430
rect 72710 42360 72790 42370
rect 73550 42370 73560 42430
rect 73620 42420 73630 42430
rect 73620 42390 73930 42420
rect 73620 42370 73630 42390
rect 73930 42370 73990 42380
rect 77500 42440 77560 42450
rect 78120 42440 78130 42500
rect 78190 42480 78770 42500
rect 78190 42440 78200 42480
rect 78770 42460 78830 42470
rect 78920 42440 78980 42450
rect 77700 42430 77780 42440
rect 78120 42430 78200 42440
rect 78540 42430 78620 42440
rect 77700 42420 77710 42430
rect 77560 42390 77710 42420
rect 77500 42370 77560 42380
rect 77700 42370 77710 42390
rect 77770 42370 77780 42430
rect 73550 42360 73630 42370
rect 77700 42360 77780 42370
rect 78540 42370 78550 42430
rect 78610 42420 78620 42430
rect 78610 42390 78920 42420
rect 78610 42370 78620 42390
rect 78920 42370 78980 42380
rect 78540 42360 78620 42370
rect 73120 42340 73220 42350
rect 73120 42270 73140 42340
rect 73210 42270 73220 42340
rect 73120 42230 73220 42270
rect 73120 42160 73140 42230
rect 73210 42160 73220 42230
rect 73120 42140 73220 42160
rect 78110 42340 78210 42350
rect 78110 42270 78130 42340
rect 78200 42270 78210 42340
rect 78110 42230 78210 42270
rect 78110 42160 78130 42230
rect 78200 42160 78210 42230
rect 78110 42140 78210 42160
rect 72490 42120 72570 42130
rect 72490 42060 72500 42120
rect 72560 42110 72570 42120
rect 72710 42120 72790 42130
rect 72710 42110 72720 42120
rect 72560 42080 72720 42110
rect 72560 42060 72570 42080
rect 72490 42050 72570 42060
rect 72710 42060 72720 42080
rect 72780 42060 72790 42120
rect 73550 42120 73630 42130
rect 73550 42060 73560 42120
rect 73620 42110 73630 42120
rect 73930 42120 74010 42130
rect 73930 42110 73940 42120
rect 73620 42080 73940 42110
rect 73620 42060 73630 42080
rect 72710 42050 72790 42060
rect 73130 42050 73210 42060
rect 73550 42050 73630 42060
rect 73930 42060 73940 42080
rect 74000 42060 74010 42120
rect 73930 42050 74010 42060
rect 77480 42120 77560 42130
rect 77480 42060 77490 42120
rect 77550 42110 77560 42120
rect 77700 42120 77780 42130
rect 77700 42110 77710 42120
rect 77550 42080 77710 42110
rect 77550 42060 77560 42080
rect 77480 42050 77560 42060
rect 77700 42060 77710 42080
rect 77770 42060 77780 42120
rect 78540 42120 78620 42130
rect 78540 42060 78550 42120
rect 78610 42110 78620 42120
rect 78920 42120 79000 42130
rect 78920 42110 78930 42120
rect 78610 42080 78930 42110
rect 78610 42060 78620 42080
rect 77700 42050 77780 42060
rect 78120 42050 78200 42060
rect 78540 42050 78620 42060
rect 78920 42060 78930 42080
rect 78990 42060 79000 42120
rect 78920 42050 79000 42060
rect 73130 41990 73140 42050
rect 73200 42010 73210 42050
rect 73200 42000 73900 42010
rect 73200 41990 73840 42000
rect 73130 41980 73840 41990
rect 78120 41990 78130 42050
rect 78190 42010 78200 42050
rect 78190 42000 78890 42010
rect 78190 41990 78830 42000
rect 78120 41980 78830 41990
rect 73840 41930 73900 41940
rect 78830 41930 78890 41940
rect 73780 40820 73840 40830
rect 73130 40790 73780 40800
rect 72510 40730 72570 40740
rect 73130 40730 73140 40790
rect 73200 40770 73780 40790
rect 73200 40730 73210 40770
rect 78770 40820 78830 40830
rect 73780 40750 73840 40760
rect 78120 40790 78770 40800
rect 73930 40730 73990 40740
rect 72710 40720 72790 40730
rect 73130 40720 73210 40730
rect 73550 40720 73630 40730
rect 72710 40710 72720 40720
rect 72570 40680 72720 40710
rect 72510 40660 72570 40670
rect 72710 40660 72720 40680
rect 72780 40660 72790 40720
rect 72710 40650 72790 40660
rect 73550 40660 73560 40720
rect 73620 40710 73630 40720
rect 73620 40680 73930 40710
rect 73620 40660 73630 40680
rect 73930 40660 73990 40670
rect 77500 40730 77560 40740
rect 78120 40730 78130 40790
rect 78190 40770 78770 40790
rect 78190 40730 78200 40770
rect 78770 40750 78830 40760
rect 78920 40730 78980 40740
rect 77700 40720 77780 40730
rect 78120 40720 78200 40730
rect 78540 40720 78620 40730
rect 77700 40710 77710 40720
rect 77560 40680 77710 40710
rect 77500 40660 77560 40670
rect 77700 40660 77710 40680
rect 77770 40660 77780 40720
rect 73550 40650 73630 40660
rect 77700 40650 77780 40660
rect 78540 40660 78550 40720
rect 78610 40710 78620 40720
rect 78610 40680 78920 40710
rect 78610 40660 78620 40680
rect 78920 40660 78980 40670
rect 78540 40650 78620 40660
rect 73120 40630 73220 40640
rect 73120 40560 73140 40630
rect 73210 40560 73220 40630
rect 73120 40520 73220 40560
rect 73120 40450 73140 40520
rect 73210 40450 73220 40520
rect 73120 40430 73220 40450
rect 78110 40630 78210 40640
rect 78110 40560 78130 40630
rect 78200 40560 78210 40630
rect 78110 40520 78210 40560
rect 78110 40450 78130 40520
rect 78200 40450 78210 40520
rect 78110 40430 78210 40450
rect 72490 40410 72570 40420
rect 72490 40350 72500 40410
rect 72560 40400 72570 40410
rect 72710 40410 72790 40420
rect 72710 40400 72720 40410
rect 72560 40370 72720 40400
rect 72560 40350 72570 40370
rect 72490 40340 72570 40350
rect 72710 40350 72720 40370
rect 72780 40350 72790 40410
rect 73550 40410 73630 40420
rect 73550 40350 73560 40410
rect 73620 40400 73630 40410
rect 73930 40410 74010 40420
rect 73930 40400 73940 40410
rect 73620 40370 73940 40400
rect 73620 40350 73630 40370
rect 72710 40340 72790 40350
rect 73130 40340 73210 40350
rect 73550 40340 73630 40350
rect 73930 40350 73940 40370
rect 74000 40350 74010 40410
rect 73930 40340 74010 40350
rect 77480 40410 77560 40420
rect 77480 40350 77490 40410
rect 77550 40400 77560 40410
rect 77700 40410 77780 40420
rect 77700 40400 77710 40410
rect 77550 40370 77710 40400
rect 77550 40350 77560 40370
rect 77480 40340 77560 40350
rect 77700 40350 77710 40370
rect 77770 40350 77780 40410
rect 78540 40410 78620 40420
rect 78540 40350 78550 40410
rect 78610 40400 78620 40410
rect 78920 40410 79000 40420
rect 78920 40400 78930 40410
rect 78610 40370 78930 40400
rect 78610 40350 78620 40370
rect 77700 40340 77780 40350
rect 78120 40340 78200 40350
rect 78540 40340 78620 40350
rect 78920 40350 78930 40370
rect 78990 40350 79000 40410
rect 78920 40340 79000 40350
rect 69060 39270 69290 39300
rect 68940 39210 69110 39240
rect 68680 38690 68760 38700
rect 68680 38630 68690 38690
rect 68750 38630 68760 38690
rect 68830 38640 68840 38700
rect 68900 38640 68910 38700
rect 68680 38620 68760 38630
rect 69080 36320 69110 39210
rect 69140 39230 69200 39240
rect 69140 39160 69200 39170
rect 67380 36310 67460 36320
rect 67380 36250 67390 36310
rect 67450 36250 67460 36310
rect 69060 36260 69070 36320
rect 69130 36260 69140 36320
rect 67380 36240 67460 36250
rect 69170 36180 69200 39160
rect 69260 36600 69290 39270
rect 69320 39290 69380 39300
rect 72540 39240 72570 40340
rect 73130 40280 73140 40340
rect 73200 40300 73210 40340
rect 73200 40290 73900 40300
rect 73200 40280 73840 40290
rect 73130 40270 73840 40280
rect 73840 40220 73900 40230
rect 69320 39220 69380 39230
rect 69240 36540 69250 36600
rect 69310 36540 69320 36600
rect 69350 36460 69380 39220
rect 69300 36400 69310 36460
rect 69370 36400 69380 36460
rect 72310 39230 72370 39240
rect 72310 39160 72370 39170
rect 72400 39210 72570 39240
rect 72600 39680 72680 39690
rect 72600 39620 72610 39680
rect 72670 39620 72680 39680
rect 73670 39680 73750 39690
rect 73670 39620 73680 39680
rect 73740 39620 73750 39680
rect 67320 36170 67400 36180
rect 62330 36100 62410 36110
rect 67320 36110 67330 36170
rect 67390 36110 67400 36170
rect 69120 36120 69130 36180
rect 69190 36120 69200 36180
rect 72310 36180 72340 39160
rect 72400 36320 72430 39210
rect 72600 38840 72670 39620
rect 73670 39610 73750 39620
rect 73840 39680 73900 39690
rect 73840 39610 73900 39620
rect 72600 38830 72680 38840
rect 72600 38770 72610 38830
rect 72670 38770 72680 38830
rect 72600 38760 72680 38770
rect 73680 38700 73750 39610
rect 73870 38700 73900 39610
rect 73930 39240 73960 40340
rect 77530 39240 77560 40340
rect 78120 40280 78130 40340
rect 78190 40300 78200 40340
rect 78190 40290 78890 40300
rect 78190 40280 78830 40290
rect 78120 40270 78830 40280
rect 78830 40220 78890 40230
rect 73930 39210 74100 39240
rect 73670 38690 73750 38700
rect 73670 38630 73680 38690
rect 73740 38630 73750 38690
rect 73820 38640 73830 38700
rect 73890 38640 73900 38700
rect 73670 38620 73750 38630
rect 74070 36320 74100 39210
rect 74130 39230 74190 39240
rect 74130 39160 74190 39170
rect 72370 36310 72450 36320
rect 72370 36250 72380 36310
rect 72440 36250 72450 36310
rect 74050 36260 74060 36320
rect 74120 36260 74130 36320
rect 72370 36240 72450 36250
rect 74160 36180 74190 39160
rect 72310 36170 72390 36180
rect 67320 36100 67400 36110
rect 72310 36110 72320 36170
rect 72380 36110 72390 36170
rect 74110 36120 74120 36180
rect 74180 36120 74190 36180
rect 77300 39230 77360 39240
rect 77300 39160 77360 39170
rect 77390 39210 77560 39240
rect 77590 39680 77670 39690
rect 77590 39620 77600 39680
rect 77660 39620 77670 39680
rect 78660 39680 78740 39690
rect 78660 39620 78670 39680
rect 78730 39620 78740 39680
rect 77300 36180 77330 39160
rect 77390 36320 77420 39210
rect 77590 38840 77660 39620
rect 78660 39610 78740 39620
rect 78830 39680 78890 39690
rect 78830 39610 78890 39620
rect 77590 38830 77670 38840
rect 77590 38770 77600 38830
rect 77660 38770 77670 38830
rect 77590 38760 77670 38770
rect 78670 38700 78740 39610
rect 78860 38700 78890 39610
rect 78920 39240 78950 40340
rect 78920 39210 79090 39240
rect 78660 38690 78740 38700
rect 78660 38630 78670 38690
rect 78730 38630 78740 38690
rect 78810 38640 78820 38700
rect 78880 38640 78890 38700
rect 78660 38620 78740 38630
rect 79060 36320 79090 39210
rect 79120 39230 79180 39240
rect 79120 39160 79180 39170
rect 77360 36310 77440 36320
rect 77360 36250 77370 36310
rect 77430 36250 77440 36310
rect 79040 36260 79050 36320
rect 79110 36260 79120 36320
rect 77360 36240 77440 36250
rect 79150 36180 79180 39160
rect 77300 36170 77380 36180
rect 72310 36100 72390 36110
rect 77300 36110 77310 36170
rect 77370 36110 77380 36170
rect 79100 36120 79110 36180
rect 79170 36120 79180 36180
rect 77300 36100 77380 36110
rect 2350 30940 2430 30950
rect 2350 30880 2360 30940
rect 2420 30880 2430 30940
rect 7340 30940 7420 30950
rect 2350 30870 2430 30880
rect 4150 30870 4160 30930
rect 4220 30870 4230 30930
rect 2350 27890 2380 30870
rect 2410 30800 2490 30810
rect 2410 30740 2420 30800
rect 2480 30740 2490 30800
rect 2410 30730 2490 30740
rect 4090 30730 4100 30790
rect 4160 30730 4170 30790
rect 2350 27880 2410 27890
rect 2350 27810 2410 27820
rect 2440 27840 2470 30730
rect 3710 28420 3790 28430
rect 3710 28360 3720 28420
rect 3780 28360 3790 28420
rect 3710 28350 3790 28360
rect 3860 28350 3870 28410
rect 3930 28350 3940 28410
rect 2640 28280 2720 28290
rect 2640 28220 2650 28280
rect 2710 28220 2720 28280
rect 2640 28210 2720 28220
rect 2440 27810 2610 27840
rect 2580 27360 2610 27810
rect 2640 27430 2710 28210
rect 3720 27440 3790 28350
rect 3910 27440 3940 28350
rect 4110 27840 4140 30730
rect 4200 27890 4230 30870
rect 3710 27430 3790 27440
rect 2640 27370 2650 27430
rect 2710 27370 2720 27430
rect 2640 27360 2720 27370
rect 3710 27370 3720 27430
rect 3780 27370 3790 27430
rect 3710 27360 3790 27370
rect 3880 27430 3940 27440
rect 3880 27360 3940 27370
rect 3970 27810 4140 27840
rect 4170 27880 4230 27890
rect 4170 27810 4230 27820
rect 7340 30880 7350 30940
rect 7410 30880 7420 30940
rect 12330 30940 12410 30950
rect 7340 30870 7420 30880
rect 9140 30870 9150 30930
rect 9210 30870 9220 30930
rect 7340 27890 7370 30870
rect 7400 30800 7480 30810
rect 7400 30740 7410 30800
rect 7470 30740 7480 30800
rect 7400 30730 7480 30740
rect 9080 30730 9090 30790
rect 9150 30730 9160 30790
rect 7340 27880 7400 27890
rect 7340 27810 7400 27820
rect 7430 27840 7460 30730
rect 8700 28420 8780 28430
rect 8700 28360 8710 28420
rect 8770 28360 8780 28420
rect 8700 28350 8780 28360
rect 8850 28350 8860 28410
rect 8920 28350 8930 28410
rect 7630 28280 7710 28290
rect 7630 28220 7640 28280
rect 7700 28220 7710 28280
rect 7630 28210 7710 28220
rect 7430 27810 7600 27840
rect 3970 27360 4000 27810
rect 7570 27360 7600 27810
rect 7630 27430 7700 28210
rect 8710 27440 8780 28350
rect 8900 27440 8930 28350
rect 9100 27840 9130 30730
rect 9190 27890 9220 30870
rect 12330 30880 12340 30940
rect 12400 30880 12410 30940
rect 17320 30940 17400 30950
rect 12330 30870 12410 30880
rect 14130 30870 14140 30930
rect 14200 30870 14210 30930
rect 8700 27430 8780 27440
rect 7630 27370 7640 27430
rect 7700 27370 7710 27430
rect 7630 27360 7710 27370
rect 8700 27370 8710 27430
rect 8770 27370 8780 27430
rect 8700 27360 8780 27370
rect 8870 27430 8930 27440
rect 8870 27360 8930 27370
rect 8960 27810 9130 27840
rect 9160 27880 9220 27890
rect 9160 27810 9220 27820
rect 12150 30660 12230 30670
rect 12150 30600 12160 30660
rect 12220 30600 12230 30660
rect 12150 30590 12230 30600
rect 12150 27830 12180 30590
rect 12210 30520 12290 30530
rect 12210 30460 12220 30520
rect 12280 30460 12290 30520
rect 12210 30450 12290 30460
rect 12150 27820 12210 27830
rect 8960 27360 8990 27810
rect 12150 27750 12210 27760
rect 12240 27780 12270 30450
rect 12330 27890 12360 30870
rect 12390 30800 12470 30810
rect 12390 30740 12400 30800
rect 12460 30740 12470 30800
rect 12390 30730 12470 30740
rect 14070 30730 14080 30790
rect 14140 30730 14150 30790
rect 12330 27880 12390 27890
rect 12330 27810 12390 27820
rect 12420 27840 12450 30730
rect 13690 28420 13770 28430
rect 13690 28360 13700 28420
rect 13760 28360 13770 28420
rect 13690 28350 13770 28360
rect 13840 28350 13850 28410
rect 13910 28350 13920 28410
rect 12620 28280 12700 28290
rect 12620 28220 12630 28280
rect 12690 28220 12700 28280
rect 12620 28210 12700 28220
rect 12420 27810 12590 27840
rect 12240 27750 12470 27780
rect 12440 27360 12470 27750
rect 12560 27360 12590 27810
rect 12620 27430 12690 28210
rect 13700 27440 13770 28350
rect 13890 27440 13920 28350
rect 14090 27840 14120 30730
rect 14180 27890 14210 30870
rect 17320 30880 17330 30940
rect 17390 30880 17400 30940
rect 22310 30940 22390 30950
rect 17320 30870 17400 30880
rect 19120 30870 19130 30930
rect 19190 30870 19200 30930
rect 17140 30660 17220 30670
rect 14310 30590 14320 30650
rect 14380 30590 14390 30650
rect 14250 30450 14260 30510
rect 14320 30450 14330 30510
rect 13690 27430 13770 27440
rect 12620 27370 12630 27430
rect 12690 27370 12700 27430
rect 12620 27360 12700 27370
rect 13690 27370 13700 27430
rect 13760 27370 13770 27430
rect 13690 27360 13770 27370
rect 13860 27430 13920 27440
rect 13860 27360 13920 27370
rect 13950 27810 14120 27840
rect 14150 27880 14210 27890
rect 14150 27810 14210 27820
rect 13950 27360 13980 27810
rect 14270 27780 14300 30450
rect 14360 27830 14390 30590
rect 14070 27750 14300 27780
rect 14330 27820 14390 27830
rect 14330 27750 14390 27760
rect 17140 30600 17150 30660
rect 17210 30600 17220 30660
rect 17140 30590 17220 30600
rect 17140 27830 17170 30590
rect 17200 30520 17280 30530
rect 17200 30460 17210 30520
rect 17270 30460 17280 30520
rect 17200 30450 17280 30460
rect 17140 27820 17200 27830
rect 17140 27750 17200 27760
rect 17230 27780 17260 30450
rect 17320 27890 17350 30870
rect 17380 30800 17460 30810
rect 17380 30740 17390 30800
rect 17450 30740 17460 30800
rect 17380 30730 17460 30740
rect 19060 30730 19070 30790
rect 19130 30730 19140 30790
rect 17320 27880 17380 27890
rect 17320 27810 17380 27820
rect 17410 27840 17440 30730
rect 18680 28420 18760 28430
rect 18680 28360 18690 28420
rect 18750 28360 18760 28420
rect 18680 28350 18760 28360
rect 18830 28350 18840 28410
rect 18900 28350 18910 28410
rect 17610 28280 17690 28290
rect 17610 28220 17620 28280
rect 17680 28220 17690 28280
rect 17610 28210 17690 28220
rect 17410 27810 17580 27840
rect 17230 27750 17460 27780
rect 14070 27360 14100 27750
rect 17430 27360 17460 27750
rect 17550 27360 17580 27810
rect 17610 27430 17680 28210
rect 18690 27440 18760 28350
rect 18880 27440 18910 28350
rect 19080 27840 19110 30730
rect 19170 27890 19200 30870
rect 22310 30880 22320 30940
rect 22380 30880 22390 30940
rect 27300 30940 27380 30950
rect 22310 30870 22390 30880
rect 24110 30870 24120 30930
rect 24180 30870 24190 30930
rect 22130 30660 22210 30670
rect 19300 30590 19310 30650
rect 19370 30590 19380 30650
rect 19240 30450 19250 30510
rect 19310 30450 19320 30510
rect 18680 27430 18760 27440
rect 17610 27370 17620 27430
rect 17680 27370 17690 27430
rect 17610 27360 17690 27370
rect 18680 27370 18690 27430
rect 18750 27370 18760 27430
rect 18680 27360 18760 27370
rect 18850 27430 18910 27440
rect 18850 27360 18910 27370
rect 18940 27810 19110 27840
rect 19140 27880 19200 27890
rect 19140 27810 19200 27820
rect 18940 27360 18970 27810
rect 19260 27780 19290 30450
rect 19350 27830 19380 30590
rect 22130 30600 22140 30660
rect 22200 30600 22210 30660
rect 22130 30590 22210 30600
rect 19060 27750 19290 27780
rect 19320 27820 19380 27830
rect 19320 27750 19380 27760
rect 21770 30380 21850 30390
rect 21770 30320 21780 30380
rect 21840 30320 21850 30380
rect 21770 30310 21850 30320
rect 19060 27360 19090 27750
rect 21770 27710 21800 30310
rect 21830 30240 21910 30250
rect 21830 30180 21840 30240
rect 21900 30180 21910 30240
rect 21830 30170 21910 30180
rect 21770 27700 21830 27710
rect 21770 27630 21830 27640
rect 21860 27660 21890 30170
rect 21950 30100 22030 30110
rect 21950 30040 21960 30100
rect 22020 30040 22030 30100
rect 21950 30030 22030 30040
rect 21950 27770 21980 30030
rect 22010 29960 22090 29970
rect 22010 29900 22020 29960
rect 22080 29900 22090 29960
rect 22010 29890 22090 29900
rect 21950 27760 22010 27770
rect 21950 27690 22010 27700
rect 22040 27720 22070 29890
rect 22130 27830 22160 30590
rect 22190 30520 22270 30530
rect 22190 30460 22200 30520
rect 22260 30460 22270 30520
rect 22190 30450 22270 30460
rect 22130 27820 22190 27830
rect 22130 27750 22190 27760
rect 22220 27780 22250 30450
rect 22310 27890 22340 30870
rect 22370 30800 22450 30810
rect 22370 30740 22380 30800
rect 22440 30740 22450 30800
rect 22370 30730 22450 30740
rect 24050 30730 24060 30790
rect 24120 30730 24130 30790
rect 22310 27880 22370 27890
rect 22310 27810 22370 27820
rect 22400 27840 22430 30730
rect 23670 28420 23750 28430
rect 23670 28360 23680 28420
rect 23740 28360 23750 28420
rect 23670 28350 23750 28360
rect 23820 28350 23830 28410
rect 23890 28350 23900 28410
rect 22600 28280 22680 28290
rect 22600 28220 22610 28280
rect 22670 28220 22680 28280
rect 22600 28210 22680 28220
rect 22400 27810 22570 27840
rect 22220 27750 22450 27780
rect 22040 27690 22330 27720
rect 21860 27630 22210 27660
rect 22180 27360 22210 27630
rect 22300 27360 22330 27690
rect 22420 27360 22450 27750
rect 22540 27360 22570 27810
rect 22600 27430 22670 28210
rect 23680 27440 23750 28350
rect 23870 27440 23900 28350
rect 24070 27840 24100 30730
rect 24160 27890 24190 30870
rect 27300 30880 27310 30940
rect 27370 30880 27380 30940
rect 32290 30940 32370 30950
rect 27300 30870 27380 30880
rect 29100 30870 29110 30930
rect 29170 30870 29180 30930
rect 27120 30660 27200 30670
rect 24290 30590 24300 30650
rect 24360 30590 24370 30650
rect 24230 30450 24240 30510
rect 24300 30450 24310 30510
rect 23670 27430 23750 27440
rect 22600 27370 22610 27430
rect 22670 27370 22680 27430
rect 22600 27360 22680 27370
rect 23670 27370 23680 27430
rect 23740 27370 23750 27430
rect 23670 27360 23750 27370
rect 23840 27430 23900 27440
rect 23840 27360 23900 27370
rect 23930 27810 24100 27840
rect 24130 27880 24190 27890
rect 24130 27810 24190 27820
rect 23930 27360 23960 27810
rect 24250 27780 24280 30450
rect 24340 27830 24370 30590
rect 27120 30600 27130 30660
rect 27190 30600 27200 30660
rect 27120 30590 27200 30600
rect 26760 30380 26840 30390
rect 24650 30310 24660 30370
rect 24720 30310 24730 30370
rect 24590 30170 24600 30230
rect 24660 30170 24670 30230
rect 24470 30030 24480 30090
rect 24540 30030 24550 30090
rect 24410 29890 24420 29950
rect 24480 29890 24490 29950
rect 24050 27750 24280 27780
rect 24310 27820 24370 27830
rect 24310 27750 24370 27760
rect 24050 27360 24080 27750
rect 24430 27720 24460 29890
rect 24520 27770 24550 30030
rect 24170 27690 24460 27720
rect 24490 27760 24550 27770
rect 24490 27690 24550 27700
rect 24170 27360 24200 27690
rect 24610 27660 24640 30170
rect 24700 27710 24730 30310
rect 24290 27630 24640 27660
rect 24670 27700 24730 27710
rect 24670 27630 24730 27640
rect 26760 30320 26770 30380
rect 26830 30320 26840 30380
rect 26760 30310 26840 30320
rect 26760 27710 26790 30310
rect 26820 30240 26900 30250
rect 26820 30180 26830 30240
rect 26890 30180 26900 30240
rect 26820 30170 26900 30180
rect 26760 27700 26820 27710
rect 26760 27630 26820 27640
rect 26850 27660 26880 30170
rect 26940 30100 27020 30110
rect 26940 30040 26950 30100
rect 27010 30040 27020 30100
rect 26940 30030 27020 30040
rect 26940 27770 26970 30030
rect 27000 29960 27080 29970
rect 27000 29900 27010 29960
rect 27070 29900 27080 29960
rect 27000 29890 27080 29900
rect 26940 27760 27000 27770
rect 26940 27690 27000 27700
rect 27030 27720 27060 29890
rect 27120 27830 27150 30590
rect 27180 30520 27260 30530
rect 27180 30460 27190 30520
rect 27250 30460 27260 30520
rect 27180 30450 27260 30460
rect 27120 27820 27180 27830
rect 27120 27750 27180 27760
rect 27210 27780 27240 30450
rect 27300 27890 27330 30870
rect 27360 30800 27440 30810
rect 27360 30740 27370 30800
rect 27430 30740 27440 30800
rect 27360 30730 27440 30740
rect 29040 30730 29050 30790
rect 29110 30730 29120 30790
rect 27300 27880 27360 27890
rect 27300 27810 27360 27820
rect 27390 27840 27420 30730
rect 28660 28420 28740 28430
rect 28660 28360 28670 28420
rect 28730 28360 28740 28420
rect 28660 28350 28740 28360
rect 28810 28350 28820 28410
rect 28880 28350 28890 28410
rect 27590 28280 27670 28290
rect 27590 28220 27600 28280
rect 27660 28220 27670 28280
rect 27590 28210 27670 28220
rect 27390 27810 27560 27840
rect 27210 27750 27440 27780
rect 27030 27690 27320 27720
rect 26850 27630 27200 27660
rect 24290 27360 24320 27630
rect 27170 27360 27200 27630
rect 27290 27360 27320 27690
rect 27410 27360 27440 27750
rect 27530 27360 27560 27810
rect 27590 27430 27660 28210
rect 28670 27440 28740 28350
rect 28860 27440 28890 28350
rect 29060 27840 29090 30730
rect 29150 27890 29180 30870
rect 32290 30880 32300 30940
rect 32360 30880 32370 30940
rect 37280 30940 37360 30950
rect 32290 30870 32370 30880
rect 34090 30870 34100 30930
rect 34160 30870 34170 30930
rect 32110 30660 32190 30670
rect 29280 30590 29290 30650
rect 29350 30590 29360 30650
rect 29220 30450 29230 30510
rect 29290 30450 29300 30510
rect 28660 27430 28740 27440
rect 27590 27370 27600 27430
rect 27660 27370 27670 27430
rect 27590 27360 27670 27370
rect 28660 27370 28670 27430
rect 28730 27370 28740 27430
rect 28660 27360 28740 27370
rect 28830 27430 28890 27440
rect 28830 27360 28890 27370
rect 28920 27810 29090 27840
rect 29120 27880 29180 27890
rect 29120 27810 29180 27820
rect 28920 27360 28950 27810
rect 29240 27780 29270 30450
rect 29330 27830 29360 30590
rect 32110 30600 32120 30660
rect 32180 30600 32190 30660
rect 32110 30590 32190 30600
rect 31930 30380 32010 30390
rect 29640 30310 29650 30370
rect 29710 30310 29720 30370
rect 29580 30170 29590 30230
rect 29650 30170 29660 30230
rect 29460 30030 29470 30090
rect 29530 30030 29540 30090
rect 29400 29890 29410 29950
rect 29470 29890 29480 29950
rect 29040 27750 29270 27780
rect 29300 27820 29360 27830
rect 29300 27750 29360 27760
rect 29040 27360 29070 27750
rect 29420 27720 29450 29890
rect 29510 27770 29540 30030
rect 29160 27690 29450 27720
rect 29480 27760 29540 27770
rect 29480 27690 29540 27700
rect 29160 27360 29190 27690
rect 29600 27660 29630 30170
rect 29690 27710 29720 30310
rect 31930 30320 31940 30380
rect 32000 30320 32010 30380
rect 31930 30310 32010 30320
rect 31750 30100 31830 30110
rect 31750 30040 31760 30100
rect 31820 30040 31830 30100
rect 31750 30030 31830 30040
rect 29280 27630 29630 27660
rect 29660 27700 29720 27710
rect 29660 27630 29720 27640
rect 31390 29820 31470 29830
rect 31390 29760 31400 29820
rect 31460 29760 31470 29820
rect 31390 29750 31470 29760
rect 29280 27360 29310 27630
rect 31390 27590 31420 29750
rect 31450 29680 31530 29690
rect 31450 29620 31460 29680
rect 31520 29620 31530 29680
rect 31450 29610 31530 29620
rect 31390 27580 31450 27590
rect 31390 27510 31450 27520
rect 31480 27540 31510 29610
rect 31570 29540 31650 29550
rect 31570 29480 31580 29540
rect 31640 29480 31650 29540
rect 31570 29470 31650 29480
rect 31570 27650 31600 29470
rect 31630 29400 31710 29410
rect 31630 29340 31640 29400
rect 31700 29340 31710 29400
rect 31630 29330 31710 29340
rect 31570 27640 31630 27650
rect 31570 27570 31630 27580
rect 31660 27600 31690 29330
rect 31750 27710 31780 30030
rect 31810 29960 31890 29970
rect 31810 29900 31820 29960
rect 31880 29900 31890 29960
rect 31810 29890 31890 29900
rect 31750 27700 31810 27710
rect 31750 27630 31810 27640
rect 31840 27660 31870 29890
rect 31930 27770 31960 30310
rect 31990 30240 32070 30250
rect 31990 30180 32000 30240
rect 32060 30180 32070 30240
rect 31990 30170 32070 30180
rect 31930 27760 31990 27770
rect 31930 27690 31990 27700
rect 32020 27720 32050 30170
rect 32110 27830 32140 30590
rect 32170 30520 32250 30530
rect 32170 30460 32180 30520
rect 32240 30460 32250 30520
rect 32170 30450 32250 30460
rect 32110 27820 32170 27830
rect 32110 27750 32170 27760
rect 32200 27780 32230 30450
rect 32290 27890 32320 30870
rect 32350 30800 32430 30810
rect 32350 30740 32360 30800
rect 32420 30740 32430 30800
rect 32350 30730 32430 30740
rect 34030 30730 34040 30790
rect 34100 30730 34110 30790
rect 32290 27880 32350 27890
rect 32290 27810 32350 27820
rect 32380 27840 32410 30730
rect 33650 28420 33730 28430
rect 33650 28360 33660 28420
rect 33720 28360 33730 28420
rect 33650 28350 33730 28360
rect 33800 28350 33810 28410
rect 33870 28350 33880 28410
rect 32580 28280 32660 28290
rect 32580 28220 32590 28280
rect 32650 28220 32660 28280
rect 32580 28210 32660 28220
rect 32380 27810 32550 27840
rect 32200 27750 32430 27780
rect 32020 27690 32310 27720
rect 31840 27630 32190 27660
rect 31660 27570 32070 27600
rect 31480 27510 31950 27540
rect 31920 27360 31950 27510
rect 32040 27360 32070 27570
rect 32160 27360 32190 27630
rect 32280 27360 32310 27690
rect 32400 27360 32430 27750
rect 32520 27360 32550 27810
rect 32580 27430 32650 28210
rect 33660 27440 33730 28350
rect 33850 27440 33880 28350
rect 34050 27840 34080 30730
rect 34140 27890 34170 30870
rect 37280 30880 37290 30940
rect 37350 30880 37360 30940
rect 42270 30940 42350 30950
rect 37280 30870 37360 30880
rect 39080 30870 39090 30930
rect 39150 30870 39160 30930
rect 37100 30660 37180 30670
rect 34270 30590 34280 30650
rect 34340 30590 34350 30650
rect 34210 30450 34220 30510
rect 34280 30450 34290 30510
rect 33650 27430 33730 27440
rect 32580 27370 32590 27430
rect 32650 27370 32660 27430
rect 32580 27360 32660 27370
rect 33650 27370 33660 27430
rect 33720 27370 33730 27430
rect 33650 27360 33730 27370
rect 33820 27430 33880 27440
rect 33820 27360 33880 27370
rect 33910 27810 34080 27840
rect 34110 27880 34170 27890
rect 34110 27810 34170 27820
rect 33910 27360 33940 27810
rect 34230 27780 34260 30450
rect 34320 27830 34350 30590
rect 37100 30600 37110 30660
rect 37170 30600 37180 30660
rect 37100 30590 37180 30600
rect 36920 30380 37000 30390
rect 34450 30310 34460 30370
rect 34520 30310 34530 30370
rect 34390 30170 34400 30230
rect 34460 30170 34470 30230
rect 34030 27750 34260 27780
rect 34290 27820 34350 27830
rect 34290 27750 34350 27760
rect 34030 27360 34060 27750
rect 34410 27720 34440 30170
rect 34500 27770 34530 30310
rect 36920 30320 36930 30380
rect 36990 30320 37000 30380
rect 36920 30310 37000 30320
rect 36740 30100 36820 30110
rect 34630 30030 34640 30090
rect 34700 30030 34710 30090
rect 34570 29890 34580 29950
rect 34640 29890 34650 29950
rect 34150 27690 34440 27720
rect 34470 27760 34530 27770
rect 34470 27690 34530 27700
rect 34150 27360 34180 27690
rect 34590 27660 34620 29890
rect 34680 27710 34710 30030
rect 36740 30040 36750 30100
rect 36810 30040 36820 30100
rect 36740 30030 36820 30040
rect 36560 29820 36640 29830
rect 34990 29750 35000 29810
rect 35060 29750 35070 29810
rect 34930 29610 34940 29670
rect 35000 29610 35010 29670
rect 34810 29470 34820 29530
rect 34880 29470 34890 29530
rect 34750 29330 34760 29390
rect 34820 29330 34830 29390
rect 34270 27630 34620 27660
rect 34650 27700 34710 27710
rect 34650 27630 34710 27640
rect 34270 27360 34300 27630
rect 34770 27600 34800 29330
rect 34860 27650 34890 29470
rect 34390 27570 34800 27600
rect 34830 27640 34890 27650
rect 34830 27570 34890 27580
rect 34390 27360 34420 27570
rect 34950 27540 34980 29610
rect 35040 27590 35070 29750
rect 36560 29760 36570 29820
rect 36630 29760 36640 29820
rect 36560 29750 36640 29760
rect 36380 29260 36460 29270
rect 36380 29200 36390 29260
rect 36450 29200 36460 29260
rect 36380 29190 36460 29200
rect 34510 27510 34980 27540
rect 35010 27580 35070 27590
rect 35010 27510 35070 27520
rect 36200 28700 36280 28710
rect 36200 28640 36210 28700
rect 36270 28640 36280 28700
rect 36200 28630 36280 28640
rect 36200 27530 36230 28630
rect 36260 28560 36340 28570
rect 36260 28500 36270 28560
rect 36330 28500 36340 28560
rect 36260 28490 36340 28500
rect 36200 27520 36260 27530
rect 34510 27360 34540 27510
rect 36200 27450 36260 27460
rect 36290 27480 36320 28490
rect 36380 27590 36410 29190
rect 36440 29120 36520 29130
rect 36440 29060 36450 29120
rect 36510 29060 36520 29120
rect 36440 29050 36520 29060
rect 36380 27580 36440 27590
rect 36380 27510 36440 27520
rect 36470 27540 36500 29050
rect 36560 27650 36590 29750
rect 36620 29680 36700 29690
rect 36620 29620 36630 29680
rect 36690 29620 36700 29680
rect 36620 29610 36700 29620
rect 36560 27640 36620 27650
rect 36560 27570 36620 27580
rect 36650 27600 36680 29610
rect 36740 27710 36770 30030
rect 36800 29960 36880 29970
rect 36800 29900 36810 29960
rect 36870 29900 36880 29960
rect 36800 29890 36880 29900
rect 36740 27700 36800 27710
rect 36740 27630 36800 27640
rect 36830 27660 36860 29890
rect 36920 27770 36950 30310
rect 36980 30240 37060 30250
rect 36980 30180 36990 30240
rect 37050 30180 37060 30240
rect 36980 30170 37060 30180
rect 36920 27760 36980 27770
rect 36920 27690 36980 27700
rect 37010 27720 37040 30170
rect 37100 27830 37130 30590
rect 37160 30520 37240 30530
rect 37160 30460 37170 30520
rect 37230 30460 37240 30520
rect 37160 30450 37240 30460
rect 37100 27820 37160 27830
rect 37100 27750 37160 27760
rect 37190 27780 37220 30450
rect 37280 27890 37310 30870
rect 37340 30800 37420 30810
rect 37340 30740 37350 30800
rect 37410 30740 37420 30800
rect 37340 30730 37420 30740
rect 39020 30730 39030 30790
rect 39090 30730 39100 30790
rect 37280 27880 37340 27890
rect 37280 27810 37340 27820
rect 37370 27840 37400 30730
rect 38640 28420 38720 28430
rect 38640 28360 38650 28420
rect 38710 28360 38720 28420
rect 38640 28350 38720 28360
rect 38790 28350 38800 28410
rect 38860 28350 38870 28410
rect 37570 28280 37650 28290
rect 37570 28220 37580 28280
rect 37640 28220 37650 28280
rect 37570 28210 37650 28220
rect 37370 27810 37540 27840
rect 37190 27750 37420 27780
rect 37010 27690 37300 27720
rect 36830 27630 37180 27660
rect 36650 27570 37060 27600
rect 36470 27510 36940 27540
rect 36290 27450 36820 27480
rect 36790 27360 36820 27450
rect 36910 27360 36940 27510
rect 37030 27360 37060 27570
rect 37150 27360 37180 27630
rect 37270 27360 37300 27690
rect 37390 27360 37420 27750
rect 37510 27360 37540 27810
rect 37570 27430 37640 28210
rect 38650 27440 38720 28350
rect 38840 27440 38870 28350
rect 39040 27840 39070 30730
rect 39130 27890 39160 30870
rect 42270 30880 42280 30940
rect 42340 30880 42350 30940
rect 47260 30940 47340 30950
rect 42270 30870 42350 30880
rect 44070 30870 44080 30930
rect 44140 30870 44150 30930
rect 42090 30660 42170 30670
rect 39260 30590 39270 30650
rect 39330 30590 39340 30650
rect 39200 30450 39210 30510
rect 39270 30450 39280 30510
rect 38640 27430 38720 27440
rect 37570 27370 37580 27430
rect 37640 27370 37650 27430
rect 37570 27360 37650 27370
rect 38640 27370 38650 27430
rect 38710 27370 38720 27430
rect 38640 27360 38720 27370
rect 38810 27430 38870 27440
rect 38810 27360 38870 27370
rect 38900 27810 39070 27840
rect 39100 27880 39160 27890
rect 39100 27810 39160 27820
rect 38900 27360 38930 27810
rect 39220 27780 39250 30450
rect 39310 27830 39340 30590
rect 42090 30600 42100 30660
rect 42160 30600 42170 30660
rect 42090 30590 42170 30600
rect 41910 30380 41990 30390
rect 39440 30310 39450 30370
rect 39510 30310 39520 30370
rect 39380 30170 39390 30230
rect 39450 30170 39460 30230
rect 39020 27750 39250 27780
rect 39280 27820 39340 27830
rect 39280 27750 39340 27760
rect 39020 27360 39050 27750
rect 39400 27720 39430 30170
rect 39490 27770 39520 30310
rect 41910 30320 41920 30380
rect 41980 30320 41990 30380
rect 41910 30310 41990 30320
rect 41730 30100 41810 30110
rect 39620 30030 39630 30090
rect 39690 30030 39700 30090
rect 39560 29890 39570 29950
rect 39630 29890 39640 29950
rect 39140 27690 39430 27720
rect 39460 27760 39520 27770
rect 39460 27690 39520 27700
rect 39140 27360 39170 27690
rect 39580 27660 39610 29890
rect 39670 27710 39700 30030
rect 41730 30040 41740 30100
rect 41800 30040 41810 30100
rect 41730 30030 41810 30040
rect 41550 29820 41630 29830
rect 39800 29750 39810 29810
rect 39870 29750 39880 29810
rect 39740 29610 39750 29670
rect 39810 29610 39820 29670
rect 39260 27630 39610 27660
rect 39640 27700 39700 27710
rect 39640 27630 39700 27640
rect 39260 27360 39290 27630
rect 39760 27600 39790 29610
rect 39850 27650 39880 29750
rect 41550 29760 41560 29820
rect 41620 29760 41630 29820
rect 41550 29750 41630 29760
rect 41190 29260 41270 29270
rect 39980 29190 39990 29250
rect 40050 29190 40060 29250
rect 39920 29050 39930 29110
rect 39990 29050 40000 29110
rect 39380 27570 39790 27600
rect 39820 27640 39880 27650
rect 39820 27570 39880 27580
rect 39380 27360 39410 27570
rect 39940 27540 39970 29050
rect 40030 27590 40060 29190
rect 41190 29200 41200 29260
rect 41260 29200 41270 29260
rect 41190 29190 41270 29200
rect 40160 28630 40170 28690
rect 40230 28630 40240 28690
rect 40090 28490 40100 28550
rect 40160 28490 40170 28550
rect 39500 27510 39970 27540
rect 40000 27580 40060 27590
rect 40000 27510 40060 27520
rect 39500 27360 39530 27510
rect 40120 27480 40150 28490
rect 40210 27530 40240 28630
rect 39620 27450 40150 27480
rect 40180 27520 40240 27530
rect 40180 27450 40240 27460
rect 41190 27530 41220 29190
rect 41250 29120 41330 29130
rect 41250 29060 41260 29120
rect 41320 29060 41330 29120
rect 41250 29050 41330 29060
rect 41190 27520 41250 27530
rect 41190 27450 41250 27460
rect 41280 27480 41310 29050
rect 41340 28980 41420 28990
rect 41340 28920 41350 28980
rect 41410 28920 41420 28980
rect 41340 28910 41420 28920
rect 41370 27590 41400 28910
rect 41430 28840 41510 28850
rect 41430 28780 41440 28840
rect 41500 28780 41510 28840
rect 41430 28770 41510 28780
rect 41370 27580 41430 27590
rect 41370 27510 41430 27520
rect 41460 27540 41490 28770
rect 41550 27650 41580 29750
rect 41610 29680 41690 29690
rect 41610 29620 41620 29680
rect 41680 29620 41690 29680
rect 41610 29610 41690 29620
rect 41550 27640 41610 27650
rect 41550 27570 41610 27580
rect 41640 27600 41670 29610
rect 41730 27710 41760 30030
rect 41790 29960 41870 29970
rect 41790 29900 41800 29960
rect 41860 29900 41870 29960
rect 41790 29890 41870 29900
rect 41730 27700 41790 27710
rect 41730 27630 41790 27640
rect 41820 27660 41850 29890
rect 41910 27770 41940 30310
rect 41970 30240 42050 30250
rect 41970 30180 41980 30240
rect 42040 30180 42050 30240
rect 41970 30170 42050 30180
rect 41910 27760 41970 27770
rect 41910 27690 41970 27700
rect 42000 27720 42030 30170
rect 42090 27830 42120 30590
rect 42150 30520 42230 30530
rect 42150 30460 42160 30520
rect 42220 30460 42230 30520
rect 42150 30450 42230 30460
rect 42090 27820 42150 27830
rect 42090 27750 42150 27760
rect 42180 27780 42210 30450
rect 42270 27890 42300 30870
rect 42330 30800 42410 30810
rect 42330 30740 42340 30800
rect 42400 30740 42410 30800
rect 42330 30730 42410 30740
rect 44010 30730 44020 30790
rect 44080 30730 44090 30790
rect 42270 27880 42330 27890
rect 42270 27810 42330 27820
rect 42360 27840 42390 30730
rect 43630 28420 43710 28430
rect 43630 28360 43640 28420
rect 43700 28360 43710 28420
rect 43630 28350 43710 28360
rect 43780 28350 43790 28410
rect 43850 28350 43860 28410
rect 42560 28280 42640 28290
rect 42560 28220 42570 28280
rect 42630 28220 42640 28280
rect 42560 28210 42640 28220
rect 42360 27810 42530 27840
rect 42180 27750 42410 27780
rect 42000 27690 42290 27720
rect 41820 27630 42170 27660
rect 41640 27570 42050 27600
rect 41460 27510 41930 27540
rect 41280 27450 41810 27480
rect 39620 27360 39650 27450
rect 41780 27360 41810 27450
rect 41900 27360 41930 27510
rect 42020 27360 42050 27570
rect 42140 27360 42170 27630
rect 42260 27360 42290 27690
rect 42380 27360 42410 27750
rect 42500 27360 42530 27810
rect 42560 27430 42630 28210
rect 43640 27440 43710 28350
rect 43830 27440 43860 28350
rect 44030 27840 44060 30730
rect 44120 27890 44150 30870
rect 47260 30880 47270 30940
rect 47330 30880 47340 30940
rect 52250 30940 52330 30950
rect 47260 30870 47340 30880
rect 49060 30870 49070 30930
rect 49130 30870 49140 30930
rect 47080 30660 47160 30670
rect 44250 30590 44260 30650
rect 44320 30590 44330 30650
rect 44190 30450 44200 30510
rect 44260 30450 44270 30510
rect 43630 27430 43710 27440
rect 42560 27370 42570 27430
rect 42630 27370 42640 27430
rect 42560 27360 42640 27370
rect 43630 27370 43640 27430
rect 43700 27370 43710 27430
rect 43630 27360 43710 27370
rect 43800 27430 43860 27440
rect 43800 27360 43860 27370
rect 43890 27810 44060 27840
rect 44090 27880 44150 27890
rect 44090 27810 44150 27820
rect 43890 27360 43920 27810
rect 44210 27780 44240 30450
rect 44300 27830 44330 30590
rect 47080 30600 47090 30660
rect 47150 30600 47160 30660
rect 47080 30590 47160 30600
rect 46900 30380 46980 30390
rect 44430 30310 44440 30370
rect 44500 30310 44510 30370
rect 44370 30170 44380 30230
rect 44440 30170 44450 30230
rect 44010 27750 44240 27780
rect 44270 27820 44330 27830
rect 44270 27750 44330 27760
rect 44010 27360 44040 27750
rect 44390 27720 44420 30170
rect 44480 27770 44510 30310
rect 46900 30320 46910 30380
rect 46970 30320 46980 30380
rect 46900 30310 46980 30320
rect 46720 30100 46800 30110
rect 44610 30030 44620 30090
rect 44680 30030 44690 30090
rect 44550 29890 44560 29950
rect 44620 29890 44630 29950
rect 44130 27690 44420 27720
rect 44450 27760 44510 27770
rect 44450 27690 44510 27700
rect 44130 27360 44160 27690
rect 44570 27660 44600 29890
rect 44660 27710 44690 30030
rect 46720 30040 46730 30100
rect 46790 30040 46800 30100
rect 46720 30030 46800 30040
rect 46360 29820 46440 29830
rect 44790 29750 44800 29810
rect 44860 29750 44870 29810
rect 44730 29610 44740 29670
rect 44800 29610 44810 29670
rect 44250 27630 44600 27660
rect 44630 27700 44690 27710
rect 44630 27630 44690 27640
rect 44250 27360 44280 27630
rect 44750 27600 44780 29610
rect 44840 27650 44870 29750
rect 46360 29760 46370 29820
rect 46430 29760 46440 29820
rect 46360 29750 46440 29760
rect 45150 29190 45160 29250
rect 45220 29190 45230 29250
rect 45090 29050 45100 29110
rect 45160 29050 45170 29110
rect 45000 28910 45010 28970
rect 45070 28910 45080 28970
rect 44910 28770 44920 28830
rect 44980 28770 44990 28830
rect 44370 27570 44780 27600
rect 44810 27640 44870 27650
rect 44810 27570 44870 27580
rect 44370 27330 44400 27570
rect 44930 27540 44960 28770
rect 45020 27590 45050 28910
rect 44490 27510 44960 27540
rect 44990 27580 45050 27590
rect 44990 27510 45050 27520
rect 44490 27360 44520 27510
rect 45110 27480 45140 29050
rect 45200 27530 45230 29190
rect 44610 27450 45140 27480
rect 45170 27520 45230 27530
rect 46360 27590 46390 29750
rect 46420 29680 46500 29690
rect 46420 29620 46430 29680
rect 46490 29620 46500 29680
rect 46420 29610 46500 29620
rect 46360 27580 46420 27590
rect 46360 27510 46420 27520
rect 46450 27540 46480 29610
rect 46540 29540 46620 29550
rect 46540 29480 46550 29540
rect 46610 29480 46620 29540
rect 46540 29470 46620 29480
rect 46540 27650 46570 29470
rect 46600 29400 46680 29410
rect 46600 29340 46610 29400
rect 46670 29340 46680 29400
rect 46600 29330 46680 29340
rect 46540 27640 46600 27650
rect 46540 27570 46600 27580
rect 46630 27600 46660 29330
rect 46720 27710 46750 30030
rect 46780 29960 46860 29970
rect 46780 29900 46790 29960
rect 46850 29900 46860 29960
rect 46780 29890 46860 29900
rect 46720 27700 46780 27710
rect 46720 27630 46780 27640
rect 46810 27660 46840 29890
rect 46900 27770 46930 30310
rect 46960 30240 47040 30250
rect 46960 30180 46970 30240
rect 47030 30180 47040 30240
rect 46960 30170 47040 30180
rect 46900 27760 46960 27770
rect 46900 27690 46960 27700
rect 46990 27720 47020 30170
rect 47080 27830 47110 30590
rect 47140 30520 47220 30530
rect 47140 30460 47150 30520
rect 47210 30460 47220 30520
rect 47140 30450 47220 30460
rect 47080 27820 47140 27830
rect 47080 27750 47140 27760
rect 47170 27780 47200 30450
rect 47260 27890 47290 30870
rect 47320 30800 47400 30810
rect 47320 30740 47330 30800
rect 47390 30740 47400 30800
rect 47320 30730 47400 30740
rect 49000 30730 49010 30790
rect 49070 30730 49080 30790
rect 47260 27880 47320 27890
rect 47260 27810 47320 27820
rect 47350 27840 47380 30730
rect 48620 28420 48700 28430
rect 48620 28360 48630 28420
rect 48690 28360 48700 28420
rect 48620 28350 48700 28360
rect 48770 28350 48780 28410
rect 48840 28350 48850 28410
rect 47550 28280 47630 28290
rect 47550 28220 47560 28280
rect 47620 28220 47630 28280
rect 47550 28210 47630 28220
rect 47350 27810 47520 27840
rect 47170 27750 47400 27780
rect 46990 27690 47280 27720
rect 46810 27630 47160 27660
rect 46630 27570 47040 27600
rect 46450 27510 46920 27540
rect 45170 27450 45230 27460
rect 44610 27360 44640 27450
rect 46890 27360 46920 27510
rect 47010 27360 47040 27570
rect 47130 27360 47160 27630
rect 47250 27360 47280 27690
rect 47370 27360 47400 27750
rect 47490 27360 47520 27810
rect 47550 27430 47620 28210
rect 48630 27440 48700 28350
rect 48820 27440 48850 28350
rect 49020 27840 49050 30730
rect 49110 27890 49140 30870
rect 52250 30880 52260 30940
rect 52320 30880 52330 30940
rect 57240 30940 57320 30950
rect 52250 30870 52330 30880
rect 54050 30870 54060 30930
rect 54120 30870 54130 30930
rect 52070 30660 52150 30670
rect 49240 30590 49250 30650
rect 49310 30590 49320 30650
rect 49180 30450 49190 30510
rect 49250 30450 49260 30510
rect 48620 27430 48700 27440
rect 47550 27370 47560 27430
rect 47620 27370 47630 27430
rect 47550 27360 47630 27370
rect 48620 27370 48630 27430
rect 48690 27370 48700 27430
rect 48620 27360 48700 27370
rect 48790 27430 48850 27440
rect 48790 27360 48850 27370
rect 48880 27810 49050 27840
rect 49080 27880 49140 27890
rect 49080 27810 49140 27820
rect 48880 27360 48910 27810
rect 49200 27780 49230 30450
rect 49290 27830 49320 30590
rect 52070 30600 52080 30660
rect 52140 30600 52150 30660
rect 52070 30590 52150 30600
rect 51710 30380 51790 30390
rect 49420 30310 49430 30370
rect 49490 30310 49500 30370
rect 49360 30170 49370 30230
rect 49430 30170 49440 30230
rect 49000 27750 49230 27780
rect 49260 27820 49320 27830
rect 49260 27750 49320 27760
rect 49000 27360 49030 27750
rect 49380 27720 49410 30170
rect 49470 27770 49500 30310
rect 51710 30320 51720 30380
rect 51780 30320 51790 30380
rect 51710 30310 51790 30320
rect 49600 30030 49610 30090
rect 49670 30030 49680 30090
rect 49540 29890 49550 29950
rect 49610 29890 49620 29950
rect 49120 27690 49410 27720
rect 49440 27760 49500 27770
rect 49440 27690 49500 27700
rect 49120 27360 49150 27690
rect 49560 27660 49590 29890
rect 49650 27710 49680 30030
rect 49960 29750 49970 29810
rect 50030 29750 50040 29810
rect 49900 29610 49910 29670
rect 49970 29610 49980 29670
rect 49780 29470 49790 29530
rect 49850 29470 49860 29530
rect 49720 29330 49730 29390
rect 49790 29330 49800 29390
rect 49240 27630 49590 27660
rect 49620 27700 49680 27710
rect 49620 27630 49680 27640
rect 49240 27360 49270 27630
rect 49740 27600 49770 29330
rect 49830 27650 49860 29470
rect 49360 27570 49770 27600
rect 49800 27640 49860 27650
rect 49800 27570 49860 27580
rect 49360 27360 49390 27570
rect 49920 27540 49950 29610
rect 50010 27590 50040 29750
rect 51710 27710 51740 30310
rect 51770 30240 51850 30250
rect 51770 30180 51780 30240
rect 51840 30180 51850 30240
rect 51770 30170 51850 30180
rect 51710 27700 51770 27710
rect 51710 27630 51770 27640
rect 51800 27660 51830 30170
rect 51890 30100 51970 30110
rect 51890 30040 51900 30100
rect 51960 30040 51970 30100
rect 51890 30030 51970 30040
rect 51890 27770 51920 30030
rect 51950 29960 52030 29970
rect 51950 29900 51960 29960
rect 52020 29900 52030 29960
rect 51950 29890 52030 29900
rect 51890 27760 51950 27770
rect 51890 27690 51950 27700
rect 51980 27720 52010 29890
rect 52070 27830 52100 30590
rect 52130 30520 52210 30530
rect 52130 30460 52140 30520
rect 52200 30460 52210 30520
rect 52130 30450 52210 30460
rect 52070 27820 52130 27830
rect 52070 27750 52130 27760
rect 52160 27780 52190 30450
rect 52250 27890 52280 30870
rect 52310 30800 52390 30810
rect 52310 30740 52320 30800
rect 52380 30740 52390 30800
rect 52310 30730 52390 30740
rect 53990 30730 54000 30790
rect 54060 30730 54070 30790
rect 52250 27880 52310 27890
rect 52250 27810 52310 27820
rect 52340 27840 52370 30730
rect 53610 28420 53690 28430
rect 53610 28360 53620 28420
rect 53680 28360 53690 28420
rect 53610 28350 53690 28360
rect 53760 28350 53770 28410
rect 53830 28350 53840 28410
rect 52540 28280 52620 28290
rect 52540 28220 52550 28280
rect 52610 28220 52620 28280
rect 52540 28210 52620 28220
rect 52340 27810 52510 27840
rect 52160 27750 52390 27780
rect 51980 27690 52270 27720
rect 51800 27630 52150 27660
rect 49480 27510 49950 27540
rect 49980 27580 50040 27590
rect 49980 27510 50040 27520
rect 49480 27360 49510 27510
rect 52120 27360 52150 27630
rect 52240 27360 52270 27690
rect 52360 27360 52390 27750
rect 52480 27360 52510 27810
rect 52540 27430 52610 28210
rect 53620 27440 53690 28350
rect 53810 27440 53840 28350
rect 54010 27840 54040 30730
rect 54100 27890 54130 30870
rect 57240 30880 57250 30940
rect 57310 30880 57320 30940
rect 62230 30940 62310 30950
rect 57240 30870 57320 30880
rect 59040 30870 59050 30930
rect 59110 30870 59120 30930
rect 57060 30660 57140 30670
rect 54230 30590 54240 30650
rect 54300 30590 54310 30650
rect 54170 30450 54180 30510
rect 54240 30450 54250 30510
rect 53610 27430 53690 27440
rect 52540 27370 52550 27430
rect 52610 27370 52620 27430
rect 52540 27360 52620 27370
rect 53610 27370 53620 27430
rect 53680 27370 53690 27430
rect 53610 27360 53690 27370
rect 53780 27430 53840 27440
rect 53780 27360 53840 27370
rect 53870 27810 54040 27840
rect 54070 27880 54130 27890
rect 54070 27810 54130 27820
rect 53870 27360 53900 27810
rect 54190 27780 54220 30450
rect 54280 27830 54310 30590
rect 57060 30600 57070 30660
rect 57130 30600 57140 30660
rect 57060 30590 57140 30600
rect 56700 30380 56780 30390
rect 54590 30310 54600 30370
rect 54660 30310 54670 30370
rect 54530 30170 54540 30230
rect 54600 30170 54610 30230
rect 54410 30030 54420 30090
rect 54480 30030 54490 30090
rect 54350 29890 54360 29950
rect 54420 29890 54430 29950
rect 53990 27750 54220 27780
rect 54250 27820 54310 27830
rect 54250 27750 54310 27760
rect 53990 27360 54020 27750
rect 54370 27720 54400 29890
rect 54460 27770 54490 30030
rect 54110 27690 54400 27720
rect 54430 27760 54490 27770
rect 54430 27690 54490 27700
rect 54110 27360 54140 27690
rect 54550 27660 54580 30170
rect 54640 27710 54670 30310
rect 54230 27630 54580 27660
rect 54610 27700 54670 27710
rect 54610 27630 54670 27640
rect 56700 30320 56710 30380
rect 56770 30320 56780 30380
rect 56700 30310 56780 30320
rect 56700 27710 56730 30310
rect 56760 30240 56840 30250
rect 56760 30180 56770 30240
rect 56830 30180 56840 30240
rect 56760 30170 56840 30180
rect 56700 27700 56760 27710
rect 56700 27630 56760 27640
rect 56790 27660 56820 30170
rect 56880 30100 56960 30110
rect 56880 30040 56890 30100
rect 56950 30040 56960 30100
rect 56880 30030 56960 30040
rect 56880 27770 56910 30030
rect 56940 29960 57020 29970
rect 56940 29900 56950 29960
rect 57010 29900 57020 29960
rect 56940 29890 57020 29900
rect 56880 27760 56940 27770
rect 56880 27690 56940 27700
rect 56970 27720 57000 29890
rect 57060 27830 57090 30590
rect 57120 30520 57200 30530
rect 57120 30460 57130 30520
rect 57190 30460 57200 30520
rect 57120 30450 57200 30460
rect 57060 27820 57120 27830
rect 57060 27750 57120 27760
rect 57150 27780 57180 30450
rect 57240 27890 57270 30870
rect 57300 30800 57380 30810
rect 57300 30740 57310 30800
rect 57370 30740 57380 30800
rect 57300 30730 57380 30740
rect 58980 30730 58990 30790
rect 59050 30730 59060 30790
rect 57240 27880 57300 27890
rect 57240 27810 57300 27820
rect 57330 27840 57360 30730
rect 58600 28420 58680 28430
rect 58600 28360 58610 28420
rect 58670 28360 58680 28420
rect 58600 28350 58680 28360
rect 58750 28350 58760 28410
rect 58820 28350 58830 28410
rect 57530 28280 57610 28290
rect 57530 28220 57540 28280
rect 57600 28220 57610 28280
rect 57530 28210 57610 28220
rect 57330 27810 57500 27840
rect 57150 27750 57380 27780
rect 56970 27690 57260 27720
rect 56790 27630 57140 27660
rect 54230 27360 54260 27630
rect 57110 27360 57140 27630
rect 57230 27360 57260 27690
rect 57350 27360 57380 27750
rect 57470 27360 57500 27810
rect 57530 27430 57600 28210
rect 58610 27440 58680 28350
rect 58800 27440 58830 28350
rect 59000 27840 59030 30730
rect 59090 27890 59120 30870
rect 62230 30880 62240 30940
rect 62300 30880 62310 30940
rect 67220 30940 67300 30950
rect 62230 30870 62310 30880
rect 64030 30870 64040 30930
rect 64100 30870 64110 30930
rect 62050 30660 62130 30670
rect 59220 30590 59230 30650
rect 59290 30590 59300 30650
rect 59160 30450 59170 30510
rect 59230 30450 59240 30510
rect 58600 27430 58680 27440
rect 57530 27370 57540 27430
rect 57600 27370 57610 27430
rect 57530 27360 57610 27370
rect 58600 27370 58610 27430
rect 58670 27370 58680 27430
rect 58600 27360 58680 27370
rect 58770 27430 58830 27440
rect 58770 27360 58830 27370
rect 58860 27810 59030 27840
rect 59060 27880 59120 27890
rect 59060 27810 59120 27820
rect 58860 27360 58890 27810
rect 59180 27780 59210 30450
rect 59270 27830 59300 30590
rect 62050 30600 62060 30660
rect 62120 30600 62130 30660
rect 62050 30590 62130 30600
rect 59580 30310 59590 30370
rect 59650 30310 59660 30370
rect 59520 30170 59530 30230
rect 59590 30170 59600 30230
rect 59400 30030 59410 30090
rect 59470 30030 59480 30090
rect 59340 29890 59350 29950
rect 59410 29890 59420 29950
rect 58980 27750 59210 27780
rect 59240 27820 59300 27830
rect 59240 27750 59300 27760
rect 58980 27360 59010 27750
rect 59360 27720 59390 29890
rect 59450 27770 59480 30030
rect 59100 27690 59390 27720
rect 59420 27760 59480 27770
rect 59420 27690 59480 27700
rect 59100 27360 59130 27690
rect 59540 27660 59570 30170
rect 59630 27710 59660 30310
rect 62050 27830 62080 30590
rect 62110 30520 62190 30530
rect 62110 30460 62120 30520
rect 62180 30460 62190 30520
rect 62110 30450 62190 30460
rect 62050 27820 62110 27830
rect 62050 27750 62110 27760
rect 62140 27780 62170 30450
rect 62230 27890 62260 30870
rect 62290 30800 62370 30810
rect 62290 30740 62300 30800
rect 62360 30740 62370 30800
rect 62290 30730 62370 30740
rect 63970 30730 63980 30790
rect 64040 30730 64050 30790
rect 62230 27880 62290 27890
rect 62230 27810 62290 27820
rect 62320 27840 62350 30730
rect 63590 28420 63670 28430
rect 63590 28360 63600 28420
rect 63660 28360 63670 28420
rect 63590 28350 63670 28360
rect 63740 28350 63750 28410
rect 63810 28350 63820 28410
rect 62520 28280 62600 28290
rect 62520 28220 62530 28280
rect 62590 28220 62600 28280
rect 62520 28210 62600 28220
rect 62320 27810 62490 27840
rect 62140 27750 62370 27780
rect 59220 27630 59570 27660
rect 59600 27700 59660 27710
rect 59600 27630 59660 27640
rect 59220 27360 59250 27630
rect 62340 27360 62370 27750
rect 62460 27360 62490 27810
rect 62520 27430 62590 28210
rect 63600 27440 63670 28350
rect 63790 27440 63820 28350
rect 63990 27840 64020 30730
rect 64080 27890 64110 30870
rect 67220 30880 67230 30940
rect 67290 30880 67300 30940
rect 72210 30940 72290 30950
rect 67220 30870 67300 30880
rect 69020 30870 69030 30930
rect 69090 30870 69100 30930
rect 67040 30660 67120 30670
rect 64210 30590 64220 30650
rect 64280 30590 64290 30650
rect 64150 30450 64160 30510
rect 64220 30450 64230 30510
rect 63590 27430 63670 27440
rect 62520 27370 62530 27430
rect 62590 27370 62600 27430
rect 62520 27360 62600 27370
rect 63590 27370 63600 27430
rect 63660 27370 63670 27430
rect 63590 27360 63670 27370
rect 63760 27430 63820 27440
rect 63760 27360 63820 27370
rect 63850 27810 64020 27840
rect 64050 27880 64110 27890
rect 64050 27810 64110 27820
rect 63850 27360 63880 27810
rect 64170 27780 64200 30450
rect 64260 27830 64290 30590
rect 63970 27750 64200 27780
rect 64230 27820 64290 27830
rect 64230 27750 64290 27760
rect 67040 30600 67050 30660
rect 67110 30600 67120 30660
rect 67040 30590 67120 30600
rect 67040 27830 67070 30590
rect 67100 30520 67180 30530
rect 67100 30460 67110 30520
rect 67170 30460 67180 30520
rect 67100 30450 67180 30460
rect 67040 27820 67100 27830
rect 67040 27750 67100 27760
rect 67130 27780 67160 30450
rect 67220 27890 67250 30870
rect 67280 30800 67360 30810
rect 67280 30740 67290 30800
rect 67350 30740 67360 30800
rect 67280 30730 67360 30740
rect 68960 30730 68970 30790
rect 69030 30730 69040 30790
rect 67220 27880 67280 27890
rect 67220 27810 67280 27820
rect 67310 27840 67340 30730
rect 68580 28420 68660 28430
rect 68580 28360 68590 28420
rect 68650 28360 68660 28420
rect 68580 28350 68660 28360
rect 68730 28350 68740 28410
rect 68800 28350 68810 28410
rect 67510 28280 67590 28290
rect 67510 28220 67520 28280
rect 67580 28220 67590 28280
rect 67510 28210 67590 28220
rect 67310 27810 67480 27840
rect 67130 27750 67360 27780
rect 63970 27360 64000 27750
rect 67330 27360 67360 27750
rect 67450 27360 67480 27810
rect 67510 27430 67580 28210
rect 68590 27440 68660 28350
rect 68780 27440 68810 28350
rect 68980 27840 69010 30730
rect 69070 27890 69100 30870
rect 72210 30880 72220 30940
rect 72280 30880 72290 30940
rect 77200 30940 77280 30950
rect 72210 30870 72290 30880
rect 74010 30870 74020 30930
rect 74080 30870 74090 30930
rect 69200 30590 69210 30650
rect 69270 30590 69280 30650
rect 69140 30450 69150 30510
rect 69210 30450 69220 30510
rect 68580 27430 68660 27440
rect 67510 27370 67520 27430
rect 67580 27370 67590 27430
rect 67510 27360 67590 27370
rect 68580 27370 68590 27430
rect 68650 27370 68660 27430
rect 68580 27360 68660 27370
rect 68750 27430 68810 27440
rect 68750 27360 68810 27370
rect 68840 27810 69010 27840
rect 69040 27880 69100 27890
rect 69040 27810 69100 27820
rect 68840 27360 68870 27810
rect 69160 27780 69190 30450
rect 69250 27830 69280 30590
rect 68960 27750 69190 27780
rect 69220 27820 69280 27830
rect 72210 27890 72240 30870
rect 72270 30800 72350 30810
rect 72270 30740 72280 30800
rect 72340 30740 72350 30800
rect 72270 30730 72350 30740
rect 73950 30730 73960 30790
rect 74020 30730 74030 30790
rect 72210 27880 72270 27890
rect 72210 27810 72270 27820
rect 72300 27840 72330 30730
rect 73570 28420 73650 28430
rect 73570 28360 73580 28420
rect 73640 28360 73650 28420
rect 73570 28350 73650 28360
rect 73720 28350 73730 28410
rect 73790 28350 73800 28410
rect 72500 28280 72580 28290
rect 72500 28220 72510 28280
rect 72570 28220 72580 28280
rect 72500 28210 72580 28220
rect 72300 27810 72470 27840
rect 69220 27750 69280 27760
rect 68960 27360 68990 27750
rect 72440 27360 72470 27810
rect 72500 27430 72570 28210
rect 73580 27440 73650 28350
rect 73770 27440 73800 28350
rect 73970 27840 74000 30730
rect 74060 27890 74090 30870
rect 73570 27430 73650 27440
rect 72500 27370 72510 27430
rect 72570 27370 72580 27430
rect 72500 27360 72580 27370
rect 73570 27370 73580 27430
rect 73640 27370 73650 27430
rect 73570 27360 73650 27370
rect 73740 27430 73800 27440
rect 73740 27360 73800 27370
rect 73830 27810 74000 27840
rect 74030 27880 74090 27890
rect 74030 27810 74090 27820
rect 77200 30880 77210 30940
rect 77270 30880 77280 30940
rect 77200 30870 77280 30880
rect 79000 30870 79010 30930
rect 79070 30870 79080 30930
rect 77200 27890 77230 30870
rect 77260 30800 77340 30810
rect 77260 30740 77270 30800
rect 77330 30740 77340 30800
rect 77260 30730 77340 30740
rect 78940 30730 78950 30790
rect 79010 30730 79020 30790
rect 77200 27880 77260 27890
rect 77200 27810 77260 27820
rect 77290 27840 77320 30730
rect 78560 28420 78640 28430
rect 78560 28360 78570 28420
rect 78630 28360 78640 28420
rect 78560 28350 78640 28360
rect 78710 28350 78720 28410
rect 78780 28350 78790 28410
rect 77490 28280 77570 28290
rect 77490 28220 77500 28280
rect 77560 28220 77570 28280
rect 77490 28210 77570 28220
rect 77290 27810 77460 27840
rect 73830 27360 73860 27810
rect 77430 27360 77460 27810
rect 77490 27430 77560 28210
rect 78570 27440 78640 28350
rect 78760 27440 78790 28350
rect 78960 27840 78990 30730
rect 79050 27890 79080 30870
rect 78560 27430 78640 27440
rect 77490 27370 77500 27430
rect 77560 27370 77570 27430
rect 77490 27360 77570 27370
rect 78560 27370 78570 27430
rect 78630 27370 78640 27430
rect 78560 27360 78640 27370
rect 78730 27430 78790 27440
rect 78730 27360 78790 27370
rect 78820 27810 78990 27840
rect 79020 27880 79080 27890
rect 79020 27810 79080 27820
rect 78820 27360 78850 27810
<< via2 >>
rect 2640 66520 2700 66580
rect 4080 66520 4140 66580
rect 7630 66520 7690 66580
rect 9070 66520 9130 66580
rect 3280 66270 3350 66280
rect 3280 66210 3340 66270
rect 3340 66210 3350 66270
rect 3280 66160 3350 66170
rect 3280 66100 3340 66160
rect 3340 66100 3350 66160
rect 8270 66270 8340 66280
rect 8270 66210 8330 66270
rect 8330 66210 8340 66270
rect 8270 66160 8340 66170
rect 8270 66100 8330 66160
rect 8330 66100 8340 66160
rect 2640 66000 2700 66060
rect 4080 66000 4140 66060
rect 7630 66000 7690 66060
rect 9070 66000 9130 66060
rect 3280 64560 3350 64570
rect 3280 64500 3340 64560
rect 3340 64500 3350 64560
rect 3280 64450 3350 64460
rect 3280 64390 3340 64450
rect 3340 64390 3350 64450
rect 8270 64560 8340 64570
rect 8270 64500 8330 64560
rect 8330 64500 8340 64560
rect 8270 64450 8340 64460
rect 8270 64390 8330 64450
rect 8330 64390 8340 64450
rect 2640 64290 2700 64350
rect 4080 64290 4140 64350
rect 7630 64290 7690 64350
rect 9070 64290 9130 64350
rect 3280 62850 3350 62860
rect 3280 62790 3340 62850
rect 3340 62790 3350 62850
rect 3280 62740 3350 62750
rect 3280 62680 3340 62740
rect 3340 62680 3350 62740
rect 8270 62850 8340 62860
rect 8270 62790 8330 62850
rect 8330 62790 8340 62850
rect 8270 62740 8340 62750
rect 8270 62680 8330 62740
rect 8330 62680 8340 62740
rect 2640 62580 2700 62640
rect 4080 62580 4140 62640
rect 7630 62580 7690 62640
rect 9070 62580 9130 62640
rect 3280 61140 3350 61150
rect 3280 61080 3340 61140
rect 3340 61080 3350 61140
rect 3280 61030 3350 61040
rect 3280 60970 3340 61030
rect 3340 60970 3350 61030
rect 8270 61140 8340 61150
rect 8270 61080 8330 61140
rect 8330 61080 8340 61140
rect 8270 61030 8340 61040
rect 8270 60970 8330 61030
rect 8330 60970 8340 61030
rect 2640 60870 2700 60930
rect 4080 60870 4140 60930
rect 7630 60870 7690 60930
rect 9070 60870 9130 60930
rect 12620 66520 12680 66580
rect 14060 66520 14120 66580
rect 13260 66270 13330 66280
rect 13260 66210 13320 66270
rect 13320 66210 13330 66270
rect 13260 66160 13330 66170
rect 13260 66100 13320 66160
rect 13320 66100 13330 66160
rect 12620 66000 12680 66060
rect 14060 66000 14120 66060
rect 13260 64560 13330 64570
rect 13260 64500 13320 64560
rect 13320 64500 13330 64560
rect 13260 64450 13330 64460
rect 13260 64390 13320 64450
rect 13320 64390 13330 64450
rect 12620 64290 12680 64350
rect 14060 64290 14120 64350
rect 13260 62850 13330 62860
rect 13260 62790 13320 62850
rect 13320 62790 13330 62850
rect 13260 62740 13330 62750
rect 13260 62680 13320 62740
rect 13320 62680 13330 62740
rect 12620 62580 12680 62640
rect 14060 62580 14120 62640
rect 13260 61140 13330 61150
rect 13260 61080 13320 61140
rect 13320 61080 13330 61140
rect 13260 61030 13330 61040
rect 13260 60970 13320 61030
rect 13320 60970 13330 61030
rect 12620 60870 12680 60930
rect 14060 60870 14120 60930
rect 12500 59680 12560 59740
rect 17610 66520 17670 66580
rect 19050 66520 19110 66580
rect 18250 66270 18320 66280
rect 18250 66210 18310 66270
rect 18310 66210 18320 66270
rect 18250 66160 18320 66170
rect 18250 66100 18310 66160
rect 18310 66100 18320 66160
rect 17610 66000 17670 66060
rect 19050 66000 19110 66060
rect 18250 64560 18320 64570
rect 18250 64500 18310 64560
rect 18310 64500 18320 64560
rect 18250 64450 18320 64460
rect 18250 64390 18310 64450
rect 18310 64390 18320 64450
rect 17610 64290 17670 64350
rect 19050 64290 19110 64350
rect 18250 62850 18320 62860
rect 18250 62790 18310 62850
rect 18310 62790 18320 62850
rect 18250 62740 18320 62750
rect 18250 62680 18310 62740
rect 18310 62680 18320 62740
rect 17610 62580 17670 62640
rect 19050 62580 19110 62640
rect 18250 61140 18320 61150
rect 18250 61080 18310 61140
rect 18310 61080 18320 61140
rect 18250 61030 18320 61040
rect 18250 60970 18310 61030
rect 18310 60970 18320 61030
rect 17610 60870 17670 60930
rect 19050 60870 19110 60930
rect 14180 59680 14240 59740
rect 17490 59680 17550 59740
rect 19170 59680 19230 59740
rect 3280 59430 3350 59440
rect 3280 59370 3340 59430
rect 3340 59370 3350 59430
rect 3280 59320 3350 59330
rect 3280 59260 3340 59320
rect 3340 59260 3350 59320
rect 8270 59430 8340 59440
rect 8270 59370 8330 59430
rect 8330 59370 8340 59430
rect 8270 59320 8340 59330
rect 8270 59260 8330 59320
rect 8330 59260 8340 59320
rect 13260 59430 13330 59440
rect 13260 59370 13320 59430
rect 13320 59370 13330 59430
rect 13260 59320 13330 59330
rect 13260 59260 13320 59320
rect 13320 59260 13330 59320
rect 18250 59430 18320 59440
rect 18250 59370 18310 59430
rect 18310 59370 18320 59430
rect 18250 59320 18320 59330
rect 18250 59260 18310 59320
rect 18310 59260 18320 59320
rect 2640 59160 2700 59220
rect 4080 59160 4140 59220
rect 7630 59160 7690 59220
rect 9070 59160 9130 59220
rect 12500 59160 12560 59220
rect 14180 59160 14240 59220
rect 17490 59160 17550 59220
rect 19170 59160 19230 59220
rect 22600 66520 22660 66580
rect 24040 66520 24100 66580
rect 23240 66270 23310 66280
rect 23240 66210 23300 66270
rect 23300 66210 23310 66270
rect 23240 66160 23310 66170
rect 23240 66100 23300 66160
rect 23300 66100 23310 66160
rect 22600 66000 22660 66060
rect 24040 66000 24100 66060
rect 23240 64560 23310 64570
rect 23240 64500 23300 64560
rect 23300 64500 23310 64560
rect 23240 64450 23310 64460
rect 23240 64390 23300 64450
rect 23300 64390 23310 64450
rect 22600 64290 22660 64350
rect 24040 64290 24100 64350
rect 22480 63100 22540 63160
rect 24160 63100 24220 63160
rect 23240 62850 23310 62860
rect 23240 62790 23300 62850
rect 23300 62790 23310 62850
rect 23240 62740 23310 62750
rect 23240 62680 23300 62740
rect 23300 62680 23310 62740
rect 22480 62580 22540 62640
rect 24160 62580 24220 62640
rect 23240 61140 23310 61150
rect 23240 61080 23300 61140
rect 23300 61080 23310 61140
rect 23240 61030 23310 61040
rect 23240 60970 23300 61030
rect 23300 60970 23310 61030
rect 22480 60860 22540 60920
rect 24160 60860 24220 60920
rect 22360 59680 22420 59740
rect 24280 59680 24340 59740
rect 23240 59430 23310 59440
rect 23240 59370 23300 59430
rect 23300 59370 23310 59430
rect 23240 59320 23310 59330
rect 23240 59260 23300 59320
rect 23300 59260 23310 59320
rect 22360 59160 22420 59220
rect 24280 59160 24340 59220
rect 22240 57970 22300 58030
rect 27590 66520 27650 66580
rect 29030 66520 29090 66580
rect 28230 66270 28300 66280
rect 28230 66210 28290 66270
rect 28290 66210 28300 66270
rect 28230 66160 28300 66170
rect 28230 66100 28290 66160
rect 28290 66100 28300 66160
rect 27590 66000 27650 66060
rect 29030 66000 29090 66060
rect 28230 64560 28300 64570
rect 28230 64500 28290 64560
rect 28290 64500 28300 64560
rect 28230 64450 28300 64460
rect 28230 64390 28290 64450
rect 28290 64390 28300 64450
rect 27590 64290 27650 64350
rect 29030 64290 29090 64350
rect 27470 63100 27530 63160
rect 29150 63100 29210 63160
rect 28230 62850 28300 62860
rect 28230 62790 28290 62850
rect 28290 62790 28300 62850
rect 28230 62740 28300 62750
rect 28230 62680 28290 62740
rect 28290 62680 28300 62740
rect 27470 62580 27530 62640
rect 29150 62580 29210 62640
rect 28230 61140 28300 61150
rect 28230 61080 28290 61140
rect 28290 61080 28300 61140
rect 28230 61030 28300 61040
rect 28230 60970 28290 61030
rect 28290 60970 28300 61030
rect 27470 60860 27530 60920
rect 29150 60860 29210 60920
rect 27350 59680 27410 59740
rect 29270 59680 29330 59740
rect 28230 59430 28300 59440
rect 28230 59370 28290 59430
rect 28290 59370 28300 59430
rect 28230 59320 28300 59330
rect 28230 59260 28290 59320
rect 28290 59260 28300 59320
rect 27350 59160 27410 59220
rect 29270 59160 29330 59220
rect 24400 57970 24460 58030
rect 27230 57970 27290 58030
rect 29390 57970 29450 58030
rect 3280 57720 3350 57730
rect 3280 57660 3340 57720
rect 3340 57660 3350 57720
rect 3280 57610 3350 57620
rect 3280 57550 3340 57610
rect 3340 57550 3350 57610
rect 8270 57720 8340 57730
rect 8270 57660 8330 57720
rect 8330 57660 8340 57720
rect 8270 57610 8340 57620
rect 8270 57550 8330 57610
rect 8330 57550 8340 57610
rect 13260 57720 13330 57730
rect 13260 57660 13320 57720
rect 13320 57660 13330 57720
rect 13260 57610 13330 57620
rect 13260 57550 13320 57610
rect 13320 57550 13330 57610
rect 18250 57720 18320 57730
rect 18250 57660 18310 57720
rect 18310 57660 18320 57720
rect 18250 57610 18320 57620
rect 18250 57550 18310 57610
rect 18310 57550 18320 57610
rect 23240 57720 23310 57730
rect 23240 57660 23300 57720
rect 23300 57660 23310 57720
rect 23240 57610 23310 57620
rect 23240 57550 23300 57610
rect 23300 57550 23310 57610
rect 28230 57720 28300 57730
rect 28230 57660 28290 57720
rect 28290 57660 28300 57720
rect 28230 57610 28300 57620
rect 28230 57550 28290 57610
rect 28290 57550 28300 57610
rect 2640 57450 2700 57510
rect 4080 57450 4140 57510
rect 7630 57450 7690 57510
rect 9070 57450 9130 57510
rect 12500 57450 12560 57510
rect 14180 57450 14240 57510
rect 17490 57450 17550 57510
rect 19170 57450 19230 57510
rect 22240 57450 22300 57510
rect 24400 57450 24460 57510
rect 27230 57450 27290 57510
rect 29390 57450 29450 57510
rect 3280 56010 3350 56020
rect 3280 55950 3340 56010
rect 3340 55950 3350 56010
rect 3280 55900 3350 55910
rect 3280 55840 3340 55900
rect 3340 55840 3350 55900
rect 8270 56010 8340 56020
rect 8270 55950 8330 56010
rect 8330 55950 8340 56010
rect 8270 55900 8340 55910
rect 8270 55840 8330 55900
rect 8330 55840 8340 55900
rect 13260 56010 13330 56020
rect 13260 55950 13320 56010
rect 13320 55950 13330 56010
rect 13260 55900 13330 55910
rect 13260 55840 13320 55900
rect 13320 55840 13330 55900
rect 18250 56010 18320 56020
rect 18250 55950 18310 56010
rect 18310 55950 18320 56010
rect 18250 55900 18320 55910
rect 18250 55840 18310 55900
rect 18310 55840 18320 55900
rect 23240 56010 23310 56020
rect 23240 55950 23300 56010
rect 23300 55950 23310 56010
rect 23240 55900 23310 55910
rect 23240 55840 23300 55900
rect 23300 55840 23310 55900
rect 28230 56010 28300 56020
rect 28230 55950 28290 56010
rect 28290 55950 28300 56010
rect 28230 55900 28300 55910
rect 28230 55840 28290 55900
rect 28290 55840 28300 55900
rect 2640 55740 2700 55800
rect 4080 55740 4140 55800
rect 7630 55740 7690 55800
rect 9070 55740 9130 55800
rect 12500 55740 12560 55800
rect 14180 55740 14240 55800
rect 17490 55740 17550 55800
rect 19170 55740 19230 55800
rect 22240 55740 22300 55800
rect 24400 55740 24460 55800
rect 27230 55740 27290 55800
rect 29390 55740 29450 55800
rect 32580 66520 32640 66580
rect 34020 66520 34080 66580
rect 33220 66270 33290 66280
rect 33220 66210 33280 66270
rect 33280 66210 33290 66270
rect 33220 66160 33290 66170
rect 33220 66100 33280 66160
rect 33280 66100 33290 66160
rect 32580 66000 32640 66060
rect 34020 66000 34080 66060
rect 33220 64560 33290 64570
rect 33220 64500 33280 64560
rect 33280 64500 33290 64560
rect 33220 64450 33290 64460
rect 33220 64390 33280 64450
rect 33280 64390 33290 64450
rect 32580 64290 32640 64350
rect 34020 64290 34080 64350
rect 32460 63100 32520 63160
rect 34140 63100 34200 63160
rect 33220 62850 33290 62860
rect 33220 62790 33280 62850
rect 33280 62790 33290 62850
rect 33220 62740 33290 62750
rect 33220 62680 33280 62740
rect 33280 62680 33290 62740
rect 32460 62580 32520 62640
rect 34140 62580 34200 62640
rect 33220 61140 33290 61150
rect 33220 61080 33280 61140
rect 33280 61080 33290 61140
rect 33220 61030 33290 61040
rect 33220 60970 33280 61030
rect 33280 60970 33290 61030
rect 32460 60870 32520 60930
rect 34140 60870 34200 60930
rect 32340 59680 32400 59740
rect 34260 59680 34320 59740
rect 33220 59430 33290 59440
rect 33220 59370 33280 59430
rect 33280 59370 33290 59430
rect 33220 59320 33290 59330
rect 33220 59260 33280 59320
rect 33280 59260 33290 59320
rect 32340 59160 32400 59220
rect 34260 59160 34320 59220
rect 32220 57970 32280 58030
rect 34380 57970 34440 58030
rect 33220 57720 33290 57730
rect 33220 57660 33280 57720
rect 33280 57660 33290 57720
rect 33220 57610 33290 57620
rect 33220 57550 33280 57610
rect 33280 57550 33290 57610
rect 32220 57450 32280 57510
rect 34380 57450 34440 57510
rect 32100 56260 32160 56320
rect 34500 56260 34560 56320
rect 33220 56010 33290 56020
rect 33220 55950 33280 56010
rect 33280 55950 33290 56010
rect 33220 55900 33290 55910
rect 33220 55840 33280 55900
rect 33280 55840 33290 55900
rect 32100 55740 32160 55800
rect 34500 55740 34560 55800
rect 31980 54550 32040 54610
rect 34620 54550 34680 54610
rect 37570 66530 37630 66590
rect 39010 66530 39070 66590
rect 38210 66270 38280 66280
rect 38210 66210 38270 66270
rect 38270 66210 38280 66270
rect 38210 66160 38280 66170
rect 38210 66100 38270 66160
rect 38270 66100 38280 66160
rect 37570 66010 37630 66070
rect 39010 66010 39070 66070
rect 38210 64560 38280 64570
rect 38210 64500 38270 64560
rect 38270 64500 38280 64560
rect 38210 64450 38280 64460
rect 38210 64390 38270 64450
rect 38270 64390 38280 64450
rect 37570 64300 37630 64360
rect 39010 64300 39070 64360
rect 37450 63110 37510 63170
rect 39130 63110 39190 63170
rect 38210 62850 38280 62860
rect 38210 62790 38270 62850
rect 38270 62790 38280 62850
rect 38210 62740 38280 62750
rect 38210 62680 38270 62740
rect 38270 62680 38280 62740
rect 37450 62590 37510 62650
rect 39130 62590 39190 62650
rect 38210 61140 38280 61150
rect 38210 61080 38270 61140
rect 38270 61080 38280 61140
rect 38210 61030 38280 61040
rect 38210 60970 38270 61030
rect 38270 60970 38280 61030
rect 37450 60880 37510 60940
rect 39130 60880 39190 60940
rect 37330 59690 37390 59750
rect 39250 59690 39310 59750
rect 38210 59430 38280 59440
rect 38210 59370 38270 59430
rect 38270 59370 38280 59430
rect 38210 59320 38280 59330
rect 38210 59260 38270 59320
rect 38270 59260 38280 59320
rect 37330 59170 37390 59230
rect 39250 59170 39310 59230
rect 37210 57980 37270 58040
rect 39370 57980 39430 58040
rect 38210 57720 38280 57730
rect 38210 57660 38270 57720
rect 38270 57660 38280 57720
rect 38210 57610 38280 57620
rect 38210 57550 38270 57610
rect 38270 57550 38280 57610
rect 37210 57460 37270 57520
rect 39370 57460 39430 57520
rect 37090 56270 37150 56330
rect 39490 56270 39550 56330
rect 38210 56010 38280 56020
rect 38210 55950 38270 56010
rect 38270 55950 38280 56010
rect 38210 55900 38280 55910
rect 38210 55840 38270 55900
rect 38270 55840 38280 55900
rect 37090 55750 37150 55810
rect 39490 55750 39550 55810
rect 36970 54550 37030 54610
rect 39610 54600 39670 54660
rect 3280 54300 3350 54310
rect 3280 54240 3340 54300
rect 3340 54240 3350 54300
rect 3280 54190 3350 54200
rect 3280 54130 3340 54190
rect 3340 54130 3350 54190
rect 8270 54300 8340 54310
rect 8270 54240 8330 54300
rect 8330 54240 8340 54300
rect 8270 54190 8340 54200
rect 8270 54130 8330 54190
rect 8330 54130 8340 54190
rect 13260 54300 13330 54310
rect 13260 54240 13320 54300
rect 13320 54240 13330 54300
rect 13260 54190 13330 54200
rect 13260 54130 13320 54190
rect 13320 54130 13330 54190
rect 18250 54300 18320 54310
rect 18250 54240 18310 54300
rect 18310 54240 18320 54300
rect 18250 54190 18320 54200
rect 18250 54130 18310 54190
rect 18310 54130 18320 54190
rect 23240 54300 23310 54310
rect 23240 54240 23300 54300
rect 23300 54240 23310 54300
rect 23240 54190 23310 54200
rect 23240 54130 23300 54190
rect 23300 54130 23310 54190
rect 28230 54300 28300 54310
rect 28230 54240 28290 54300
rect 28290 54240 28300 54300
rect 28230 54190 28300 54200
rect 28230 54130 28290 54190
rect 28290 54130 28300 54190
rect 33220 54300 33290 54310
rect 33220 54240 33280 54300
rect 33280 54240 33290 54300
rect 42560 66530 42620 66590
rect 44000 66530 44060 66590
rect 43200 66270 43270 66280
rect 43200 66210 43260 66270
rect 43260 66210 43270 66270
rect 43200 66160 43270 66170
rect 43200 66100 43260 66160
rect 43260 66100 43270 66160
rect 42560 66010 42620 66070
rect 44000 66010 44060 66070
rect 43200 64560 43270 64570
rect 43200 64500 43260 64560
rect 43260 64500 43270 64560
rect 43200 64450 43270 64460
rect 43200 64390 43260 64450
rect 43260 64390 43270 64450
rect 42560 64300 42620 64360
rect 44000 64300 44060 64360
rect 42440 63110 42500 63170
rect 44120 63110 44180 63170
rect 43200 62850 43270 62860
rect 43200 62790 43260 62850
rect 43260 62790 43270 62850
rect 43200 62740 43270 62750
rect 43200 62680 43260 62740
rect 43260 62680 43270 62740
rect 42440 62590 42500 62650
rect 44120 62590 44180 62650
rect 43200 61140 43270 61150
rect 43200 61080 43260 61140
rect 43260 61080 43270 61140
rect 43200 61030 43270 61040
rect 43200 60970 43260 61030
rect 43260 60970 43270 61030
rect 42440 60880 42500 60940
rect 44120 60880 44180 60940
rect 42320 59690 42380 59750
rect 44240 59690 44300 59750
rect 43200 59430 43270 59440
rect 43200 59370 43260 59430
rect 43260 59370 43270 59430
rect 43200 59320 43270 59330
rect 43200 59260 43260 59320
rect 43260 59260 43270 59320
rect 42320 59170 42380 59230
rect 44240 59170 44300 59230
rect 42200 57980 42260 58040
rect 44360 57980 44420 58040
rect 43200 57720 43270 57730
rect 43200 57660 43260 57720
rect 43260 57660 43270 57720
rect 43200 57610 43270 57620
rect 43200 57550 43260 57610
rect 43260 57550 43270 57610
rect 42200 57460 42260 57520
rect 44360 57460 44420 57520
rect 42080 56270 42140 56330
rect 44480 56270 44540 56330
rect 43200 56010 43270 56020
rect 43200 55950 43260 56010
rect 43260 55950 43270 56010
rect 43200 55900 43270 55910
rect 43200 55840 43260 55900
rect 43260 55840 43270 55900
rect 42080 55750 42140 55810
rect 44480 55750 44540 55810
rect 41960 54550 42020 54610
rect 44600 54600 44660 54660
rect 33220 54190 33290 54200
rect 33220 54130 33280 54190
rect 33280 54130 33290 54190
rect 2640 54030 2700 54090
rect 4080 54030 4140 54090
rect 7630 54030 7690 54090
rect 9070 54030 9130 54090
rect 12500 54030 12560 54090
rect 14180 54030 14240 54090
rect 17490 54030 17550 54090
rect 19170 54030 19230 54090
rect 22240 54030 22300 54090
rect 24400 54030 24460 54090
rect 27230 54030 27290 54090
rect 29390 54030 29450 54090
rect 31980 54030 32040 54090
rect 34620 54030 34680 54090
rect 38210 54300 38280 54310
rect 38210 54240 38270 54300
rect 38270 54240 38280 54300
rect 38210 54190 38280 54200
rect 38210 54130 38270 54190
rect 38270 54130 38280 54190
rect 47550 66520 47610 66580
rect 48990 66520 49050 66580
rect 48190 66270 48260 66280
rect 48190 66210 48250 66270
rect 48250 66210 48260 66270
rect 48190 66160 48260 66170
rect 48190 66100 48250 66160
rect 48250 66100 48260 66160
rect 47550 66000 47610 66060
rect 48990 66000 49050 66060
rect 48190 64560 48260 64570
rect 48190 64500 48250 64560
rect 48250 64500 48260 64560
rect 48190 64450 48260 64460
rect 48190 64390 48250 64450
rect 48250 64390 48260 64450
rect 47550 64290 47610 64350
rect 48990 64290 49050 64350
rect 47430 63100 47490 63160
rect 49110 63100 49170 63160
rect 48190 62850 48260 62860
rect 48190 62790 48250 62850
rect 48250 62790 48260 62850
rect 48190 62740 48260 62750
rect 48190 62680 48250 62740
rect 48250 62680 48260 62740
rect 47430 62580 47490 62640
rect 49110 62580 49170 62640
rect 48190 61140 48260 61150
rect 48190 61080 48250 61140
rect 48250 61080 48260 61140
rect 48190 61030 48260 61040
rect 48190 60970 48250 61030
rect 48250 60970 48260 61030
rect 47430 60870 47490 60930
rect 49110 60870 49170 60930
rect 47310 59680 47370 59740
rect 49230 59680 49290 59740
rect 48190 59430 48260 59440
rect 48190 59370 48250 59430
rect 48250 59370 48260 59430
rect 48190 59320 48260 59330
rect 48190 59260 48250 59320
rect 48250 59260 48260 59320
rect 47310 59160 47370 59220
rect 49230 59160 49290 59220
rect 47190 57970 47250 58030
rect 49350 57970 49410 58030
rect 48190 57720 48260 57730
rect 48190 57660 48250 57720
rect 48250 57660 48260 57720
rect 48190 57610 48260 57620
rect 48190 57550 48250 57610
rect 48250 57550 48260 57610
rect 47190 57450 47250 57510
rect 49350 57450 49410 57510
rect 47070 56260 47130 56320
rect 49470 56260 49530 56320
rect 48190 56010 48260 56020
rect 48190 55950 48250 56010
rect 48250 55950 48260 56010
rect 48190 55900 48260 55910
rect 48190 55840 48250 55900
rect 48250 55840 48260 55900
rect 47070 55740 47130 55800
rect 49470 55740 49530 55800
rect 46950 54550 47010 54610
rect 52540 66520 52600 66580
rect 53980 66520 54040 66580
rect 53180 66270 53250 66280
rect 53180 66210 53240 66270
rect 53240 66210 53250 66270
rect 53180 66160 53250 66170
rect 53180 66100 53240 66160
rect 53240 66100 53250 66160
rect 52540 66000 52600 66060
rect 53980 66000 54040 66060
rect 53180 64560 53250 64570
rect 53180 64500 53240 64560
rect 53240 64500 53250 64560
rect 53180 64450 53250 64460
rect 53180 64390 53240 64450
rect 53240 64390 53250 64450
rect 52540 64290 52600 64350
rect 53980 64290 54040 64350
rect 52420 63100 52480 63160
rect 54100 63100 54160 63160
rect 53180 62850 53250 62860
rect 53180 62790 53240 62850
rect 53240 62790 53250 62850
rect 53180 62740 53250 62750
rect 53180 62680 53240 62740
rect 53240 62680 53250 62740
rect 52420 62580 52480 62640
rect 54100 62580 54160 62640
rect 53180 61140 53250 61150
rect 53180 61080 53240 61140
rect 53240 61080 53250 61140
rect 53180 61030 53250 61040
rect 53180 60970 53240 61030
rect 53240 60970 53250 61030
rect 52420 60860 52480 60920
rect 54100 60860 54160 60920
rect 52300 59680 52360 59740
rect 54220 59680 54280 59740
rect 53180 59430 53250 59440
rect 53180 59370 53240 59430
rect 53240 59370 53250 59430
rect 53180 59320 53250 59330
rect 53180 59260 53240 59320
rect 53240 59260 53250 59320
rect 52300 59160 52360 59220
rect 54220 59160 54280 59220
rect 52180 57970 52240 58030
rect 57530 66520 57590 66580
rect 58970 66520 59030 66580
rect 58170 66270 58240 66280
rect 58170 66210 58230 66270
rect 58230 66210 58240 66270
rect 58170 66160 58240 66170
rect 58170 66100 58230 66160
rect 58230 66100 58240 66160
rect 57530 66000 57590 66060
rect 58970 66000 59030 66060
rect 58170 64560 58240 64570
rect 58170 64500 58230 64560
rect 58230 64500 58240 64560
rect 58170 64450 58240 64460
rect 58170 64390 58230 64450
rect 58230 64390 58240 64450
rect 57530 64290 57590 64350
rect 58970 64290 59030 64350
rect 57410 63100 57470 63160
rect 59090 63100 59150 63160
rect 58170 62850 58240 62860
rect 58170 62790 58230 62850
rect 58230 62790 58240 62850
rect 58170 62740 58240 62750
rect 58170 62680 58230 62740
rect 58230 62680 58240 62740
rect 57410 62580 57470 62640
rect 59090 62580 59150 62640
rect 58170 61140 58240 61150
rect 58170 61080 58230 61140
rect 58230 61080 58240 61140
rect 58170 61030 58240 61040
rect 58170 60970 58230 61030
rect 58230 60970 58240 61030
rect 57410 60860 57470 60920
rect 59090 60860 59150 60920
rect 57290 59680 57350 59740
rect 59210 59680 59270 59740
rect 58170 59430 58240 59440
rect 58170 59370 58230 59430
rect 58230 59370 58240 59430
rect 58170 59320 58240 59330
rect 58170 59260 58230 59320
rect 58230 59260 58240 59320
rect 57290 59160 57350 59220
rect 59210 59160 59270 59220
rect 54340 57970 54400 58030
rect 57170 57970 57230 58030
rect 62520 66520 62580 66580
rect 63960 66520 64020 66580
rect 63160 66270 63230 66280
rect 63160 66210 63220 66270
rect 63220 66210 63230 66270
rect 63160 66160 63230 66170
rect 63160 66100 63220 66160
rect 63220 66100 63230 66160
rect 62520 66000 62580 66060
rect 63960 66000 64020 66060
rect 63160 64560 63230 64570
rect 63160 64500 63220 64560
rect 63220 64500 63230 64560
rect 63160 64450 63230 64460
rect 63160 64390 63220 64450
rect 63220 64390 63230 64450
rect 62520 64290 62580 64350
rect 63960 64290 64020 64350
rect 63160 62850 63230 62860
rect 63160 62790 63220 62850
rect 63220 62790 63230 62850
rect 63160 62740 63230 62750
rect 63160 62680 63220 62740
rect 63220 62680 63230 62740
rect 62520 62580 62580 62640
rect 63960 62580 64020 62640
rect 63160 61140 63230 61150
rect 63160 61080 63220 61140
rect 63220 61080 63230 61140
rect 63160 61030 63230 61040
rect 63160 60970 63220 61030
rect 63220 60970 63230 61030
rect 62520 60870 62580 60930
rect 63960 60870 64020 60930
rect 62400 59680 62460 59740
rect 67510 66520 67570 66580
rect 68950 66520 69010 66580
rect 68150 66270 68220 66280
rect 68150 66210 68210 66270
rect 68210 66210 68220 66270
rect 68150 66160 68220 66170
rect 68150 66100 68210 66160
rect 68210 66100 68220 66160
rect 67510 66000 67570 66060
rect 68950 66000 69010 66060
rect 68150 64560 68220 64570
rect 68150 64500 68210 64560
rect 68210 64500 68220 64560
rect 68150 64450 68220 64460
rect 68150 64390 68210 64450
rect 68210 64390 68220 64450
rect 67510 64290 67570 64350
rect 68950 64290 69010 64350
rect 68150 62850 68220 62860
rect 68150 62790 68210 62850
rect 68210 62790 68220 62850
rect 68150 62740 68220 62750
rect 68150 62680 68210 62740
rect 68210 62680 68220 62740
rect 67510 62580 67570 62640
rect 68950 62580 69010 62640
rect 68150 61140 68220 61150
rect 68150 61080 68210 61140
rect 68210 61080 68220 61140
rect 68150 61030 68220 61040
rect 68150 60970 68210 61030
rect 68210 60970 68220 61030
rect 67510 60870 67570 60930
rect 68950 60870 69010 60930
rect 64080 59680 64140 59740
rect 67390 59680 67450 59740
rect 72500 66520 72560 66580
rect 73940 66520 74000 66580
rect 77490 66520 77550 66580
rect 78930 66520 78990 66580
rect 73140 66270 73210 66280
rect 73140 66210 73200 66270
rect 73200 66210 73210 66270
rect 73140 66160 73210 66170
rect 73140 66100 73200 66160
rect 73200 66100 73210 66160
rect 78130 66270 78200 66280
rect 78130 66210 78190 66270
rect 78190 66210 78200 66270
rect 78130 66160 78200 66170
rect 78130 66100 78190 66160
rect 78190 66100 78200 66160
rect 72500 66000 72560 66060
rect 73940 66000 74000 66060
rect 77490 66000 77550 66060
rect 78930 66000 78990 66060
rect 73140 64560 73210 64570
rect 73140 64500 73200 64560
rect 73200 64500 73210 64560
rect 73140 64450 73210 64460
rect 73140 64390 73200 64450
rect 73200 64390 73210 64450
rect 78130 64560 78200 64570
rect 78130 64500 78190 64560
rect 78190 64500 78200 64560
rect 78130 64450 78200 64460
rect 78130 64390 78190 64450
rect 78190 64390 78200 64450
rect 72500 64290 72560 64350
rect 73940 64290 74000 64350
rect 77490 64290 77550 64350
rect 78930 64290 78990 64350
rect 73140 62850 73210 62860
rect 73140 62790 73200 62850
rect 73200 62790 73210 62850
rect 73140 62740 73210 62750
rect 73140 62680 73200 62740
rect 73200 62680 73210 62740
rect 78130 62850 78200 62860
rect 78130 62790 78190 62850
rect 78190 62790 78200 62850
rect 78130 62740 78200 62750
rect 78130 62680 78190 62740
rect 78190 62680 78200 62740
rect 72500 62580 72560 62640
rect 73940 62580 74000 62640
rect 77490 62580 77550 62640
rect 78930 62580 78990 62640
rect 73140 61140 73210 61150
rect 73140 61080 73200 61140
rect 73200 61080 73210 61140
rect 73140 61030 73210 61040
rect 73140 60970 73200 61030
rect 73200 60970 73210 61030
rect 78130 61140 78200 61150
rect 78130 61080 78190 61140
rect 78190 61080 78200 61140
rect 78130 61030 78200 61040
rect 78130 60970 78190 61030
rect 78190 60970 78200 61030
rect 72500 60870 72560 60930
rect 73940 60870 74000 60930
rect 77490 60870 77550 60930
rect 78930 60870 78990 60930
rect 69070 59680 69130 59740
rect 63160 59430 63230 59440
rect 63160 59370 63220 59430
rect 63220 59370 63230 59430
rect 63160 59320 63230 59330
rect 63160 59260 63220 59320
rect 63220 59260 63230 59320
rect 68150 59430 68220 59440
rect 68150 59370 68210 59430
rect 68210 59370 68220 59430
rect 68150 59320 68220 59330
rect 68150 59260 68210 59320
rect 68210 59260 68220 59320
rect 73140 59430 73210 59440
rect 73140 59370 73200 59430
rect 73200 59370 73210 59430
rect 73140 59320 73210 59330
rect 73140 59260 73200 59320
rect 73200 59260 73210 59320
rect 78130 59430 78200 59440
rect 78130 59370 78190 59430
rect 78190 59370 78200 59430
rect 78130 59320 78200 59330
rect 78130 59260 78190 59320
rect 78190 59260 78200 59320
rect 62400 59160 62460 59220
rect 64080 59160 64140 59220
rect 67390 59160 67450 59220
rect 69070 59160 69130 59220
rect 72500 59160 72560 59220
rect 73940 59160 74000 59220
rect 77490 59160 77550 59220
rect 78930 59160 78990 59220
rect 59330 57970 59390 58030
rect 53180 57720 53250 57730
rect 53180 57660 53240 57720
rect 53240 57660 53250 57720
rect 53180 57610 53250 57620
rect 53180 57550 53240 57610
rect 53240 57550 53250 57610
rect 58170 57720 58240 57730
rect 58170 57660 58230 57720
rect 58230 57660 58240 57720
rect 58170 57610 58240 57620
rect 58170 57550 58230 57610
rect 58230 57550 58240 57610
rect 63160 57720 63230 57730
rect 63160 57660 63220 57720
rect 63220 57660 63230 57720
rect 63160 57610 63230 57620
rect 63160 57550 63220 57610
rect 63220 57550 63230 57610
rect 68150 57720 68220 57730
rect 68150 57660 68210 57720
rect 68210 57660 68220 57720
rect 68150 57610 68220 57620
rect 68150 57550 68210 57610
rect 68210 57550 68220 57610
rect 73140 57720 73210 57730
rect 73140 57660 73200 57720
rect 73200 57660 73210 57720
rect 73140 57610 73210 57620
rect 73140 57550 73200 57610
rect 73200 57550 73210 57610
rect 78130 57720 78200 57730
rect 78130 57660 78190 57720
rect 78190 57660 78200 57720
rect 78130 57610 78200 57620
rect 78130 57550 78190 57610
rect 78190 57550 78200 57610
rect 52180 57450 52240 57510
rect 54340 57450 54400 57510
rect 57170 57450 57230 57510
rect 59330 57450 59390 57510
rect 62400 57450 62460 57510
rect 64080 57450 64140 57510
rect 67390 57450 67450 57510
rect 69070 57450 69130 57510
rect 72500 57450 72560 57510
rect 73940 57450 74000 57510
rect 77490 57450 77550 57510
rect 78930 57450 78990 57510
rect 53180 56010 53250 56020
rect 53180 55950 53240 56010
rect 53240 55950 53250 56010
rect 53180 55900 53250 55910
rect 53180 55840 53240 55900
rect 53240 55840 53250 55900
rect 58170 56010 58240 56020
rect 58170 55950 58230 56010
rect 58230 55950 58240 56010
rect 58170 55900 58240 55910
rect 58170 55840 58230 55900
rect 58230 55840 58240 55900
rect 63160 56010 63230 56020
rect 63160 55950 63220 56010
rect 63220 55950 63230 56010
rect 63160 55900 63230 55910
rect 63160 55840 63220 55900
rect 63220 55840 63230 55900
rect 68150 56010 68220 56020
rect 68150 55950 68210 56010
rect 68210 55950 68220 56010
rect 68150 55900 68220 55910
rect 68150 55840 68210 55900
rect 68210 55840 68220 55900
rect 73140 56010 73210 56020
rect 73140 55950 73200 56010
rect 73200 55950 73210 56010
rect 73140 55900 73210 55910
rect 73140 55840 73200 55900
rect 73200 55840 73210 55900
rect 78130 56010 78200 56020
rect 78130 55950 78190 56010
rect 78190 55950 78200 56010
rect 78130 55900 78200 55910
rect 78130 55840 78190 55900
rect 78190 55840 78200 55900
rect 52180 55740 52240 55800
rect 54340 55740 54400 55800
rect 57170 55740 57230 55800
rect 59330 55740 59390 55800
rect 62400 55740 62460 55800
rect 64080 55740 64140 55800
rect 67390 55740 67450 55800
rect 69070 55740 69130 55800
rect 72500 55740 72560 55800
rect 73940 55740 74000 55800
rect 77490 55740 77550 55800
rect 78930 55740 78990 55800
rect 49590 54550 49650 54610
rect 3280 52590 3350 52600
rect 3280 52530 3340 52590
rect 3340 52530 3350 52590
rect 3280 52480 3350 52490
rect 3280 52420 3340 52480
rect 3340 52420 3350 52480
rect 8270 52590 8340 52600
rect 8270 52530 8330 52590
rect 8330 52530 8340 52590
rect 8270 52480 8340 52490
rect 8270 52420 8330 52480
rect 8330 52420 8340 52480
rect 13260 52590 13330 52600
rect 13260 52530 13320 52590
rect 13320 52530 13330 52590
rect 13260 52480 13330 52490
rect 13260 52420 13320 52480
rect 13320 52420 13330 52480
rect 18250 52590 18320 52600
rect 18250 52530 18310 52590
rect 18310 52530 18320 52590
rect 18250 52480 18320 52490
rect 18250 52420 18310 52480
rect 18310 52420 18320 52480
rect 23240 52590 23310 52600
rect 23240 52530 23300 52590
rect 23300 52530 23310 52590
rect 23240 52480 23310 52490
rect 23240 52420 23300 52480
rect 23300 52420 23310 52480
rect 28230 52590 28300 52600
rect 28230 52530 28290 52590
rect 28290 52530 28300 52590
rect 28230 52480 28300 52490
rect 28230 52420 28290 52480
rect 28290 52420 28300 52480
rect 33220 52590 33290 52600
rect 33220 52530 33280 52590
rect 33280 52530 33290 52590
rect 33220 52480 33290 52490
rect 33220 52420 33280 52480
rect 33280 52420 33290 52480
rect 2640 52320 2700 52380
rect 4080 52320 4140 52380
rect 7630 52320 7690 52380
rect 9070 52320 9130 52380
rect 12500 52320 12560 52380
rect 14180 52320 14240 52380
rect 17490 52320 17550 52380
rect 19170 52320 19230 52380
rect 22240 52320 22300 52380
rect 24400 52320 24460 52380
rect 27230 52320 27290 52380
rect 29390 52320 29450 52380
rect 31980 52320 32040 52380
rect 34620 52320 34680 52380
rect 3280 50880 3350 50890
rect 3280 50820 3340 50880
rect 3340 50820 3350 50880
rect 3280 50770 3350 50780
rect 3280 50710 3340 50770
rect 3340 50710 3350 50770
rect 8270 50880 8340 50890
rect 8270 50820 8330 50880
rect 8330 50820 8340 50880
rect 8270 50770 8340 50780
rect 8270 50710 8330 50770
rect 8330 50710 8340 50770
rect 13260 50880 13330 50890
rect 13260 50820 13320 50880
rect 13320 50820 13330 50880
rect 13260 50770 13330 50780
rect 13260 50710 13320 50770
rect 13320 50710 13330 50770
rect 18250 50880 18320 50890
rect 18250 50820 18310 50880
rect 18310 50820 18320 50880
rect 18250 50770 18320 50780
rect 18250 50710 18310 50770
rect 18310 50710 18320 50770
rect 23240 50880 23310 50890
rect 23240 50820 23300 50880
rect 23300 50820 23310 50880
rect 23240 50770 23310 50780
rect 23240 50710 23300 50770
rect 23300 50710 23310 50770
rect 28230 50880 28300 50890
rect 28230 50820 28290 50880
rect 28290 50820 28300 50880
rect 28230 50770 28300 50780
rect 28230 50710 28290 50770
rect 28290 50710 28300 50770
rect 2640 50610 2700 50670
rect 4080 50610 4140 50670
rect 7630 50610 7690 50670
rect 9070 50610 9130 50670
rect 12500 50610 12560 50670
rect 14180 50610 14240 50670
rect 17490 50610 17550 50670
rect 19170 50610 19230 50670
rect 22240 50610 22300 50670
rect 24400 50610 24460 50670
rect 27230 50610 27290 50670
rect 29390 50610 29450 50670
rect 3280 49170 3350 49180
rect 3280 49110 3340 49170
rect 3340 49110 3350 49170
rect 3280 49060 3350 49070
rect 3280 49000 3340 49060
rect 3340 49000 3350 49060
rect 8270 49170 8340 49180
rect 8270 49110 8330 49170
rect 8330 49110 8340 49170
rect 8270 49060 8340 49070
rect 8270 49000 8330 49060
rect 8330 49000 8340 49060
rect 13260 49170 13330 49180
rect 13260 49110 13320 49170
rect 13320 49110 13330 49170
rect 13260 49060 13330 49070
rect 13260 49000 13320 49060
rect 13320 49000 13330 49060
rect 18250 49170 18320 49180
rect 18250 49110 18310 49170
rect 18310 49110 18320 49170
rect 18250 49060 18320 49070
rect 18250 49000 18310 49060
rect 18310 49000 18320 49060
rect 23240 49170 23310 49180
rect 23240 49110 23300 49170
rect 23300 49110 23310 49170
rect 23240 49060 23310 49070
rect 23240 49000 23300 49060
rect 23300 49000 23310 49060
rect 28230 49170 28300 49180
rect 28230 49110 28290 49170
rect 28290 49110 28300 49170
rect 28230 49060 28300 49070
rect 28230 49000 28290 49060
rect 28290 49000 28300 49060
rect 2640 48900 2700 48960
rect 4080 48900 4140 48960
rect 7630 48900 7690 48960
rect 9070 48900 9130 48960
rect 12500 48900 12560 48960
rect 14180 48900 14240 48960
rect 17490 48900 17550 48960
rect 19170 48900 19230 48960
rect 22240 48900 22300 48960
rect 24400 48900 24460 48960
rect 27230 48900 27290 48960
rect 29390 48900 29450 48960
rect 3280 47460 3350 47470
rect 3280 47400 3340 47460
rect 3340 47400 3350 47460
rect 3280 47350 3350 47360
rect 3280 47290 3340 47350
rect 3340 47290 3350 47350
rect 8270 47460 8340 47470
rect 8270 47400 8330 47460
rect 8330 47400 8340 47460
rect 8270 47350 8340 47360
rect 8270 47290 8330 47350
rect 8330 47290 8340 47350
rect 13260 47460 13330 47470
rect 13260 47400 13320 47460
rect 13320 47400 13330 47460
rect 13260 47350 13330 47360
rect 13260 47290 13320 47350
rect 13320 47290 13330 47350
rect 18250 47460 18320 47470
rect 18250 47400 18310 47460
rect 18310 47400 18320 47460
rect 18250 47350 18320 47360
rect 18250 47290 18310 47350
rect 18310 47290 18320 47350
rect 2640 47190 2700 47250
rect 4080 47190 4140 47250
rect 7630 47190 7690 47250
rect 9070 47190 9130 47250
rect 12500 47190 12560 47250
rect 14180 47190 14240 47250
rect 17490 47190 17550 47250
rect 19170 47190 19230 47250
rect 3280 45750 3350 45760
rect 3280 45690 3340 45750
rect 3340 45690 3350 45750
rect 3280 45640 3350 45650
rect 3280 45580 3340 45640
rect 3340 45580 3350 45640
rect 8270 45750 8340 45760
rect 8270 45690 8330 45750
rect 8330 45690 8340 45750
rect 8270 45640 8340 45650
rect 8270 45580 8330 45640
rect 8330 45580 8340 45640
rect 2640 45480 2700 45540
rect 4080 45480 4140 45540
rect 7630 45480 7690 45540
rect 9070 45480 9130 45540
rect 3280 44040 3350 44050
rect 3280 43980 3340 44040
rect 3340 43980 3350 44040
rect 3280 43930 3350 43940
rect 3280 43870 3340 43930
rect 3340 43870 3350 43930
rect 8270 44040 8340 44050
rect 8270 43980 8330 44040
rect 8330 43980 8340 44040
rect 8270 43930 8340 43940
rect 8270 43870 8330 43930
rect 8330 43870 8340 43930
rect 2640 43770 2700 43830
rect 4080 43770 4140 43830
rect 7630 43770 7690 43830
rect 9070 43770 9130 43830
rect 3280 42330 3350 42340
rect 3280 42270 3340 42330
rect 3340 42270 3350 42330
rect 3280 42220 3350 42230
rect 3280 42160 3340 42220
rect 3340 42160 3350 42220
rect 8270 42330 8340 42340
rect 8270 42270 8330 42330
rect 8330 42270 8340 42330
rect 8270 42220 8340 42230
rect 8270 42160 8330 42220
rect 8330 42160 8340 42220
rect 2640 42060 2700 42120
rect 4080 42060 4140 42120
rect 7630 42060 7690 42120
rect 9070 42060 9130 42120
rect 3280 40620 3350 40630
rect 3280 40560 3340 40620
rect 3340 40560 3350 40620
rect 3280 40510 3350 40520
rect 3280 40450 3340 40510
rect 3340 40450 3350 40510
rect 8270 40620 8340 40630
rect 8270 40560 8330 40620
rect 8330 40560 8340 40620
rect 8270 40510 8340 40520
rect 8270 40450 8330 40510
rect 8330 40450 8340 40510
rect 2640 40350 2700 40410
rect 4080 40350 4140 40410
rect 7630 40350 7690 40410
rect 9070 40350 9130 40410
rect 2750 38770 2810 38830
rect 3820 38630 3880 38690
rect 2520 36250 2580 36310
rect 2460 36110 2520 36170
rect 7740 38770 7800 38830
rect 13260 45750 13330 45760
rect 13260 45690 13320 45750
rect 13320 45690 13330 45750
rect 13260 45640 13330 45650
rect 13260 45580 13320 45640
rect 13320 45580 13330 45640
rect 12620 45480 12680 45540
rect 14060 45480 14120 45540
rect 13260 44040 13330 44050
rect 13260 43980 13320 44040
rect 13320 43980 13330 44040
rect 13260 43930 13330 43940
rect 13260 43870 13320 43930
rect 13320 43870 13330 43930
rect 12620 43770 12680 43830
rect 14060 43770 14120 43830
rect 13260 42330 13330 42340
rect 13260 42270 13320 42330
rect 13320 42270 13330 42330
rect 13260 42220 13330 42230
rect 13260 42160 13320 42220
rect 13320 42160 13330 42220
rect 12620 42060 12680 42120
rect 14060 42060 14120 42120
rect 13260 40620 13330 40630
rect 13260 40560 13320 40620
rect 13320 40560 13330 40620
rect 13260 40510 13330 40520
rect 13260 40450 13320 40510
rect 13320 40450 13330 40510
rect 12620 40350 12680 40410
rect 14060 40350 14120 40410
rect 8810 38630 8870 38690
rect 7510 36250 7570 36310
rect 12320 36530 12380 36590
rect 12260 36390 12320 36450
rect 7450 36110 7510 36170
rect 12730 38770 12790 38830
rect 18250 45750 18320 45760
rect 18250 45690 18310 45750
rect 18310 45690 18320 45750
rect 18250 45640 18320 45650
rect 18250 45580 18310 45640
rect 18310 45580 18320 45640
rect 17610 45480 17670 45540
rect 19050 45480 19110 45540
rect 18250 44040 18320 44050
rect 18250 43980 18310 44040
rect 18310 43980 18320 44040
rect 18250 43930 18320 43940
rect 18250 43870 18310 43930
rect 18310 43870 18320 43930
rect 17610 43770 17670 43830
rect 19050 43770 19110 43830
rect 18250 42330 18320 42340
rect 18250 42270 18310 42330
rect 18310 42270 18320 42330
rect 18250 42220 18320 42230
rect 18250 42160 18310 42220
rect 18310 42160 18320 42220
rect 17610 42060 17670 42120
rect 19050 42060 19110 42120
rect 18250 40620 18320 40630
rect 18250 40560 18310 40620
rect 18310 40560 18320 40620
rect 18250 40510 18320 40520
rect 18250 40450 18310 40510
rect 18310 40450 18320 40510
rect 17610 40350 17670 40410
rect 19050 40350 19110 40410
rect 13800 38630 13860 38690
rect 12500 36250 12560 36310
rect 17310 36530 17370 36590
rect 17250 36390 17310 36450
rect 12440 36110 12500 36170
rect 17720 38770 17780 38830
rect 23240 47460 23310 47470
rect 23240 47400 23300 47460
rect 23300 47400 23310 47460
rect 23240 47350 23310 47360
rect 23240 47290 23300 47350
rect 23300 47290 23310 47350
rect 22360 47190 22420 47250
rect 24280 47190 24340 47250
rect 18790 38630 18850 38690
rect 17490 36250 17550 36310
rect 23240 45750 23310 45760
rect 23240 45690 23300 45750
rect 23300 45690 23310 45750
rect 23240 45640 23310 45650
rect 23240 45580 23300 45640
rect 23300 45580 23310 45640
rect 22480 45480 22540 45540
rect 24160 45480 24220 45540
rect 23240 44040 23310 44050
rect 23240 43980 23300 44040
rect 23300 43980 23310 44040
rect 23240 43930 23310 43940
rect 23240 43870 23300 43930
rect 23300 43870 23310 43930
rect 22480 43770 22540 43830
rect 24160 43770 24220 43830
rect 23240 42330 23310 42340
rect 23240 42270 23300 42330
rect 23300 42270 23310 42330
rect 23240 42220 23310 42230
rect 23240 42160 23300 42220
rect 23300 42160 23310 42220
rect 22600 42060 22660 42120
rect 24040 42060 24100 42120
rect 23240 40620 23310 40630
rect 23240 40560 23300 40620
rect 23300 40560 23310 40620
rect 23240 40510 23310 40520
rect 23240 40450 23300 40510
rect 23300 40450 23310 40510
rect 22600 40350 22660 40410
rect 24040 40350 24100 40410
rect 22120 37090 22180 37150
rect 22060 36950 22120 37010
rect 21940 36810 22000 36870
rect 21880 36670 21940 36730
rect 22300 36530 22360 36590
rect 22240 36390 22300 36450
rect 17430 36110 17490 36170
rect 22710 38770 22770 38830
rect 28230 47460 28300 47470
rect 28230 47400 28290 47460
rect 28290 47400 28300 47460
rect 28230 47350 28300 47360
rect 28230 47290 28290 47350
rect 28290 47290 28300 47350
rect 27350 47190 27410 47250
rect 29270 47190 29330 47250
rect 23780 38630 23840 38690
rect 22480 36250 22540 36310
rect 28230 45750 28300 45760
rect 28230 45690 28290 45750
rect 28290 45690 28300 45750
rect 28230 45640 28300 45650
rect 28230 45580 28290 45640
rect 28290 45580 28300 45640
rect 27470 45480 27530 45540
rect 29150 45480 29210 45540
rect 28230 44040 28300 44050
rect 28230 43980 28290 44040
rect 28290 43980 28300 44040
rect 28230 43930 28300 43940
rect 28230 43870 28290 43930
rect 28290 43870 28300 43930
rect 27470 43770 27530 43830
rect 29150 43770 29210 43830
rect 28230 42330 28300 42340
rect 28230 42270 28290 42330
rect 28290 42270 28300 42330
rect 28230 42220 28300 42230
rect 28230 42160 28290 42220
rect 28290 42160 28300 42220
rect 27590 42060 27650 42120
rect 29030 42060 29090 42120
rect 28230 40620 28300 40630
rect 28230 40560 28290 40620
rect 28290 40560 28300 40620
rect 28230 40510 28300 40520
rect 28230 40450 28290 40510
rect 28290 40450 28300 40510
rect 27590 40350 27650 40410
rect 29030 40350 29090 40410
rect 27110 37090 27170 37150
rect 27050 36950 27110 37010
rect 26930 36810 26990 36870
rect 26870 36670 26930 36730
rect 27290 36530 27350 36590
rect 27230 36390 27290 36450
rect 22420 36110 22480 36170
rect 27700 38770 27760 38830
rect 33220 50880 33290 50890
rect 33220 50820 33280 50880
rect 33280 50820 33290 50880
rect 33220 50770 33290 50780
rect 33220 50710 33280 50770
rect 33280 50710 33290 50770
rect 32100 50610 32160 50670
rect 34500 50610 34560 50670
rect 28770 38630 28830 38690
rect 27470 36250 27530 36310
rect 33220 49170 33290 49180
rect 33220 49110 33280 49170
rect 33280 49110 33290 49170
rect 33220 49060 33290 49070
rect 33220 49000 33280 49060
rect 33280 49000 33290 49060
rect 32220 48900 32280 48960
rect 34380 48900 34440 48960
rect 33220 47460 33290 47470
rect 33220 47400 33280 47460
rect 33280 47400 33290 47460
rect 33220 47350 33290 47360
rect 33220 47290 33280 47350
rect 33280 47290 33290 47350
rect 32340 47190 32400 47250
rect 34260 47190 34320 47250
rect 31740 37650 31800 37710
rect 31680 37510 31740 37570
rect 31560 37370 31620 37430
rect 31500 37230 31560 37290
rect 33220 45750 33290 45760
rect 33220 45690 33280 45750
rect 33280 45690 33290 45750
rect 33220 45640 33290 45650
rect 33220 45580 33280 45640
rect 33280 45580 33290 45640
rect 32460 45480 32520 45540
rect 34140 45480 34200 45540
rect 33220 44040 33290 44050
rect 33220 43980 33280 44040
rect 33280 43980 33290 44040
rect 33220 43930 33290 43940
rect 33220 43870 33280 43930
rect 33280 43870 33290 43930
rect 32460 43770 32520 43830
rect 34140 43770 34200 43830
rect 31920 37090 31980 37150
rect 31860 36950 31920 37010
rect 33220 42330 33290 42340
rect 33220 42270 33280 42330
rect 33280 42270 33290 42330
rect 33220 42220 33290 42230
rect 33220 42160 33280 42220
rect 33280 42160 33290 42220
rect 32580 42060 32640 42120
rect 34020 42060 34080 42120
rect 33220 40620 33290 40630
rect 33220 40560 33280 40620
rect 33280 40560 33290 40620
rect 33220 40510 33290 40520
rect 33220 40450 33280 40510
rect 33280 40450 33290 40510
rect 32580 40350 32640 40410
rect 34020 40350 34080 40410
rect 32100 36810 32160 36870
rect 32040 36670 32100 36730
rect 32280 36530 32340 36590
rect 32220 36390 32280 36450
rect 27410 36110 27470 36170
rect 32690 38770 32750 38830
rect 38210 52590 38280 52600
rect 38210 52530 38270 52590
rect 38270 52530 38280 52590
rect 38210 52480 38280 52490
rect 38210 52420 38270 52480
rect 38270 52420 38280 52480
rect 36970 52330 37030 52390
rect 33760 38630 33820 38690
rect 32460 36250 32520 36310
rect 39610 52330 39670 52390
rect 38210 50880 38280 50890
rect 38210 50820 38270 50880
rect 38270 50820 38280 50880
rect 38210 50770 38280 50780
rect 38210 50710 38270 50770
rect 38270 50710 38280 50770
rect 37090 50620 37150 50680
rect 36370 38490 36430 38550
rect 36310 38350 36370 38410
rect 39490 50620 39550 50680
rect 38210 49170 38280 49180
rect 38210 49110 38270 49170
rect 38270 49110 38280 49170
rect 38210 49060 38280 49070
rect 38210 49000 38270 49060
rect 38270 49000 38280 49060
rect 37210 48910 37270 48970
rect 36550 37930 36610 37990
rect 36490 37790 36550 37850
rect 39370 48910 39430 48970
rect 38210 47460 38280 47470
rect 38210 47400 38270 47460
rect 38270 47400 38280 47460
rect 38210 47350 38280 47360
rect 38210 47290 38270 47350
rect 38270 47290 38280 47350
rect 37330 47200 37390 47260
rect 36730 37370 36790 37430
rect 36670 37230 36730 37290
rect 39250 47200 39310 47260
rect 38210 45750 38280 45760
rect 38210 45690 38270 45750
rect 38270 45690 38280 45750
rect 38210 45640 38280 45650
rect 38210 45580 38270 45640
rect 38270 45580 38280 45640
rect 37450 45490 37510 45550
rect 39130 45490 39190 45550
rect 38210 44040 38280 44050
rect 38210 43980 38270 44040
rect 38270 43980 38280 44040
rect 38210 43930 38280 43940
rect 38210 43870 38270 43930
rect 38270 43870 38280 43930
rect 37450 43780 37510 43840
rect 36910 37090 36970 37150
rect 36850 36950 36910 37010
rect 39130 43770 39190 43830
rect 38210 42330 38280 42340
rect 38210 42270 38270 42330
rect 38270 42270 38280 42330
rect 38210 42220 38280 42230
rect 38210 42160 38270 42220
rect 38270 42160 38280 42220
rect 37570 42070 37630 42130
rect 39010 42060 39070 42120
rect 38210 40620 38280 40630
rect 38210 40560 38270 40620
rect 38270 40560 38280 40620
rect 38210 40510 38280 40520
rect 38210 40450 38270 40510
rect 38270 40450 38280 40510
rect 37570 40360 37630 40420
rect 37090 36810 37150 36870
rect 37030 36670 37090 36730
rect 39010 40360 39070 40420
rect 39010 40150 39070 40210
rect 37270 36530 37330 36590
rect 37210 36390 37270 36450
rect 32400 36110 32460 36170
rect 37680 38770 37740 38830
rect 43200 54300 43270 54310
rect 43200 54240 43260 54300
rect 43260 54240 43270 54300
rect 43200 54190 43270 54200
rect 43200 54130 43260 54190
rect 43260 54130 43270 54190
rect 48190 54300 48260 54310
rect 48190 54240 48250 54300
rect 48250 54240 48260 54300
rect 48190 54190 48260 54200
rect 48190 54130 48250 54190
rect 48250 54130 48260 54190
rect 53180 54300 53250 54310
rect 53180 54240 53240 54300
rect 53240 54240 53250 54300
rect 53180 54190 53250 54200
rect 53180 54130 53240 54190
rect 53240 54130 53250 54190
rect 58170 54300 58240 54310
rect 58170 54240 58230 54300
rect 58230 54240 58240 54300
rect 58170 54190 58240 54200
rect 58170 54130 58230 54190
rect 58230 54130 58240 54190
rect 63160 54300 63230 54310
rect 63160 54240 63220 54300
rect 63220 54240 63230 54300
rect 63160 54190 63230 54200
rect 63160 54130 63220 54190
rect 63220 54130 63230 54190
rect 68150 54300 68220 54310
rect 68150 54240 68210 54300
rect 68210 54240 68220 54300
rect 68150 54190 68220 54200
rect 68150 54130 68210 54190
rect 68210 54130 68220 54190
rect 73140 54300 73210 54310
rect 73140 54240 73200 54300
rect 73200 54240 73210 54300
rect 73140 54190 73210 54200
rect 73140 54130 73200 54190
rect 73200 54130 73210 54190
rect 78130 54300 78200 54310
rect 78130 54240 78190 54300
rect 78190 54240 78200 54300
rect 78130 54190 78200 54200
rect 78130 54130 78190 54190
rect 78190 54130 78200 54190
rect 43200 52590 43270 52600
rect 43200 52530 43260 52590
rect 43260 52530 43270 52590
rect 43200 52480 43270 52490
rect 43200 52420 43260 52480
rect 43260 52420 43270 52480
rect 41960 52330 42020 52390
rect 38750 38630 38810 38690
rect 37450 36250 37510 36310
rect 44600 52330 44660 52390
rect 43200 50880 43270 50890
rect 43200 50820 43260 50880
rect 43260 50820 43270 50880
rect 43200 50770 43270 50780
rect 43200 50710 43260 50770
rect 43260 50710 43270 50770
rect 42080 50620 42140 50680
rect 44480 50620 44540 50680
rect 43200 49170 43270 49180
rect 43200 49110 43260 49170
rect 43260 49110 43270 49170
rect 43200 49060 43270 49070
rect 43200 49000 43260 49060
rect 43260 49000 43270 49060
rect 42200 48910 42260 48970
rect 41540 38210 41600 38270
rect 41450 38070 41510 38130
rect 41360 37930 41420 37990
rect 41300 37790 41360 37850
rect 44360 48910 44420 48970
rect 43200 47460 43270 47470
rect 43200 47400 43260 47460
rect 43260 47400 43270 47460
rect 43200 47350 43270 47360
rect 43200 47290 43260 47350
rect 43260 47290 43270 47350
rect 42320 47200 42380 47260
rect 41720 37370 41780 37430
rect 41660 37230 41720 37290
rect 44240 47200 44300 47260
rect 43200 45750 43270 45760
rect 43200 45690 43260 45750
rect 43260 45690 43270 45750
rect 43200 45640 43270 45650
rect 43200 45580 43260 45640
rect 43260 45580 43270 45640
rect 42440 45490 42500 45550
rect 44120 45490 44180 45550
rect 43200 44040 43270 44050
rect 43200 43980 43260 44040
rect 43260 43980 43270 44040
rect 43200 43930 43270 43940
rect 43200 43870 43260 43930
rect 43260 43870 43270 43930
rect 42440 43780 42500 43840
rect 41900 37090 41960 37150
rect 41840 36950 41900 37010
rect 44120 43770 44180 43830
rect 43200 42330 43270 42340
rect 43200 42270 43260 42330
rect 43260 42270 43270 42330
rect 43200 42220 43270 42230
rect 43200 42160 43260 42220
rect 43260 42160 43270 42220
rect 42560 42070 42620 42130
rect 44000 42060 44060 42120
rect 43200 40620 43270 40630
rect 43200 40560 43260 40620
rect 43260 40560 43270 40620
rect 43200 40510 43270 40520
rect 43200 40450 43260 40510
rect 43260 40450 43270 40510
rect 42560 40360 42620 40420
rect 42080 36810 42140 36870
rect 42020 36670 42080 36730
rect 44000 40360 44060 40420
rect 44000 40150 44060 40210
rect 42260 36530 42320 36590
rect 42200 36390 42260 36450
rect 37390 36110 37450 36170
rect 42670 38770 42730 38830
rect 46950 54030 47010 54090
rect 49590 54030 49650 54090
rect 52180 54030 52240 54090
rect 54340 54030 54400 54090
rect 57170 54030 57230 54090
rect 59330 54030 59390 54090
rect 62400 54030 62460 54090
rect 64080 54030 64140 54090
rect 67390 54030 67450 54090
rect 69070 54030 69130 54090
rect 72500 54030 72560 54090
rect 73940 54030 74000 54090
rect 77490 54030 77550 54090
rect 78930 54030 78990 54090
rect 48190 52590 48260 52600
rect 48190 52530 48250 52590
rect 48250 52530 48260 52590
rect 48190 52480 48260 52490
rect 48190 52420 48250 52480
rect 48250 52420 48260 52480
rect 53180 52590 53250 52600
rect 53180 52530 53240 52590
rect 53240 52530 53250 52590
rect 53180 52480 53250 52490
rect 53180 52420 53240 52480
rect 53240 52420 53250 52480
rect 58170 52590 58240 52600
rect 58170 52530 58230 52590
rect 58230 52530 58240 52590
rect 58170 52480 58240 52490
rect 58170 52420 58230 52480
rect 58230 52420 58240 52480
rect 63160 52590 63230 52600
rect 63160 52530 63220 52590
rect 63220 52530 63230 52590
rect 63160 52480 63230 52490
rect 63160 52420 63220 52480
rect 63220 52420 63230 52480
rect 68150 52590 68220 52600
rect 68150 52530 68210 52590
rect 68210 52530 68220 52590
rect 68150 52480 68220 52490
rect 68150 52420 68210 52480
rect 68210 52420 68220 52480
rect 73140 52590 73210 52600
rect 73140 52530 73200 52590
rect 73200 52530 73210 52590
rect 73140 52480 73210 52490
rect 73140 52420 73200 52480
rect 73200 52420 73210 52480
rect 78130 52590 78200 52600
rect 78130 52530 78190 52590
rect 78190 52530 78200 52590
rect 78130 52480 78200 52490
rect 78130 52420 78190 52480
rect 78190 52420 78200 52480
rect 46950 52320 47010 52380
rect 49590 52320 49650 52380
rect 52180 52320 52240 52380
rect 54340 52320 54400 52380
rect 57170 52320 57230 52380
rect 59330 52320 59390 52380
rect 62400 52320 62460 52380
rect 64080 52320 64140 52380
rect 67390 52320 67450 52380
rect 69070 52320 69130 52380
rect 72500 52320 72560 52380
rect 73940 52320 74000 52380
rect 77490 52320 77550 52380
rect 78930 52320 78990 52380
rect 43740 38630 43800 38690
rect 42440 36250 42500 36310
rect 48190 50880 48260 50890
rect 48190 50820 48250 50880
rect 48250 50820 48260 50880
rect 48190 50770 48260 50780
rect 48190 50710 48250 50770
rect 48250 50710 48260 50770
rect 47070 50610 47130 50670
rect 49470 50610 49530 50670
rect 48190 49170 48260 49180
rect 48190 49110 48250 49170
rect 48250 49110 48260 49170
rect 48190 49060 48260 49070
rect 48190 49000 48250 49060
rect 48250 49000 48260 49060
rect 47190 48900 47250 48960
rect 49350 48900 49410 48960
rect 48190 47460 48260 47470
rect 48190 47400 48250 47460
rect 48250 47400 48260 47460
rect 48190 47350 48260 47360
rect 48190 47290 48250 47350
rect 48250 47290 48260 47350
rect 47310 47190 47370 47250
rect 49230 47190 49290 47250
rect 46710 37650 46770 37710
rect 46650 37510 46710 37570
rect 46530 37370 46590 37430
rect 46470 37230 46530 37290
rect 48190 45750 48260 45760
rect 48190 45690 48250 45750
rect 48250 45690 48260 45750
rect 48190 45640 48260 45650
rect 48190 45580 48250 45640
rect 48250 45580 48260 45640
rect 47430 45480 47490 45540
rect 49110 45480 49170 45540
rect 48190 44040 48260 44050
rect 48190 43980 48250 44040
rect 48250 43980 48260 44040
rect 48190 43930 48260 43940
rect 48190 43870 48250 43930
rect 48250 43870 48260 43930
rect 47430 43770 47490 43830
rect 49110 43770 49170 43830
rect 46890 37090 46950 37150
rect 46830 36950 46890 37010
rect 48190 42330 48260 42340
rect 48190 42270 48250 42330
rect 48250 42270 48260 42330
rect 48190 42220 48260 42230
rect 48190 42160 48250 42220
rect 48250 42160 48260 42220
rect 47550 42060 47610 42120
rect 48990 42060 49050 42120
rect 48190 40620 48260 40630
rect 48190 40560 48250 40620
rect 48250 40560 48260 40620
rect 48190 40510 48260 40520
rect 48190 40450 48250 40510
rect 48250 40450 48260 40510
rect 47550 40350 47610 40410
rect 48990 40350 49050 40410
rect 47070 36810 47130 36870
rect 47010 36670 47070 36730
rect 47250 36530 47310 36590
rect 47190 36390 47250 36450
rect 42380 36110 42440 36170
rect 47660 38770 47720 38830
rect 53180 50880 53250 50890
rect 53180 50820 53240 50880
rect 53240 50820 53250 50880
rect 53180 50770 53250 50780
rect 53180 50710 53240 50770
rect 53240 50710 53250 50770
rect 58170 50880 58240 50890
rect 58170 50820 58230 50880
rect 58230 50820 58240 50880
rect 58170 50770 58240 50780
rect 58170 50710 58230 50770
rect 58230 50710 58240 50770
rect 63160 50880 63230 50890
rect 63160 50820 63220 50880
rect 63220 50820 63230 50880
rect 63160 50770 63230 50780
rect 63160 50710 63220 50770
rect 63220 50710 63230 50770
rect 68150 50880 68220 50890
rect 68150 50820 68210 50880
rect 68210 50820 68220 50880
rect 68150 50770 68220 50780
rect 68150 50710 68210 50770
rect 68210 50710 68220 50770
rect 73140 50880 73210 50890
rect 73140 50820 73200 50880
rect 73200 50820 73210 50880
rect 73140 50770 73210 50780
rect 73140 50710 73200 50770
rect 73200 50710 73210 50770
rect 78130 50880 78200 50890
rect 78130 50820 78190 50880
rect 78190 50820 78200 50880
rect 78130 50770 78200 50780
rect 78130 50710 78190 50770
rect 78190 50710 78200 50770
rect 52180 50610 52240 50670
rect 54340 50610 54400 50670
rect 57170 50610 57230 50670
rect 59330 50610 59390 50670
rect 62400 50610 62460 50670
rect 64080 50610 64140 50670
rect 67390 50610 67450 50670
rect 69070 50610 69130 50670
rect 72500 50610 72560 50670
rect 73940 50610 74000 50670
rect 77490 50610 77550 50670
rect 78930 50610 78990 50670
rect 53180 49170 53250 49180
rect 53180 49110 53240 49170
rect 53240 49110 53250 49170
rect 53180 49060 53250 49070
rect 53180 49000 53240 49060
rect 53240 49000 53250 49060
rect 58170 49170 58240 49180
rect 58170 49110 58230 49170
rect 58230 49110 58240 49170
rect 58170 49060 58240 49070
rect 58170 49000 58230 49060
rect 58230 49000 58240 49060
rect 63160 49170 63230 49180
rect 63160 49110 63220 49170
rect 63220 49110 63230 49170
rect 63160 49060 63230 49070
rect 63160 49000 63220 49060
rect 63220 49000 63230 49060
rect 68150 49170 68220 49180
rect 68150 49110 68210 49170
rect 68210 49110 68220 49170
rect 68150 49060 68220 49070
rect 68150 49000 68210 49060
rect 68210 49000 68220 49060
rect 73140 49170 73210 49180
rect 73140 49110 73200 49170
rect 73200 49110 73210 49170
rect 73140 49060 73210 49070
rect 73140 49000 73200 49060
rect 73200 49000 73210 49060
rect 78130 49170 78200 49180
rect 78130 49110 78190 49170
rect 78190 49110 78200 49170
rect 78130 49060 78200 49070
rect 78130 49000 78190 49060
rect 78190 49000 78200 49060
rect 52180 48900 52240 48960
rect 54340 48900 54400 48960
rect 57170 48900 57230 48960
rect 59330 48900 59390 48960
rect 62400 48900 62460 48960
rect 64080 48900 64140 48960
rect 67390 48900 67450 48960
rect 69070 48900 69130 48960
rect 72500 48900 72560 48960
rect 73940 48900 74000 48960
rect 77490 48900 77550 48960
rect 78930 48900 78990 48960
rect 48730 38630 48790 38690
rect 47430 36250 47490 36310
rect 53180 47460 53250 47470
rect 53180 47400 53240 47460
rect 53240 47400 53250 47460
rect 53180 47350 53250 47360
rect 53180 47290 53240 47350
rect 53240 47290 53250 47350
rect 52300 47190 52360 47250
rect 54220 47190 54280 47250
rect 53180 45750 53250 45760
rect 53180 45690 53240 45750
rect 53240 45690 53250 45750
rect 53180 45640 53250 45650
rect 53180 45580 53240 45640
rect 53240 45580 53250 45640
rect 52420 45480 52480 45540
rect 54100 45480 54160 45540
rect 53180 44040 53250 44050
rect 53180 43980 53240 44040
rect 53240 43980 53250 44040
rect 53180 43930 53250 43940
rect 53180 43870 53240 43930
rect 53240 43870 53250 43930
rect 52420 43770 52480 43830
rect 54100 43770 54160 43830
rect 53180 42330 53250 42340
rect 53180 42270 53240 42330
rect 53240 42270 53250 42330
rect 53180 42220 53250 42230
rect 53180 42160 53240 42220
rect 53240 42160 53250 42220
rect 52540 42060 52600 42120
rect 53980 42060 54040 42120
rect 53180 40620 53250 40630
rect 53180 40560 53240 40620
rect 53240 40560 53250 40620
rect 53180 40510 53250 40520
rect 53180 40450 53240 40510
rect 53240 40450 53250 40510
rect 52540 40350 52600 40410
rect 53980 40350 54040 40410
rect 52060 37090 52120 37150
rect 52000 36950 52060 37010
rect 51880 36810 51940 36870
rect 51820 36670 51880 36730
rect 52240 36530 52300 36590
rect 52180 36390 52240 36450
rect 47370 36110 47430 36170
rect 52650 38770 52710 38830
rect 58170 47460 58240 47470
rect 58170 47400 58230 47460
rect 58230 47400 58240 47460
rect 58170 47350 58240 47360
rect 58170 47290 58230 47350
rect 58230 47290 58240 47350
rect 57290 47190 57350 47250
rect 59210 47190 59270 47250
rect 53720 38630 53780 38690
rect 52420 36250 52480 36310
rect 58170 45750 58240 45760
rect 58170 45690 58230 45750
rect 58230 45690 58240 45750
rect 58170 45640 58240 45650
rect 58170 45580 58230 45640
rect 58230 45580 58240 45640
rect 57410 45480 57470 45540
rect 59090 45480 59150 45540
rect 58170 44040 58240 44050
rect 58170 43980 58230 44040
rect 58230 43980 58240 44040
rect 58170 43930 58240 43940
rect 58170 43870 58230 43930
rect 58230 43870 58240 43930
rect 57410 43770 57470 43830
rect 59090 43770 59150 43830
rect 58170 42330 58240 42340
rect 58170 42270 58230 42330
rect 58230 42270 58240 42330
rect 58170 42220 58240 42230
rect 58170 42160 58230 42220
rect 58230 42160 58240 42220
rect 57530 42060 57590 42120
rect 58970 42060 59030 42120
rect 58170 40620 58240 40630
rect 58170 40560 58230 40620
rect 58230 40560 58240 40620
rect 58170 40510 58240 40520
rect 58170 40450 58230 40510
rect 58230 40450 58240 40510
rect 57530 40350 57590 40410
rect 58970 40350 59030 40410
rect 57050 37090 57110 37150
rect 56990 36950 57050 37010
rect 56870 36810 56930 36870
rect 56810 36670 56870 36730
rect 57230 36530 57290 36590
rect 57170 36390 57230 36450
rect 52360 36110 52420 36170
rect 57640 38770 57700 38830
rect 63160 47460 63230 47470
rect 63160 47400 63220 47460
rect 63220 47400 63230 47460
rect 63160 47350 63230 47360
rect 63160 47290 63220 47350
rect 63220 47290 63230 47350
rect 68150 47460 68220 47470
rect 68150 47400 68210 47460
rect 68210 47400 68220 47460
rect 68150 47350 68220 47360
rect 68150 47290 68210 47350
rect 68210 47290 68220 47350
rect 73140 47460 73210 47470
rect 73140 47400 73200 47460
rect 73200 47400 73210 47460
rect 73140 47350 73210 47360
rect 73140 47290 73200 47350
rect 73200 47290 73210 47350
rect 78130 47460 78200 47470
rect 78130 47400 78190 47460
rect 78190 47400 78200 47460
rect 78130 47350 78200 47360
rect 78130 47290 78190 47350
rect 78190 47290 78200 47350
rect 62400 47190 62460 47250
rect 64080 47190 64140 47250
rect 67390 47190 67450 47250
rect 69070 47190 69130 47250
rect 72500 47190 72560 47250
rect 73940 47190 74000 47250
rect 77490 47190 77550 47250
rect 78930 47190 78990 47250
rect 58710 38630 58770 38690
rect 57410 36250 57470 36310
rect 63160 45750 63230 45760
rect 63160 45690 63220 45750
rect 63220 45690 63230 45750
rect 63160 45640 63230 45650
rect 63160 45580 63220 45640
rect 63220 45580 63230 45640
rect 62520 45480 62580 45540
rect 63960 45480 64020 45540
rect 63160 44040 63230 44050
rect 63160 43980 63220 44040
rect 63220 43980 63230 44040
rect 63160 43930 63230 43940
rect 63160 43870 63220 43930
rect 63220 43870 63230 43930
rect 62520 43770 62580 43830
rect 63960 43770 64020 43830
rect 63160 42330 63230 42340
rect 63160 42270 63220 42330
rect 63220 42270 63230 42330
rect 63160 42220 63230 42230
rect 63160 42160 63220 42220
rect 63220 42160 63230 42220
rect 62520 42060 62580 42120
rect 63960 42060 64020 42120
rect 63160 40620 63230 40630
rect 63160 40560 63220 40620
rect 63220 40560 63230 40620
rect 63160 40510 63230 40520
rect 63160 40450 63220 40510
rect 63220 40450 63230 40510
rect 62520 40350 62580 40410
rect 63960 40350 64020 40410
rect 62220 36530 62280 36590
rect 62160 36390 62220 36450
rect 57350 36110 57410 36170
rect 62630 38770 62690 38830
rect 68150 45750 68220 45760
rect 68150 45690 68210 45750
rect 68210 45690 68220 45750
rect 68150 45640 68220 45650
rect 68150 45580 68210 45640
rect 68210 45580 68220 45640
rect 67510 45480 67570 45540
rect 68950 45480 69010 45540
rect 68150 44040 68220 44050
rect 68150 43980 68210 44040
rect 68210 43980 68220 44040
rect 68150 43930 68220 43940
rect 68150 43870 68210 43930
rect 68210 43870 68220 43930
rect 67510 43770 67570 43830
rect 68950 43770 69010 43830
rect 68150 42330 68220 42340
rect 68150 42270 68210 42330
rect 68210 42270 68220 42330
rect 68150 42220 68220 42230
rect 68150 42160 68210 42220
rect 68210 42160 68220 42220
rect 67510 42060 67570 42120
rect 68950 42060 69010 42120
rect 68150 40620 68220 40630
rect 68150 40560 68210 40620
rect 68210 40560 68220 40620
rect 68150 40510 68220 40520
rect 68150 40450 68210 40510
rect 68210 40450 68220 40510
rect 67510 40350 67570 40410
rect 68950 40350 69010 40410
rect 63700 38630 63760 38690
rect 62400 36250 62460 36310
rect 67210 36530 67270 36590
rect 67150 36390 67210 36450
rect 62340 36110 62400 36170
rect 67620 38770 67680 38830
rect 73140 45750 73210 45760
rect 73140 45690 73200 45750
rect 73200 45690 73210 45750
rect 73140 45640 73210 45650
rect 73140 45580 73200 45640
rect 73200 45580 73210 45640
rect 78130 45750 78200 45760
rect 78130 45690 78190 45750
rect 78190 45690 78200 45750
rect 78130 45640 78200 45650
rect 78130 45580 78190 45640
rect 78190 45580 78200 45640
rect 72500 45480 72560 45540
rect 73940 45480 74000 45540
rect 77490 45480 77550 45540
rect 78930 45480 78990 45540
rect 73140 44040 73210 44050
rect 73140 43980 73200 44040
rect 73200 43980 73210 44040
rect 73140 43930 73210 43940
rect 73140 43870 73200 43930
rect 73200 43870 73210 43930
rect 78130 44040 78200 44050
rect 78130 43980 78190 44040
rect 78190 43980 78200 44040
rect 78130 43930 78200 43940
rect 78130 43870 78190 43930
rect 78190 43870 78200 43930
rect 72500 43770 72560 43830
rect 73940 43770 74000 43830
rect 77490 43770 77550 43830
rect 78930 43770 78990 43830
rect 73140 42330 73210 42340
rect 73140 42270 73200 42330
rect 73200 42270 73210 42330
rect 73140 42220 73210 42230
rect 73140 42160 73200 42220
rect 73200 42160 73210 42220
rect 78130 42330 78200 42340
rect 78130 42270 78190 42330
rect 78190 42270 78200 42330
rect 78130 42220 78200 42230
rect 78130 42160 78190 42220
rect 78190 42160 78200 42220
rect 72500 42060 72560 42120
rect 73940 42060 74000 42120
rect 77490 42060 77550 42120
rect 78930 42060 78990 42120
rect 73140 40620 73210 40630
rect 73140 40560 73200 40620
rect 73200 40560 73210 40620
rect 73140 40510 73210 40520
rect 73140 40450 73200 40510
rect 73200 40450 73210 40510
rect 78130 40620 78200 40630
rect 78130 40560 78190 40620
rect 78190 40560 78200 40620
rect 78130 40510 78200 40520
rect 78130 40450 78190 40510
rect 78190 40450 78200 40510
rect 72500 40350 72560 40410
rect 73940 40350 74000 40410
rect 77490 40350 77550 40410
rect 78930 40350 78990 40410
rect 68690 38630 68750 38690
rect 67390 36250 67450 36310
rect 67330 36110 67390 36170
rect 72610 38770 72670 38830
rect 73680 38630 73740 38690
rect 72380 36250 72440 36310
rect 72320 36110 72380 36170
rect 77600 38770 77660 38830
rect 78670 38630 78730 38690
rect 77370 36250 77430 36310
rect 77310 36110 77370 36170
rect 2360 30880 2420 30940
rect 2420 30740 2480 30800
rect 3720 28360 3780 28420
rect 2650 28220 2710 28280
rect 7350 30880 7410 30940
rect 7410 30740 7470 30800
rect 8710 28360 8770 28420
rect 7640 28220 7700 28280
rect 12340 30880 12400 30940
rect 12160 30600 12220 30660
rect 12220 30460 12280 30520
rect 12400 30740 12460 30800
rect 13700 28360 13760 28420
rect 12630 28220 12690 28280
rect 17330 30880 17390 30940
rect 17150 30600 17210 30660
rect 17210 30460 17270 30520
rect 17390 30740 17450 30800
rect 18690 28360 18750 28420
rect 17620 28220 17680 28280
rect 22320 30880 22380 30940
rect 22140 30600 22200 30660
rect 21780 30320 21840 30380
rect 21840 30180 21900 30240
rect 21960 30040 22020 30100
rect 22020 29900 22080 29960
rect 22200 30460 22260 30520
rect 22380 30740 22440 30800
rect 23680 28360 23740 28420
rect 22610 28220 22670 28280
rect 27310 30880 27370 30940
rect 27130 30600 27190 30660
rect 26770 30320 26830 30380
rect 26830 30180 26890 30240
rect 26950 30040 27010 30100
rect 27010 29900 27070 29960
rect 27190 30460 27250 30520
rect 27370 30740 27430 30800
rect 28670 28360 28730 28420
rect 27600 28220 27660 28280
rect 32300 30880 32360 30940
rect 32120 30600 32180 30660
rect 31940 30320 32000 30380
rect 31760 30040 31820 30100
rect 31400 29760 31460 29820
rect 31460 29620 31520 29680
rect 31580 29480 31640 29540
rect 31640 29340 31700 29400
rect 31820 29900 31880 29960
rect 32000 30180 32060 30240
rect 32180 30460 32240 30520
rect 32360 30740 32420 30800
rect 33660 28360 33720 28420
rect 32590 28220 32650 28280
rect 37290 30880 37350 30940
rect 37110 30600 37170 30660
rect 36930 30320 36990 30380
rect 36750 30040 36810 30100
rect 36570 29760 36630 29820
rect 36390 29200 36450 29260
rect 36210 28640 36270 28700
rect 36270 28500 36330 28560
rect 36450 29060 36510 29120
rect 36630 29620 36690 29680
rect 36810 29900 36870 29960
rect 36990 30180 37050 30240
rect 37170 30460 37230 30520
rect 37350 30740 37410 30800
rect 38650 28360 38710 28420
rect 37580 28220 37640 28280
rect 42280 30880 42340 30940
rect 42100 30600 42160 30660
rect 41920 30320 41980 30380
rect 41740 30040 41800 30100
rect 41560 29760 41620 29820
rect 41200 29200 41260 29260
rect 41260 29060 41320 29120
rect 41350 28920 41410 28980
rect 41440 28780 41500 28840
rect 41620 29620 41680 29680
rect 41800 29900 41860 29960
rect 41980 30180 42040 30240
rect 42160 30460 42220 30520
rect 42340 30740 42400 30800
rect 43640 28360 43700 28420
rect 42570 28220 42630 28280
rect 47270 30880 47330 30940
rect 47090 30600 47150 30660
rect 46910 30320 46970 30380
rect 46730 30040 46790 30100
rect 46370 29760 46430 29820
rect 46430 29620 46490 29680
rect 46550 29480 46610 29540
rect 46610 29340 46670 29400
rect 46790 29900 46850 29960
rect 46970 30180 47030 30240
rect 47150 30460 47210 30520
rect 47330 30740 47390 30800
rect 48630 28360 48690 28420
rect 47560 28220 47620 28280
rect 52260 30880 52320 30940
rect 52080 30600 52140 30660
rect 51720 30320 51780 30380
rect 51780 30180 51840 30240
rect 51900 30040 51960 30100
rect 51960 29900 52020 29960
rect 52140 30460 52200 30520
rect 52320 30740 52380 30800
rect 53620 28360 53680 28420
rect 52550 28220 52610 28280
rect 57250 30880 57310 30940
rect 57070 30600 57130 30660
rect 56710 30320 56770 30380
rect 56770 30180 56830 30240
rect 56890 30040 56950 30100
rect 56950 29900 57010 29960
rect 57130 30460 57190 30520
rect 57310 30740 57370 30800
rect 58610 28360 58670 28420
rect 57540 28220 57600 28280
rect 62240 30880 62300 30940
rect 62060 30600 62120 30660
rect 62120 30460 62180 30520
rect 62300 30740 62360 30800
rect 63600 28360 63660 28420
rect 62530 28220 62590 28280
rect 67230 30880 67290 30940
rect 67050 30600 67110 30660
rect 67110 30460 67170 30520
rect 67290 30740 67350 30800
rect 68590 28360 68650 28420
rect 67520 28220 67580 28280
rect 72220 30880 72280 30940
rect 72280 30740 72340 30800
rect 73580 28360 73640 28420
rect 72510 28220 72570 28280
rect 77210 30880 77270 30940
rect 77270 30740 77330 30800
rect 78570 28360 78630 28420
rect 77500 28220 77560 28280
<< metal3 >>
rect 100 66902 1872 66930
rect 100 65478 1788 66902
rect 1852 65478 1872 66902
rect 5090 66902 6862 66930
rect 2630 66580 2710 66590
rect 2630 66520 2640 66580
rect 2700 66520 2710 66580
rect 2630 66510 2710 66520
rect 2650 66070 2710 66510
rect 4070 66580 4150 66590
rect 4070 66520 4080 66580
rect 4140 66520 4150 66580
rect 4070 66510 4150 66520
rect 2630 66060 2710 66070
rect 3240 66280 3380 66310
rect 3240 66210 3270 66280
rect 3350 66210 3380 66280
rect 3240 66170 3380 66210
rect 3240 66100 3270 66170
rect 3350 66100 3380 66170
rect 3240 66060 3380 66100
rect 4070 66070 4130 66510
rect 4070 66060 4150 66070
rect 2630 66000 2640 66060
rect 2700 66000 2710 66060
rect 2630 65990 2710 66000
rect 100 65450 1872 65478
rect 100 65192 1872 65220
rect 100 63768 1788 65192
rect 1852 63768 1872 65192
rect 2650 64360 2710 65990
rect 4070 66000 4080 66060
rect 4140 66000 4150 66060
rect 4070 65990 4150 66000
rect 2630 64350 2710 64360
rect 3240 64570 3380 64600
rect 3240 64500 3270 64570
rect 3350 64500 3380 64570
rect 3240 64460 3380 64500
rect 3240 64390 3270 64460
rect 3350 64390 3380 64460
rect 3240 64350 3380 64390
rect 4070 64360 4130 65990
rect 5090 65478 6778 66902
rect 6842 65478 6862 66902
rect 10080 66902 11852 66930
rect 7620 66580 7700 66590
rect 7620 66520 7630 66580
rect 7690 66520 7700 66580
rect 7620 66510 7700 66520
rect 7640 66070 7700 66510
rect 9060 66580 9140 66590
rect 9060 66520 9070 66580
rect 9130 66520 9140 66580
rect 9060 66510 9140 66520
rect 7620 66060 7700 66070
rect 8230 66280 8370 66310
rect 8230 66210 8260 66280
rect 8340 66210 8370 66280
rect 8230 66170 8370 66210
rect 8230 66100 8260 66170
rect 8340 66100 8370 66170
rect 8230 66060 8370 66100
rect 9060 66070 9120 66510
rect 9060 66060 9140 66070
rect 7620 66000 7630 66060
rect 7690 66000 7700 66060
rect 7620 65990 7700 66000
rect 5090 65450 6862 65478
rect 5090 65192 6862 65220
rect 4070 64350 4150 64360
rect 2630 64290 2640 64350
rect 2700 64290 2710 64350
rect 2630 64280 2710 64290
rect 100 63740 1872 63768
rect 100 63482 1872 63510
rect 100 62058 1788 63482
rect 1852 62058 1872 63482
rect 2650 62650 2710 64280
rect 4070 64290 4080 64350
rect 4140 64290 4150 64350
rect 4070 64280 4150 64290
rect 2630 62640 2710 62650
rect 3240 62860 3380 62890
rect 3240 62790 3270 62860
rect 3350 62790 3380 62860
rect 3240 62750 3380 62790
rect 3240 62680 3270 62750
rect 3350 62680 3380 62750
rect 3240 62640 3380 62680
rect 4070 62650 4130 64280
rect 5090 63768 6778 65192
rect 6842 63768 6862 65192
rect 7640 64360 7700 65990
rect 9060 66000 9070 66060
rect 9130 66000 9140 66060
rect 9060 65990 9140 66000
rect 7620 64350 7700 64360
rect 8230 64570 8370 64600
rect 8230 64500 8260 64570
rect 8340 64500 8370 64570
rect 8230 64460 8370 64500
rect 8230 64390 8260 64460
rect 8340 64390 8370 64460
rect 8230 64350 8370 64390
rect 9060 64360 9120 65990
rect 10080 65478 11768 66902
rect 11832 65478 11852 66902
rect 15070 66902 16842 66930
rect 12610 66580 12690 66590
rect 12610 66520 12620 66580
rect 12680 66520 12690 66580
rect 12610 66510 12690 66520
rect 12630 66070 12690 66510
rect 14050 66580 14130 66590
rect 14050 66520 14060 66580
rect 14120 66520 14130 66580
rect 14050 66510 14130 66520
rect 12610 66060 12690 66070
rect 13220 66280 13360 66310
rect 13220 66210 13250 66280
rect 13330 66210 13360 66280
rect 13220 66170 13360 66210
rect 13220 66100 13250 66170
rect 13330 66100 13360 66170
rect 13220 66060 13360 66100
rect 14050 66070 14110 66510
rect 14050 66060 14130 66070
rect 12610 66000 12620 66060
rect 12680 66000 12690 66060
rect 12610 65990 12690 66000
rect 10080 65450 11852 65478
rect 10080 65192 11852 65220
rect 9060 64350 9140 64360
rect 7620 64290 7630 64350
rect 7690 64290 7700 64350
rect 7620 64280 7700 64290
rect 5090 63740 6862 63768
rect 5090 63482 6862 63510
rect 4070 62640 4150 62650
rect 2630 62580 2640 62640
rect 2700 62580 2710 62640
rect 2630 62570 2710 62580
rect 100 62030 1872 62058
rect 100 61772 1872 61800
rect 100 60348 1788 61772
rect 1852 60348 1872 61772
rect 2650 60940 2710 62570
rect 4070 62580 4080 62640
rect 4140 62580 4150 62640
rect 4070 62570 4150 62580
rect 2630 60930 2710 60940
rect 3240 61150 3380 61180
rect 3240 61080 3270 61150
rect 3350 61080 3380 61150
rect 3240 61040 3380 61080
rect 3240 60970 3270 61040
rect 3350 60970 3380 61040
rect 3240 60930 3380 60970
rect 4070 60940 4130 62570
rect 5090 62058 6778 63482
rect 6842 62058 6862 63482
rect 7640 62650 7700 64280
rect 9060 64290 9070 64350
rect 9130 64290 9140 64350
rect 9060 64280 9140 64290
rect 7620 62640 7700 62650
rect 8230 62860 8370 62890
rect 8230 62790 8260 62860
rect 8340 62790 8370 62860
rect 8230 62750 8370 62790
rect 8230 62680 8260 62750
rect 8340 62680 8370 62750
rect 8230 62640 8370 62680
rect 9060 62650 9120 64280
rect 10080 63768 11768 65192
rect 11832 63768 11852 65192
rect 12630 64360 12690 65990
rect 14050 66000 14060 66060
rect 14120 66000 14130 66060
rect 14050 65990 14130 66000
rect 12610 64350 12690 64360
rect 13220 64570 13360 64600
rect 13220 64500 13250 64570
rect 13330 64500 13360 64570
rect 13220 64460 13360 64500
rect 13220 64390 13250 64460
rect 13330 64390 13360 64460
rect 13220 64350 13360 64390
rect 14050 64360 14110 65990
rect 15070 65478 16758 66902
rect 16822 65478 16842 66902
rect 20060 66902 21832 66930
rect 17600 66580 17680 66590
rect 17600 66520 17610 66580
rect 17670 66520 17680 66580
rect 17600 66510 17680 66520
rect 17620 66070 17680 66510
rect 19040 66580 19120 66590
rect 19040 66520 19050 66580
rect 19110 66520 19120 66580
rect 19040 66510 19120 66520
rect 17600 66060 17680 66070
rect 18210 66280 18350 66310
rect 18210 66210 18240 66280
rect 18320 66210 18350 66280
rect 18210 66170 18350 66210
rect 18210 66100 18240 66170
rect 18320 66100 18350 66170
rect 18210 66060 18350 66100
rect 19040 66070 19100 66510
rect 19040 66060 19120 66070
rect 17600 66000 17610 66060
rect 17670 66000 17680 66060
rect 17600 65990 17680 66000
rect 15070 65450 16842 65478
rect 15070 65192 16842 65220
rect 14050 64350 14130 64360
rect 12610 64290 12620 64350
rect 12680 64290 12690 64350
rect 12610 64280 12690 64290
rect 10080 63740 11852 63768
rect 10080 63482 11852 63510
rect 9060 62640 9140 62650
rect 7620 62580 7630 62640
rect 7690 62580 7700 62640
rect 7620 62570 7700 62580
rect 5090 62030 6862 62058
rect 5090 61772 6862 61800
rect 4070 60930 4150 60940
rect 2630 60870 2640 60930
rect 2700 60870 2710 60930
rect 2630 60860 2710 60870
rect 100 60320 1872 60348
rect 100 60062 1872 60090
rect 100 58638 1788 60062
rect 1852 58638 1872 60062
rect 2650 59230 2710 60860
rect 4070 60870 4080 60930
rect 4140 60870 4150 60930
rect 4070 60860 4150 60870
rect 2630 59220 2710 59230
rect 3240 59440 3380 59470
rect 3240 59370 3270 59440
rect 3350 59370 3380 59440
rect 3240 59330 3380 59370
rect 3240 59260 3270 59330
rect 3350 59260 3380 59330
rect 3240 59220 3380 59260
rect 4070 59230 4130 60860
rect 5090 60348 6778 61772
rect 6842 60348 6862 61772
rect 7640 60940 7700 62570
rect 9060 62580 9070 62640
rect 9130 62580 9140 62640
rect 9060 62570 9140 62580
rect 7620 60930 7700 60940
rect 8230 61150 8370 61180
rect 8230 61080 8260 61150
rect 8340 61080 8370 61150
rect 8230 61040 8370 61080
rect 8230 60970 8260 61040
rect 8340 60970 8370 61040
rect 8230 60930 8370 60970
rect 9060 60940 9120 62570
rect 10080 62058 11768 63482
rect 11832 62058 11852 63482
rect 12630 62650 12690 64280
rect 14050 64290 14060 64350
rect 14120 64290 14130 64350
rect 14050 64280 14130 64290
rect 12610 62640 12690 62650
rect 13220 62860 13360 62890
rect 13220 62790 13250 62860
rect 13330 62790 13360 62860
rect 13220 62750 13360 62790
rect 13220 62680 13250 62750
rect 13330 62680 13360 62750
rect 13220 62640 13360 62680
rect 14050 62650 14110 64280
rect 15070 63768 16758 65192
rect 16822 63768 16842 65192
rect 17620 64360 17680 65990
rect 19040 66000 19050 66060
rect 19110 66000 19120 66060
rect 19040 65990 19120 66000
rect 17600 64350 17680 64360
rect 18210 64570 18350 64600
rect 18210 64500 18240 64570
rect 18320 64500 18350 64570
rect 18210 64460 18350 64500
rect 18210 64390 18240 64460
rect 18320 64390 18350 64460
rect 18210 64350 18350 64390
rect 19040 64360 19100 65990
rect 20060 65478 21748 66902
rect 21812 65478 21832 66902
rect 25050 66902 26822 66930
rect 22590 66580 22670 66590
rect 22590 66520 22600 66580
rect 22660 66520 22670 66580
rect 22590 66510 22670 66520
rect 22610 66070 22670 66510
rect 24030 66580 24110 66590
rect 24030 66520 24040 66580
rect 24100 66520 24110 66580
rect 24030 66510 24110 66520
rect 22590 66060 22670 66070
rect 23200 66280 23340 66310
rect 23200 66210 23230 66280
rect 23310 66210 23340 66280
rect 23200 66170 23340 66210
rect 23200 66100 23230 66170
rect 23310 66100 23340 66170
rect 23200 66060 23340 66100
rect 24030 66070 24090 66510
rect 24030 66060 24110 66070
rect 22590 66000 22600 66060
rect 22660 66000 22670 66060
rect 22590 65990 22670 66000
rect 20060 65450 21832 65478
rect 20060 65192 21832 65220
rect 19040 64350 19120 64360
rect 17600 64290 17610 64350
rect 17670 64290 17680 64350
rect 17600 64280 17680 64290
rect 15070 63740 16842 63768
rect 15070 63482 16842 63510
rect 14050 62640 14130 62650
rect 12610 62580 12620 62640
rect 12680 62580 12690 62640
rect 12610 62570 12690 62580
rect 10080 62030 11852 62058
rect 10080 61772 11852 61800
rect 9060 60930 9140 60940
rect 7620 60870 7630 60930
rect 7690 60870 7700 60930
rect 7620 60860 7700 60870
rect 5090 60320 6862 60348
rect 5090 60062 6862 60090
rect 4070 59220 4150 59230
rect 2630 59160 2640 59220
rect 2700 59160 2710 59220
rect 2630 59150 2710 59160
rect 100 58610 1872 58638
rect 100 58352 1872 58380
rect 100 56928 1788 58352
rect 1852 56928 1872 58352
rect 2650 57520 2710 59150
rect 4070 59160 4080 59220
rect 4140 59160 4150 59220
rect 4070 59150 4150 59160
rect 2630 57510 2710 57520
rect 3240 57730 3380 57760
rect 3240 57660 3270 57730
rect 3350 57660 3380 57730
rect 3240 57620 3380 57660
rect 3240 57550 3270 57620
rect 3350 57550 3380 57620
rect 3240 57510 3380 57550
rect 4070 57520 4130 59150
rect 5090 58638 6778 60062
rect 6842 58638 6862 60062
rect 7640 59230 7700 60860
rect 9060 60870 9070 60930
rect 9130 60870 9140 60930
rect 9060 60860 9140 60870
rect 7620 59220 7700 59230
rect 8230 59440 8370 59470
rect 8230 59370 8260 59440
rect 8340 59370 8370 59440
rect 8230 59330 8370 59370
rect 8230 59260 8260 59330
rect 8340 59260 8370 59330
rect 8230 59220 8370 59260
rect 9060 59230 9120 60860
rect 10080 60348 11768 61772
rect 11832 60348 11852 61772
rect 12630 60940 12690 62570
rect 14050 62580 14060 62640
rect 14120 62580 14130 62640
rect 14050 62570 14130 62580
rect 12610 60930 12690 60940
rect 13220 61150 13360 61180
rect 13220 61080 13250 61150
rect 13330 61080 13360 61150
rect 13220 61040 13360 61080
rect 13220 60970 13250 61040
rect 13330 60970 13360 61040
rect 13220 60930 13360 60970
rect 14050 60940 14110 62570
rect 15070 62058 16758 63482
rect 16822 62058 16842 63482
rect 17620 62650 17680 64280
rect 19040 64290 19050 64350
rect 19110 64290 19120 64350
rect 19040 64280 19120 64290
rect 17600 62640 17680 62650
rect 18210 62860 18350 62890
rect 18210 62790 18240 62860
rect 18320 62790 18350 62860
rect 18210 62750 18350 62790
rect 18210 62680 18240 62750
rect 18320 62680 18350 62750
rect 18210 62640 18350 62680
rect 19040 62650 19100 64280
rect 20060 63768 21748 65192
rect 21812 63768 21832 65192
rect 22610 64360 22670 65990
rect 24030 66000 24040 66060
rect 24100 66000 24110 66060
rect 24030 65990 24110 66000
rect 22590 64350 22670 64360
rect 23200 64570 23340 64600
rect 23200 64500 23230 64570
rect 23310 64500 23340 64570
rect 23200 64460 23340 64500
rect 23200 64390 23230 64460
rect 23310 64390 23340 64460
rect 23200 64350 23340 64390
rect 24030 64360 24090 65990
rect 25050 65478 26738 66902
rect 26802 65478 26822 66902
rect 30040 66902 31812 66930
rect 27580 66580 27660 66590
rect 27580 66520 27590 66580
rect 27650 66520 27660 66580
rect 27580 66510 27660 66520
rect 27600 66070 27660 66510
rect 29020 66580 29100 66590
rect 29020 66520 29030 66580
rect 29090 66520 29100 66580
rect 29020 66510 29100 66520
rect 27580 66060 27660 66070
rect 28190 66280 28330 66310
rect 28190 66210 28220 66280
rect 28300 66210 28330 66280
rect 28190 66170 28330 66210
rect 28190 66100 28220 66170
rect 28300 66100 28330 66170
rect 28190 66060 28330 66100
rect 29020 66070 29080 66510
rect 29020 66060 29100 66070
rect 27580 66000 27590 66060
rect 27650 66000 27660 66060
rect 27580 65990 27660 66000
rect 25050 65450 26822 65478
rect 25050 65192 26822 65220
rect 24030 64350 24110 64360
rect 22590 64290 22600 64350
rect 22660 64290 22670 64350
rect 22590 64280 22670 64290
rect 20060 63740 21832 63768
rect 20060 63482 21832 63510
rect 19040 62640 19120 62650
rect 17600 62580 17610 62640
rect 17670 62580 17680 62640
rect 17600 62570 17680 62580
rect 15070 62030 16842 62058
rect 15070 61772 16842 61800
rect 14050 60930 14130 60940
rect 12610 60870 12620 60930
rect 12680 60870 12690 60930
rect 12610 60860 12690 60870
rect 10080 60320 11852 60348
rect 10080 60062 11852 60090
rect 9060 59220 9140 59230
rect 7620 59160 7630 59220
rect 7690 59160 7700 59220
rect 7620 59150 7700 59160
rect 5090 58610 6862 58638
rect 5090 58352 6862 58380
rect 4070 57510 4150 57520
rect 2630 57450 2640 57510
rect 2700 57450 2710 57510
rect 2630 57440 2710 57450
rect 100 56900 1872 56928
rect 100 56642 1872 56670
rect 100 55218 1788 56642
rect 1852 55218 1872 56642
rect 2650 55810 2710 57440
rect 4070 57450 4080 57510
rect 4140 57450 4150 57510
rect 4070 57440 4150 57450
rect 2630 55800 2710 55810
rect 3240 56020 3380 56050
rect 3240 55950 3270 56020
rect 3350 55950 3380 56020
rect 3240 55910 3380 55950
rect 3240 55840 3270 55910
rect 3350 55840 3380 55910
rect 3240 55800 3380 55840
rect 4070 55810 4130 57440
rect 5090 56928 6778 58352
rect 6842 56928 6862 58352
rect 7640 57520 7700 59150
rect 9060 59160 9070 59220
rect 9130 59160 9140 59220
rect 9060 59150 9140 59160
rect 7620 57510 7700 57520
rect 8230 57730 8370 57760
rect 8230 57660 8260 57730
rect 8340 57660 8370 57730
rect 8230 57620 8370 57660
rect 8230 57550 8260 57620
rect 8340 57550 8370 57620
rect 8230 57510 8370 57550
rect 9060 57520 9120 59150
rect 10080 58638 11768 60062
rect 11832 58638 11852 60062
rect 12490 59740 12570 59750
rect 12490 59680 12500 59740
rect 12560 59680 12570 59740
rect 12490 59670 12570 59680
rect 12510 59230 12570 59670
rect 12490 59220 12570 59230
rect 12490 59160 12500 59220
rect 12560 59160 12570 59220
rect 12490 59150 12570 59160
rect 10080 58610 11852 58638
rect 10080 58352 11852 58380
rect 9060 57510 9140 57520
rect 7620 57450 7630 57510
rect 7690 57450 7700 57510
rect 7620 57440 7700 57450
rect 5090 56900 6862 56928
rect 5090 56642 6862 56670
rect 4070 55800 4150 55810
rect 2630 55740 2640 55800
rect 2700 55740 2710 55800
rect 2630 55730 2710 55740
rect 100 55190 1872 55218
rect 100 54932 1872 54960
rect 100 53508 1788 54932
rect 1852 53508 1872 54932
rect 2650 54100 2710 55730
rect 4070 55740 4080 55800
rect 4140 55740 4150 55800
rect 4070 55730 4150 55740
rect 2630 54090 2710 54100
rect 3240 54310 3380 54340
rect 3240 54240 3270 54310
rect 3350 54240 3380 54310
rect 3240 54200 3380 54240
rect 3240 54130 3270 54200
rect 3350 54130 3380 54200
rect 3240 54090 3380 54130
rect 4070 54100 4130 55730
rect 5090 55218 6778 56642
rect 6842 55218 6862 56642
rect 7640 55810 7700 57440
rect 9060 57450 9070 57510
rect 9130 57450 9140 57510
rect 9060 57440 9140 57450
rect 7620 55800 7700 55810
rect 8230 56020 8370 56050
rect 8230 55950 8260 56020
rect 8340 55950 8370 56020
rect 8230 55910 8370 55950
rect 8230 55840 8260 55910
rect 8340 55840 8370 55910
rect 8230 55800 8370 55840
rect 9060 55810 9120 57440
rect 10080 56928 11768 58352
rect 11832 56928 11852 58352
rect 12510 57520 12570 59150
rect 12490 57510 12570 57520
rect 12490 57450 12500 57510
rect 12560 57450 12570 57510
rect 12490 57440 12570 57450
rect 10080 56900 11852 56928
rect 10080 56642 11852 56670
rect 9060 55800 9140 55810
rect 7620 55740 7630 55800
rect 7690 55740 7700 55800
rect 7620 55730 7700 55740
rect 5090 55190 6862 55218
rect 5090 54932 6862 54960
rect 4070 54090 4150 54100
rect 2630 54030 2640 54090
rect 2700 54030 2710 54090
rect 2630 54020 2710 54030
rect 100 53480 1872 53508
rect 100 53222 1872 53250
rect 100 51798 1788 53222
rect 1852 51798 1872 53222
rect 2650 52390 2710 54020
rect 4070 54030 4080 54090
rect 4140 54030 4150 54090
rect 4070 54020 4150 54030
rect 2630 52380 2710 52390
rect 3240 52600 3380 52630
rect 3240 52530 3270 52600
rect 3350 52530 3380 52600
rect 3240 52490 3380 52530
rect 3240 52420 3270 52490
rect 3350 52420 3380 52490
rect 3240 52380 3380 52420
rect 4070 52390 4130 54020
rect 5090 53508 6778 54932
rect 6842 53508 6862 54932
rect 7640 54100 7700 55730
rect 9060 55740 9070 55800
rect 9130 55740 9140 55800
rect 9060 55730 9140 55740
rect 7620 54090 7700 54100
rect 8230 54310 8370 54340
rect 8230 54240 8260 54310
rect 8340 54240 8370 54310
rect 8230 54200 8370 54240
rect 8230 54130 8260 54200
rect 8340 54130 8370 54200
rect 8230 54090 8370 54130
rect 9060 54100 9120 55730
rect 10080 55218 11768 56642
rect 11832 55218 11852 56642
rect 12510 55810 12570 57440
rect 12490 55800 12570 55810
rect 12490 55740 12500 55800
rect 12560 55740 12570 55800
rect 12490 55730 12570 55740
rect 10080 55190 11852 55218
rect 10080 54932 11852 54960
rect 9060 54090 9140 54100
rect 7620 54030 7630 54090
rect 7690 54030 7700 54090
rect 7620 54020 7700 54030
rect 5090 53480 6862 53508
rect 5090 53222 6862 53250
rect 4070 52380 4150 52390
rect 2630 52320 2640 52380
rect 2700 52320 2710 52380
rect 2630 52310 2710 52320
rect 100 51770 1872 51798
rect 100 51512 1872 51540
rect 100 50088 1788 51512
rect 1852 50088 1872 51512
rect 2650 50680 2710 52310
rect 4070 52320 4080 52380
rect 4140 52320 4150 52380
rect 4070 52310 4150 52320
rect 2630 50670 2710 50680
rect 3240 50890 3380 50920
rect 3240 50820 3270 50890
rect 3350 50820 3380 50890
rect 3240 50780 3380 50820
rect 3240 50710 3270 50780
rect 3350 50710 3380 50780
rect 3240 50670 3380 50710
rect 4070 50680 4130 52310
rect 5090 51798 6778 53222
rect 6842 51798 6862 53222
rect 7640 52390 7700 54020
rect 9060 54030 9070 54090
rect 9130 54030 9140 54090
rect 9060 54020 9140 54030
rect 7620 52380 7700 52390
rect 8230 52600 8370 52630
rect 8230 52530 8260 52600
rect 8340 52530 8370 52600
rect 8230 52490 8370 52530
rect 8230 52420 8260 52490
rect 8340 52420 8370 52490
rect 8230 52380 8370 52420
rect 9060 52390 9120 54020
rect 10080 53508 11768 54932
rect 11832 53508 11852 54932
rect 12510 54100 12570 55730
rect 12490 54090 12570 54100
rect 12490 54030 12500 54090
rect 12560 54030 12570 54090
rect 12490 54020 12570 54030
rect 10080 53480 11852 53508
rect 10080 53222 11852 53250
rect 9060 52380 9140 52390
rect 7620 52320 7630 52380
rect 7690 52320 7700 52380
rect 7620 52310 7700 52320
rect 5090 51770 6862 51798
rect 5090 51512 6862 51540
rect 4070 50670 4150 50680
rect 2630 50610 2640 50670
rect 2700 50610 2710 50670
rect 2630 50600 2710 50610
rect 100 50060 1872 50088
rect 100 49802 1872 49830
rect 100 48378 1788 49802
rect 1852 48378 1872 49802
rect 2650 48970 2710 50600
rect 4070 50610 4080 50670
rect 4140 50610 4150 50670
rect 4070 50600 4150 50610
rect 2630 48960 2710 48970
rect 3240 49180 3380 49210
rect 3240 49110 3270 49180
rect 3350 49110 3380 49180
rect 3240 49070 3380 49110
rect 3240 49000 3270 49070
rect 3350 49000 3380 49070
rect 3240 48960 3380 49000
rect 4070 48970 4130 50600
rect 5090 50088 6778 51512
rect 6842 50088 6862 51512
rect 7640 50680 7700 52310
rect 9060 52320 9070 52380
rect 9130 52320 9140 52380
rect 9060 52310 9140 52320
rect 7620 50670 7700 50680
rect 8230 50890 8370 50920
rect 8230 50820 8260 50890
rect 8340 50820 8370 50890
rect 8230 50780 8370 50820
rect 8230 50710 8260 50780
rect 8340 50710 8370 50780
rect 8230 50670 8370 50710
rect 9060 50680 9120 52310
rect 10080 51798 11768 53222
rect 11832 51798 11852 53222
rect 12510 52390 12570 54020
rect 12490 52380 12570 52390
rect 12490 52320 12500 52380
rect 12560 52320 12570 52380
rect 12490 52310 12570 52320
rect 10080 51770 11852 51798
rect 10080 51512 11852 51540
rect 9060 50670 9140 50680
rect 7620 50610 7630 50670
rect 7690 50610 7700 50670
rect 7620 50600 7700 50610
rect 5090 50060 6862 50088
rect 5090 49802 6862 49830
rect 4070 48960 4150 48970
rect 2630 48900 2640 48960
rect 2700 48900 2710 48960
rect 2630 48890 2710 48900
rect 100 48350 1872 48378
rect 100 48092 1872 48120
rect 100 46668 1788 48092
rect 1852 46668 1872 48092
rect 2650 47260 2710 48890
rect 4070 48900 4080 48960
rect 4140 48900 4150 48960
rect 4070 48890 4150 48900
rect 2630 47250 2710 47260
rect 3240 47470 3380 47500
rect 3240 47400 3270 47470
rect 3350 47400 3380 47470
rect 3240 47360 3380 47400
rect 3240 47290 3270 47360
rect 3350 47290 3380 47360
rect 3240 47250 3380 47290
rect 4070 47260 4130 48890
rect 5090 48378 6778 49802
rect 6842 48378 6862 49802
rect 7640 48970 7700 50600
rect 9060 50610 9070 50670
rect 9130 50610 9140 50670
rect 9060 50600 9140 50610
rect 7620 48960 7700 48970
rect 8230 49180 8370 49210
rect 8230 49110 8260 49180
rect 8340 49110 8370 49180
rect 8230 49070 8370 49110
rect 8230 49000 8260 49070
rect 8340 49000 8370 49070
rect 8230 48960 8370 49000
rect 9060 48970 9120 50600
rect 10080 50088 11768 51512
rect 11832 50088 11852 51512
rect 12510 50680 12570 52310
rect 12490 50670 12570 50680
rect 12490 50610 12500 50670
rect 12560 50610 12570 50670
rect 12490 50600 12570 50610
rect 10080 50060 11852 50088
rect 10080 49802 11852 49830
rect 9060 48960 9140 48970
rect 7620 48900 7630 48960
rect 7690 48900 7700 48960
rect 7620 48890 7700 48900
rect 5090 48350 6862 48378
rect 5090 48092 6862 48120
rect 4070 47250 4150 47260
rect 2630 47190 2640 47250
rect 2700 47190 2710 47250
rect 2630 47180 2710 47190
rect 100 46640 1872 46668
rect 100 46382 1872 46410
rect 100 44958 1788 46382
rect 1852 44958 1872 46382
rect 2650 45550 2710 47180
rect 4070 47190 4080 47250
rect 4140 47190 4150 47250
rect 4070 47180 4150 47190
rect 2630 45540 2710 45550
rect 3240 45760 3380 45790
rect 3240 45690 3270 45760
rect 3350 45690 3380 45760
rect 3240 45650 3380 45690
rect 3240 45580 3270 45650
rect 3350 45580 3380 45650
rect 3240 45540 3380 45580
rect 4070 45550 4130 47180
rect 5090 46668 6778 48092
rect 6842 46668 6862 48092
rect 7640 47260 7700 48890
rect 9060 48900 9070 48960
rect 9130 48900 9140 48960
rect 9060 48890 9140 48900
rect 7620 47250 7700 47260
rect 8230 47470 8370 47500
rect 8230 47400 8260 47470
rect 8340 47400 8370 47470
rect 8230 47360 8370 47400
rect 8230 47290 8260 47360
rect 8340 47290 8370 47360
rect 8230 47250 8370 47290
rect 9060 47260 9120 48890
rect 10080 48378 11768 49802
rect 11832 48378 11852 49802
rect 12510 48970 12570 50600
rect 12490 48960 12570 48970
rect 12490 48900 12500 48960
rect 12560 48900 12570 48960
rect 12490 48890 12570 48900
rect 10080 48350 11852 48378
rect 10080 48092 11852 48120
rect 9060 47250 9140 47260
rect 7620 47190 7630 47250
rect 7690 47190 7700 47250
rect 7620 47180 7700 47190
rect 5090 46640 6862 46668
rect 5090 46382 6862 46410
rect 4070 45540 4150 45550
rect 2630 45480 2640 45540
rect 2700 45480 2710 45540
rect 2630 45470 2710 45480
rect 100 44930 1872 44958
rect 100 44672 1872 44700
rect 100 43248 1788 44672
rect 1852 43248 1872 44672
rect 2650 43840 2710 45470
rect 4070 45480 4080 45540
rect 4140 45480 4150 45540
rect 4070 45470 4150 45480
rect 2630 43830 2710 43840
rect 3240 44050 3380 44080
rect 3240 43980 3270 44050
rect 3350 43980 3380 44050
rect 3240 43940 3380 43980
rect 3240 43870 3270 43940
rect 3350 43870 3380 43940
rect 3240 43830 3380 43870
rect 4070 43840 4130 45470
rect 5090 44958 6778 46382
rect 6842 44958 6862 46382
rect 7640 45550 7700 47180
rect 9060 47190 9070 47250
rect 9130 47190 9140 47250
rect 9060 47180 9140 47190
rect 7620 45540 7700 45550
rect 8230 45760 8370 45790
rect 8230 45690 8260 45760
rect 8340 45690 8370 45760
rect 8230 45650 8370 45690
rect 8230 45580 8260 45650
rect 8340 45580 8370 45650
rect 8230 45540 8370 45580
rect 9060 45550 9120 47180
rect 10080 46668 11768 48092
rect 11832 46668 11852 48092
rect 12510 47260 12570 48890
rect 12490 47250 12570 47260
rect 12490 47190 12500 47250
rect 12560 47190 12570 47250
rect 12490 47180 12570 47190
rect 10080 46640 11852 46668
rect 10080 46382 11852 46410
rect 9060 45540 9140 45550
rect 7620 45480 7630 45540
rect 7690 45480 7700 45540
rect 7620 45470 7700 45480
rect 5090 44930 6862 44958
rect 5090 44672 6862 44700
rect 4070 43830 4150 43840
rect 2630 43770 2640 43830
rect 2700 43770 2710 43830
rect 2630 43760 2710 43770
rect 100 43220 1872 43248
rect 100 42962 1872 42990
rect 100 41538 1788 42962
rect 1852 41538 1872 42962
rect 2650 42130 2710 43760
rect 4070 43770 4080 43830
rect 4140 43770 4150 43830
rect 4070 43760 4150 43770
rect 2630 42120 2710 42130
rect 3240 42340 3380 42370
rect 3240 42270 3270 42340
rect 3350 42270 3380 42340
rect 3240 42230 3380 42270
rect 3240 42160 3270 42230
rect 3350 42160 3380 42230
rect 3240 42120 3380 42160
rect 4070 42130 4130 43760
rect 5090 43248 6778 44672
rect 6842 43248 6862 44672
rect 7640 43840 7700 45470
rect 9060 45480 9070 45540
rect 9130 45480 9140 45540
rect 9060 45470 9140 45480
rect 7620 43830 7700 43840
rect 8230 44050 8370 44080
rect 8230 43980 8260 44050
rect 8340 43980 8370 44050
rect 8230 43940 8370 43980
rect 8230 43870 8260 43940
rect 8340 43870 8370 43940
rect 8230 43830 8370 43870
rect 9060 43840 9120 45470
rect 10080 44958 11768 46382
rect 11832 44958 11852 46382
rect 12630 45550 12690 60860
rect 14050 60870 14060 60930
rect 14120 60870 14130 60930
rect 14050 60860 14130 60870
rect 13220 59440 13360 59470
rect 13220 59370 13250 59440
rect 13330 59370 13360 59440
rect 13220 59330 13360 59370
rect 13220 59260 13250 59330
rect 13330 59260 13360 59330
rect 13220 59220 13360 59260
rect 13220 57730 13360 57760
rect 13220 57660 13250 57730
rect 13330 57660 13360 57730
rect 13220 57620 13360 57660
rect 13220 57550 13250 57620
rect 13330 57550 13360 57620
rect 13220 57510 13360 57550
rect 13220 56020 13360 56050
rect 13220 55950 13250 56020
rect 13330 55950 13360 56020
rect 13220 55910 13360 55950
rect 13220 55840 13250 55910
rect 13330 55840 13360 55910
rect 13220 55800 13360 55840
rect 13220 54310 13360 54340
rect 13220 54240 13250 54310
rect 13330 54240 13360 54310
rect 13220 54200 13360 54240
rect 13220 54130 13250 54200
rect 13330 54130 13360 54200
rect 13220 54090 13360 54130
rect 13220 52600 13360 52630
rect 13220 52530 13250 52600
rect 13330 52530 13360 52600
rect 13220 52490 13360 52530
rect 13220 52420 13250 52490
rect 13330 52420 13360 52490
rect 13220 52380 13360 52420
rect 13220 50890 13360 50920
rect 13220 50820 13250 50890
rect 13330 50820 13360 50890
rect 13220 50780 13360 50820
rect 13220 50710 13250 50780
rect 13330 50710 13360 50780
rect 13220 50670 13360 50710
rect 13220 49180 13360 49210
rect 13220 49110 13250 49180
rect 13330 49110 13360 49180
rect 13220 49070 13360 49110
rect 13220 49000 13250 49070
rect 13330 49000 13360 49070
rect 13220 48960 13360 49000
rect 13220 47470 13360 47500
rect 13220 47400 13250 47470
rect 13330 47400 13360 47470
rect 13220 47360 13360 47400
rect 13220 47290 13250 47360
rect 13330 47290 13360 47360
rect 13220 47250 13360 47290
rect 12610 45540 12690 45550
rect 13220 45760 13360 45790
rect 13220 45690 13250 45760
rect 13330 45690 13360 45760
rect 13220 45650 13360 45690
rect 13220 45580 13250 45650
rect 13330 45580 13360 45650
rect 13220 45540 13360 45580
rect 14050 45550 14110 60860
rect 15070 60348 16758 61772
rect 16822 60348 16842 61772
rect 17620 60940 17680 62570
rect 19040 62580 19050 62640
rect 19110 62580 19120 62640
rect 19040 62570 19120 62580
rect 17600 60930 17680 60940
rect 18210 61150 18350 61180
rect 18210 61080 18240 61150
rect 18320 61080 18350 61150
rect 18210 61040 18350 61080
rect 18210 60970 18240 61040
rect 18320 60970 18350 61040
rect 18210 60930 18350 60970
rect 19040 60940 19100 62570
rect 20060 62058 21748 63482
rect 21812 62058 21832 63482
rect 22470 63160 22550 63170
rect 22470 63100 22480 63160
rect 22540 63100 22550 63160
rect 22470 63090 22550 63100
rect 22490 62650 22550 63090
rect 22470 62640 22550 62650
rect 22470 62580 22480 62640
rect 22540 62580 22550 62640
rect 22470 62570 22550 62580
rect 20060 62030 21832 62058
rect 20060 61772 21832 61800
rect 19040 60930 19120 60940
rect 17600 60870 17610 60930
rect 17670 60870 17680 60930
rect 17600 60860 17680 60870
rect 15070 60320 16842 60348
rect 15070 60062 16842 60090
rect 14170 59740 14250 59750
rect 14170 59680 14180 59740
rect 14240 59680 14250 59740
rect 14170 59670 14250 59680
rect 14170 59230 14230 59670
rect 14170 59220 14250 59230
rect 14170 59160 14180 59220
rect 14240 59160 14250 59220
rect 14170 59150 14250 59160
rect 14170 57520 14230 59150
rect 15070 58638 16758 60062
rect 16822 58638 16842 60062
rect 17480 59740 17560 59750
rect 17480 59680 17490 59740
rect 17550 59680 17560 59740
rect 17480 59670 17560 59680
rect 17500 59230 17560 59670
rect 17480 59220 17560 59230
rect 17480 59160 17490 59220
rect 17550 59160 17560 59220
rect 17480 59150 17560 59160
rect 15070 58610 16842 58638
rect 15070 58352 16842 58380
rect 14170 57510 14250 57520
rect 14170 57450 14180 57510
rect 14240 57450 14250 57510
rect 14170 57440 14250 57450
rect 14170 55810 14230 57440
rect 15070 56928 16758 58352
rect 16822 56928 16842 58352
rect 17500 57520 17560 59150
rect 17480 57510 17560 57520
rect 17480 57450 17490 57510
rect 17550 57450 17560 57510
rect 17480 57440 17560 57450
rect 15070 56900 16842 56928
rect 15070 56642 16842 56670
rect 14170 55800 14250 55810
rect 14170 55740 14180 55800
rect 14240 55740 14250 55800
rect 14170 55730 14250 55740
rect 14170 54100 14230 55730
rect 15070 55218 16758 56642
rect 16822 55218 16842 56642
rect 17500 55810 17560 57440
rect 17480 55800 17560 55810
rect 17480 55740 17490 55800
rect 17550 55740 17560 55800
rect 17480 55730 17560 55740
rect 15070 55190 16842 55218
rect 15070 54932 16842 54960
rect 14170 54090 14250 54100
rect 14170 54030 14180 54090
rect 14240 54030 14250 54090
rect 14170 54020 14250 54030
rect 14170 52390 14230 54020
rect 15070 53508 16758 54932
rect 16822 53508 16842 54932
rect 17500 54100 17560 55730
rect 17480 54090 17560 54100
rect 17480 54030 17490 54090
rect 17550 54030 17560 54090
rect 17480 54020 17560 54030
rect 15070 53480 16842 53508
rect 15070 53222 16842 53250
rect 14170 52380 14250 52390
rect 14170 52320 14180 52380
rect 14240 52320 14250 52380
rect 14170 52310 14250 52320
rect 14170 50680 14230 52310
rect 15070 51798 16758 53222
rect 16822 51798 16842 53222
rect 17500 52390 17560 54020
rect 17480 52380 17560 52390
rect 17480 52320 17490 52380
rect 17550 52320 17560 52380
rect 17480 52310 17560 52320
rect 15070 51770 16842 51798
rect 15070 51512 16842 51540
rect 14170 50670 14250 50680
rect 14170 50610 14180 50670
rect 14240 50610 14250 50670
rect 14170 50600 14250 50610
rect 14170 48970 14230 50600
rect 15070 50088 16758 51512
rect 16822 50088 16842 51512
rect 17500 50680 17560 52310
rect 17480 50670 17560 50680
rect 17480 50610 17490 50670
rect 17550 50610 17560 50670
rect 17480 50600 17560 50610
rect 15070 50060 16842 50088
rect 15070 49802 16842 49830
rect 14170 48960 14250 48970
rect 14170 48900 14180 48960
rect 14240 48900 14250 48960
rect 14170 48890 14250 48900
rect 14170 47260 14230 48890
rect 15070 48378 16758 49802
rect 16822 48378 16842 49802
rect 17500 48970 17560 50600
rect 17480 48960 17560 48970
rect 17480 48900 17490 48960
rect 17550 48900 17560 48960
rect 17480 48890 17560 48900
rect 15070 48350 16842 48378
rect 15070 48092 16842 48120
rect 14170 47250 14250 47260
rect 14170 47190 14180 47250
rect 14240 47190 14250 47250
rect 14170 47180 14250 47190
rect 15070 46668 16758 48092
rect 16822 46668 16842 48092
rect 17500 47260 17560 48890
rect 17480 47250 17560 47260
rect 17480 47190 17490 47250
rect 17550 47190 17560 47250
rect 17480 47180 17560 47190
rect 15070 46640 16842 46668
rect 15070 46382 16842 46410
rect 14050 45540 14130 45550
rect 12610 45480 12620 45540
rect 12680 45480 12690 45540
rect 12610 45470 12690 45480
rect 10080 44930 11852 44958
rect 10080 44672 11852 44700
rect 9060 43830 9140 43840
rect 7620 43770 7630 43830
rect 7690 43770 7700 43830
rect 7620 43760 7700 43770
rect 5090 43220 6862 43248
rect 5090 42962 6862 42990
rect 4070 42120 4150 42130
rect 2630 42060 2640 42120
rect 2700 42060 2710 42120
rect 2630 42050 2710 42060
rect 100 41510 1872 41538
rect 100 41252 1872 41280
rect 100 39828 1788 41252
rect 1852 39828 1872 41252
rect 2650 40420 2710 42050
rect 4070 42060 4080 42120
rect 4140 42060 4150 42120
rect 4070 42050 4150 42060
rect 2630 40410 2710 40420
rect 3240 40630 3380 40660
rect 3240 40560 3270 40630
rect 3350 40560 3380 40630
rect 3240 40520 3380 40560
rect 3240 40450 3270 40520
rect 3350 40450 3380 40520
rect 3240 40410 3380 40450
rect 4070 40420 4130 42050
rect 5090 41538 6778 42962
rect 6842 41538 6862 42962
rect 7640 42130 7700 43760
rect 9060 43770 9070 43830
rect 9130 43770 9140 43830
rect 9060 43760 9140 43770
rect 7620 42120 7700 42130
rect 8230 42340 8370 42370
rect 8230 42270 8260 42340
rect 8340 42270 8370 42340
rect 8230 42230 8370 42270
rect 8230 42160 8260 42230
rect 8340 42160 8370 42230
rect 8230 42120 8370 42160
rect 9060 42130 9120 43760
rect 10080 43248 11768 44672
rect 11832 43248 11852 44672
rect 12630 43840 12690 45470
rect 14050 45480 14060 45540
rect 14120 45480 14130 45540
rect 14050 45470 14130 45480
rect 12610 43830 12690 43840
rect 13220 44050 13360 44080
rect 13220 43980 13250 44050
rect 13330 43980 13360 44050
rect 13220 43940 13360 43980
rect 13220 43870 13250 43940
rect 13330 43870 13360 43940
rect 13220 43830 13360 43870
rect 14050 43840 14110 45470
rect 15070 44958 16758 46382
rect 16822 44958 16842 46382
rect 17620 45550 17680 60860
rect 19040 60870 19050 60930
rect 19110 60870 19120 60930
rect 19040 60860 19120 60870
rect 18210 59440 18350 59470
rect 18210 59370 18240 59440
rect 18320 59370 18350 59440
rect 18210 59330 18350 59370
rect 18210 59260 18240 59330
rect 18320 59260 18350 59330
rect 18210 59220 18350 59260
rect 18210 57730 18350 57760
rect 18210 57660 18240 57730
rect 18320 57660 18350 57730
rect 18210 57620 18350 57660
rect 18210 57550 18240 57620
rect 18320 57550 18350 57620
rect 18210 57510 18350 57550
rect 18210 56020 18350 56050
rect 18210 55950 18240 56020
rect 18320 55950 18350 56020
rect 18210 55910 18350 55950
rect 18210 55840 18240 55910
rect 18320 55840 18350 55910
rect 18210 55800 18350 55840
rect 18210 54310 18350 54340
rect 18210 54240 18240 54310
rect 18320 54240 18350 54310
rect 18210 54200 18350 54240
rect 18210 54130 18240 54200
rect 18320 54130 18350 54200
rect 18210 54090 18350 54130
rect 18210 52600 18350 52630
rect 18210 52530 18240 52600
rect 18320 52530 18350 52600
rect 18210 52490 18350 52530
rect 18210 52420 18240 52490
rect 18320 52420 18350 52490
rect 18210 52380 18350 52420
rect 18210 50890 18350 50920
rect 18210 50820 18240 50890
rect 18320 50820 18350 50890
rect 18210 50780 18350 50820
rect 18210 50710 18240 50780
rect 18320 50710 18350 50780
rect 18210 50670 18350 50710
rect 18210 49180 18350 49210
rect 18210 49110 18240 49180
rect 18320 49110 18350 49180
rect 18210 49070 18350 49110
rect 18210 49000 18240 49070
rect 18320 49000 18350 49070
rect 18210 48960 18350 49000
rect 18210 47470 18350 47500
rect 18210 47400 18240 47470
rect 18320 47400 18350 47470
rect 18210 47360 18350 47400
rect 18210 47290 18240 47360
rect 18320 47290 18350 47360
rect 18210 47250 18350 47290
rect 17600 45540 17680 45550
rect 18210 45760 18350 45790
rect 18210 45690 18240 45760
rect 18320 45690 18350 45760
rect 18210 45650 18350 45690
rect 18210 45580 18240 45650
rect 18320 45580 18350 45650
rect 18210 45540 18350 45580
rect 19040 45550 19100 60860
rect 20060 60348 21748 61772
rect 21812 60348 21832 61772
rect 22490 60930 22550 62570
rect 22470 60920 22550 60930
rect 22470 60860 22480 60920
rect 22540 60860 22550 60920
rect 22470 60850 22550 60860
rect 20060 60320 21832 60348
rect 20060 60062 21832 60090
rect 19160 59740 19240 59750
rect 19160 59680 19170 59740
rect 19230 59680 19240 59740
rect 19160 59670 19240 59680
rect 19160 59230 19220 59670
rect 19160 59220 19240 59230
rect 19160 59160 19170 59220
rect 19230 59160 19240 59220
rect 19160 59150 19240 59160
rect 19160 57520 19220 59150
rect 20060 58638 21748 60062
rect 21812 58638 21832 60062
rect 22350 59740 22430 59750
rect 22350 59680 22360 59740
rect 22420 59680 22430 59740
rect 22350 59670 22430 59680
rect 22370 59230 22430 59670
rect 22350 59220 22430 59230
rect 22350 59160 22360 59220
rect 22420 59160 22430 59220
rect 22350 59150 22430 59160
rect 20060 58610 21832 58638
rect 20060 58352 21832 58380
rect 19160 57510 19240 57520
rect 19160 57450 19170 57510
rect 19230 57450 19240 57510
rect 19160 57440 19240 57450
rect 19160 55810 19220 57440
rect 20060 56928 21748 58352
rect 21812 56928 21832 58352
rect 22230 58030 22310 58040
rect 22230 57970 22240 58030
rect 22300 57970 22310 58030
rect 22230 57960 22310 57970
rect 22250 57520 22310 57960
rect 22230 57510 22310 57520
rect 22230 57450 22240 57510
rect 22300 57450 22310 57510
rect 22230 57440 22310 57450
rect 20060 56900 21832 56928
rect 20060 56642 21832 56670
rect 19160 55800 19240 55810
rect 19160 55740 19170 55800
rect 19230 55740 19240 55800
rect 19160 55730 19240 55740
rect 19160 54100 19220 55730
rect 20060 55218 21748 56642
rect 21812 55218 21832 56642
rect 22250 55810 22310 57440
rect 22230 55800 22310 55810
rect 22230 55740 22240 55800
rect 22300 55740 22310 55800
rect 22230 55730 22310 55740
rect 20060 55190 21832 55218
rect 20060 54932 21832 54960
rect 19160 54090 19240 54100
rect 19160 54030 19170 54090
rect 19230 54030 19240 54090
rect 19160 54020 19240 54030
rect 19160 52390 19220 54020
rect 20060 53508 21748 54932
rect 21812 53508 21832 54932
rect 22250 54100 22310 55730
rect 22230 54090 22310 54100
rect 22230 54030 22240 54090
rect 22300 54030 22310 54090
rect 22230 54020 22310 54030
rect 20060 53480 21832 53508
rect 20060 53222 21832 53250
rect 19160 52380 19240 52390
rect 19160 52320 19170 52380
rect 19230 52320 19240 52380
rect 19160 52310 19240 52320
rect 19160 50680 19220 52310
rect 20060 51798 21748 53222
rect 21812 51798 21832 53222
rect 22250 52390 22310 54020
rect 22230 52380 22310 52390
rect 22230 52320 22240 52380
rect 22300 52320 22310 52380
rect 22230 52310 22310 52320
rect 20060 51770 21832 51798
rect 20060 51512 21832 51540
rect 19160 50670 19240 50680
rect 19160 50610 19170 50670
rect 19230 50610 19240 50670
rect 19160 50600 19240 50610
rect 19160 48970 19220 50600
rect 20060 50088 21748 51512
rect 21812 50088 21832 51512
rect 22250 50680 22310 52310
rect 22230 50670 22310 50680
rect 22230 50610 22240 50670
rect 22300 50610 22310 50670
rect 22230 50600 22310 50610
rect 20060 50060 21832 50088
rect 20060 49802 21832 49830
rect 19160 48960 19240 48970
rect 19160 48900 19170 48960
rect 19230 48900 19240 48960
rect 19160 48890 19240 48900
rect 19160 47260 19220 48890
rect 20060 48378 21748 49802
rect 21812 48378 21832 49802
rect 22250 48970 22310 50600
rect 22230 48960 22310 48970
rect 22230 48900 22240 48960
rect 22300 48900 22310 48960
rect 22230 48890 22310 48900
rect 20060 48350 21832 48378
rect 20060 48092 21832 48120
rect 19160 47250 19240 47260
rect 19160 47190 19170 47250
rect 19230 47190 19240 47250
rect 19160 47180 19240 47190
rect 20060 46668 21748 48092
rect 21812 46668 21832 48092
rect 22370 47260 22430 59150
rect 22350 47250 22430 47260
rect 22350 47190 22360 47250
rect 22420 47190 22430 47250
rect 22350 47180 22430 47190
rect 20060 46640 21832 46668
rect 20060 46382 21832 46410
rect 19040 45540 19120 45550
rect 17600 45480 17610 45540
rect 17670 45480 17680 45540
rect 17600 45470 17680 45480
rect 15070 44930 16842 44958
rect 15070 44672 16842 44700
rect 14050 43830 14130 43840
rect 12610 43770 12620 43830
rect 12680 43770 12690 43830
rect 12610 43760 12690 43770
rect 10080 43220 11852 43248
rect 10080 42962 11852 42990
rect 9060 42120 9140 42130
rect 7620 42060 7630 42120
rect 7690 42060 7700 42120
rect 7620 42050 7700 42060
rect 5090 41510 6862 41538
rect 5090 41252 6862 41280
rect 4070 40410 4150 40420
rect 2630 40350 2640 40410
rect 2700 40350 2710 40410
rect 2630 40340 2710 40350
rect 4070 40350 4080 40410
rect 4140 40350 4150 40410
rect 4070 40340 4150 40350
rect 100 39800 1872 39828
rect 5090 39828 6778 41252
rect 6842 39828 6862 41252
rect 7640 40420 7700 42050
rect 9060 42060 9070 42120
rect 9130 42060 9140 42120
rect 9060 42050 9140 42060
rect 7620 40410 7700 40420
rect 8230 40630 8370 40660
rect 8230 40560 8260 40630
rect 8340 40560 8370 40630
rect 8230 40520 8370 40560
rect 8230 40450 8260 40520
rect 8340 40450 8370 40520
rect 8230 40410 8370 40450
rect 9060 40420 9120 42050
rect 10080 41538 11768 42962
rect 11832 41538 11852 42962
rect 12630 42130 12690 43760
rect 14050 43770 14060 43830
rect 14120 43770 14130 43830
rect 14050 43760 14130 43770
rect 12610 42120 12690 42130
rect 13220 42340 13360 42370
rect 13220 42270 13250 42340
rect 13330 42270 13360 42340
rect 13220 42230 13360 42270
rect 13220 42160 13250 42230
rect 13330 42160 13360 42230
rect 13220 42120 13360 42160
rect 14050 42130 14110 43760
rect 15070 43248 16758 44672
rect 16822 43248 16842 44672
rect 17620 43840 17680 45470
rect 19040 45480 19050 45540
rect 19110 45480 19120 45540
rect 19040 45470 19120 45480
rect 17600 43830 17680 43840
rect 18210 44050 18350 44080
rect 18210 43980 18240 44050
rect 18320 43980 18350 44050
rect 18210 43940 18350 43980
rect 18210 43870 18240 43940
rect 18320 43870 18350 43940
rect 18210 43830 18350 43870
rect 19040 43840 19100 45470
rect 20060 44958 21748 46382
rect 21812 44958 21832 46382
rect 22490 45550 22550 60850
rect 22470 45540 22550 45550
rect 22470 45480 22480 45540
rect 22540 45480 22550 45540
rect 22470 45470 22550 45480
rect 20060 44930 21832 44958
rect 20060 44672 21832 44700
rect 19040 43830 19120 43840
rect 17600 43770 17610 43830
rect 17670 43770 17680 43830
rect 17600 43760 17680 43770
rect 15070 43220 16842 43248
rect 15070 42962 16842 42990
rect 14050 42120 14130 42130
rect 12610 42060 12620 42120
rect 12680 42060 12690 42120
rect 12610 42050 12690 42060
rect 10080 41510 11852 41538
rect 10080 41252 11852 41280
rect 9060 40410 9140 40420
rect 7620 40350 7630 40410
rect 7690 40350 7700 40410
rect 7620 40340 7700 40350
rect 9060 40350 9070 40410
rect 9130 40350 9140 40410
rect 9060 40340 9140 40350
rect 5090 39800 6862 39828
rect 10080 39828 11768 41252
rect 11832 39828 11852 41252
rect 12630 40420 12690 42050
rect 14050 42060 14060 42120
rect 14120 42060 14130 42120
rect 14050 42050 14130 42060
rect 12610 40410 12690 40420
rect 13220 40630 13360 40660
rect 13220 40560 13250 40630
rect 13330 40560 13360 40630
rect 13220 40520 13360 40560
rect 13220 40450 13250 40520
rect 13330 40450 13360 40520
rect 13220 40410 13360 40450
rect 14050 40420 14110 42050
rect 15070 41538 16758 42962
rect 16822 41538 16842 42962
rect 17620 42130 17680 43760
rect 19040 43770 19050 43830
rect 19110 43770 19120 43830
rect 19040 43760 19120 43770
rect 17600 42120 17680 42130
rect 18210 42340 18350 42370
rect 18210 42270 18240 42340
rect 18320 42270 18350 42340
rect 18210 42230 18350 42270
rect 18210 42160 18240 42230
rect 18320 42160 18350 42230
rect 18210 42120 18350 42160
rect 19040 42130 19100 43760
rect 20060 43248 21748 44672
rect 21812 43248 21832 44672
rect 22490 43840 22550 45470
rect 22470 43830 22550 43840
rect 22470 43770 22480 43830
rect 22540 43770 22550 43830
rect 22470 43760 22550 43770
rect 20060 43220 21832 43248
rect 20060 42962 21832 42990
rect 19040 42120 19120 42130
rect 17600 42060 17610 42120
rect 17670 42060 17680 42120
rect 17600 42050 17680 42060
rect 15070 41510 16842 41538
rect 15070 41252 16842 41280
rect 14050 40410 14130 40420
rect 12610 40350 12620 40410
rect 12680 40350 12690 40410
rect 12610 40340 12690 40350
rect 14050 40350 14060 40410
rect 14120 40350 14130 40410
rect 14050 40340 14130 40350
rect 10080 39800 11852 39828
rect 15070 39828 16758 41252
rect 16822 39828 16842 41252
rect 17620 40420 17680 42050
rect 19040 42060 19050 42120
rect 19110 42060 19120 42120
rect 19040 42050 19120 42060
rect 17600 40410 17680 40420
rect 18210 40630 18350 40660
rect 18210 40560 18240 40630
rect 18320 40560 18350 40630
rect 18210 40520 18350 40560
rect 18210 40450 18240 40520
rect 18320 40450 18350 40520
rect 18210 40410 18350 40450
rect 19040 40420 19100 42050
rect 20060 41538 21748 42962
rect 21812 41538 21832 42962
rect 22610 42130 22670 64280
rect 24030 64290 24040 64350
rect 24100 64290 24110 64350
rect 24030 64280 24110 64290
rect 23200 62860 23340 62890
rect 23200 62790 23230 62860
rect 23310 62790 23340 62860
rect 23200 62750 23340 62790
rect 23200 62680 23230 62750
rect 23310 62680 23340 62750
rect 23200 62640 23340 62680
rect 23200 61150 23340 61180
rect 23200 61080 23230 61150
rect 23310 61080 23340 61150
rect 23200 61040 23340 61080
rect 23200 60970 23230 61040
rect 23310 60970 23340 61040
rect 23200 60930 23340 60970
rect 23200 59440 23340 59470
rect 23200 59370 23230 59440
rect 23310 59370 23340 59440
rect 23200 59330 23340 59370
rect 23200 59260 23230 59330
rect 23310 59260 23340 59330
rect 23200 59220 23340 59260
rect 23200 57730 23340 57760
rect 23200 57660 23230 57730
rect 23310 57660 23340 57730
rect 23200 57620 23340 57660
rect 23200 57550 23230 57620
rect 23310 57550 23340 57620
rect 23200 57510 23340 57550
rect 23200 56020 23340 56050
rect 23200 55950 23230 56020
rect 23310 55950 23340 56020
rect 23200 55910 23340 55950
rect 23200 55840 23230 55910
rect 23310 55840 23340 55910
rect 23200 55800 23340 55840
rect 23200 54310 23340 54340
rect 23200 54240 23230 54310
rect 23310 54240 23340 54310
rect 23200 54200 23340 54240
rect 23200 54130 23230 54200
rect 23310 54130 23340 54200
rect 23200 54090 23340 54130
rect 23200 52600 23340 52630
rect 23200 52530 23230 52600
rect 23310 52530 23340 52600
rect 23200 52490 23340 52530
rect 23200 52420 23230 52490
rect 23310 52420 23340 52490
rect 23200 52380 23340 52420
rect 23200 50890 23340 50920
rect 23200 50820 23230 50890
rect 23310 50820 23340 50890
rect 23200 50780 23340 50820
rect 23200 50710 23230 50780
rect 23310 50710 23340 50780
rect 23200 50670 23340 50710
rect 23200 49180 23340 49210
rect 23200 49110 23230 49180
rect 23310 49110 23340 49180
rect 23200 49070 23340 49110
rect 23200 49000 23230 49070
rect 23310 49000 23340 49070
rect 23200 48960 23340 49000
rect 23200 47470 23340 47500
rect 23200 47400 23230 47470
rect 23310 47400 23340 47470
rect 23200 47360 23340 47400
rect 23200 47290 23230 47360
rect 23310 47290 23340 47360
rect 23200 47250 23340 47290
rect 23200 45760 23340 45790
rect 23200 45690 23230 45760
rect 23310 45690 23340 45760
rect 23200 45650 23340 45690
rect 23200 45580 23230 45650
rect 23310 45580 23340 45650
rect 23200 45540 23340 45580
rect 23200 44050 23340 44080
rect 23200 43980 23230 44050
rect 23310 43980 23340 44050
rect 23200 43940 23340 43980
rect 23200 43870 23230 43940
rect 23310 43870 23340 43940
rect 23200 43830 23340 43870
rect 22590 42120 22670 42130
rect 23200 42340 23340 42370
rect 23200 42270 23230 42340
rect 23310 42270 23340 42340
rect 23200 42230 23340 42270
rect 23200 42160 23230 42230
rect 23310 42160 23340 42230
rect 23200 42120 23340 42160
rect 24030 42130 24090 64280
rect 25050 63768 26738 65192
rect 26802 63768 26822 65192
rect 27600 64360 27660 65990
rect 29020 66000 29030 66060
rect 29090 66000 29100 66060
rect 29020 65990 29100 66000
rect 27580 64350 27660 64360
rect 28190 64570 28330 64600
rect 28190 64500 28220 64570
rect 28300 64500 28330 64570
rect 28190 64460 28330 64500
rect 28190 64390 28220 64460
rect 28300 64390 28330 64460
rect 28190 64350 28330 64390
rect 29020 64360 29080 65990
rect 30040 65478 31728 66902
rect 31792 65478 31812 66902
rect 35030 66902 36802 66930
rect 32570 66580 32650 66590
rect 32570 66520 32580 66580
rect 32640 66520 32650 66580
rect 32570 66510 32650 66520
rect 32590 66070 32650 66510
rect 34010 66580 34090 66590
rect 34010 66520 34020 66580
rect 34080 66520 34090 66580
rect 34010 66510 34090 66520
rect 32570 66060 32650 66070
rect 33180 66280 33320 66310
rect 33180 66210 33210 66280
rect 33290 66210 33320 66280
rect 33180 66170 33320 66210
rect 33180 66100 33210 66170
rect 33290 66100 33320 66170
rect 33180 66060 33320 66100
rect 34010 66070 34070 66510
rect 34010 66060 34090 66070
rect 32570 66000 32580 66060
rect 32640 66000 32650 66060
rect 32570 65990 32650 66000
rect 30040 65450 31812 65478
rect 30040 65192 31812 65220
rect 29020 64350 29100 64360
rect 27580 64290 27590 64350
rect 27650 64290 27660 64350
rect 27580 64280 27660 64290
rect 25050 63740 26822 63768
rect 25050 63482 26822 63510
rect 24150 63160 24230 63170
rect 24150 63100 24160 63160
rect 24220 63100 24230 63160
rect 24150 63090 24230 63100
rect 24150 62650 24210 63090
rect 24150 62640 24230 62650
rect 24150 62580 24160 62640
rect 24220 62580 24230 62640
rect 24150 62570 24230 62580
rect 24150 60930 24210 62570
rect 25050 62058 26738 63482
rect 26802 62058 26822 63482
rect 27460 63160 27540 63170
rect 27460 63100 27470 63160
rect 27530 63100 27540 63160
rect 27460 63090 27540 63100
rect 27480 62650 27540 63090
rect 27460 62640 27540 62650
rect 27460 62580 27470 62640
rect 27530 62580 27540 62640
rect 27460 62570 27540 62580
rect 25050 62030 26822 62058
rect 25050 61772 26822 61800
rect 24150 60920 24230 60930
rect 24150 60860 24160 60920
rect 24220 60860 24230 60920
rect 24150 60850 24230 60860
rect 24150 45550 24210 60850
rect 25050 60348 26738 61772
rect 26802 60348 26822 61772
rect 27480 60930 27540 62570
rect 27460 60920 27540 60930
rect 27460 60860 27470 60920
rect 27530 60860 27540 60920
rect 27460 60850 27540 60860
rect 25050 60320 26822 60348
rect 25050 60062 26822 60090
rect 24270 59740 24350 59750
rect 24270 59680 24280 59740
rect 24340 59680 24350 59740
rect 24270 59670 24350 59680
rect 24270 59230 24330 59670
rect 24270 59220 24350 59230
rect 24270 59160 24280 59220
rect 24340 59160 24350 59220
rect 24270 59150 24350 59160
rect 24270 47260 24330 59150
rect 25050 58638 26738 60062
rect 26802 58638 26822 60062
rect 27340 59740 27420 59750
rect 27340 59680 27350 59740
rect 27410 59680 27420 59740
rect 27340 59670 27420 59680
rect 27360 59230 27420 59670
rect 27340 59220 27420 59230
rect 27340 59160 27350 59220
rect 27410 59160 27420 59220
rect 27340 59150 27420 59160
rect 25050 58610 26822 58638
rect 25050 58352 26822 58380
rect 24390 58030 24470 58040
rect 24390 57970 24400 58030
rect 24460 57970 24470 58030
rect 24390 57960 24470 57970
rect 24390 57520 24450 57960
rect 24390 57510 24470 57520
rect 24390 57450 24400 57510
rect 24460 57450 24470 57510
rect 24390 57440 24470 57450
rect 24390 55810 24450 57440
rect 25050 56928 26738 58352
rect 26802 56928 26822 58352
rect 27220 58030 27300 58040
rect 27220 57970 27230 58030
rect 27290 57970 27300 58030
rect 27220 57960 27300 57970
rect 27240 57520 27300 57960
rect 27220 57510 27300 57520
rect 27220 57450 27230 57510
rect 27290 57450 27300 57510
rect 27220 57440 27300 57450
rect 25050 56900 26822 56928
rect 25050 56642 26822 56670
rect 24390 55800 24470 55810
rect 24390 55740 24400 55800
rect 24460 55740 24470 55800
rect 24390 55730 24470 55740
rect 24390 54100 24450 55730
rect 25050 55218 26738 56642
rect 26802 55218 26822 56642
rect 27240 55810 27300 57440
rect 27220 55800 27300 55810
rect 27220 55740 27230 55800
rect 27290 55740 27300 55800
rect 27220 55730 27300 55740
rect 25050 55190 26822 55218
rect 25050 54932 26822 54960
rect 24390 54090 24470 54100
rect 24390 54030 24400 54090
rect 24460 54030 24470 54090
rect 24390 54020 24470 54030
rect 24390 52390 24450 54020
rect 25050 53508 26738 54932
rect 26802 53508 26822 54932
rect 27240 54100 27300 55730
rect 27220 54090 27300 54100
rect 27220 54030 27230 54090
rect 27290 54030 27300 54090
rect 27220 54020 27300 54030
rect 25050 53480 26822 53508
rect 25050 53222 26822 53250
rect 24390 52380 24470 52390
rect 24390 52320 24400 52380
rect 24460 52320 24470 52380
rect 24390 52310 24470 52320
rect 24390 50680 24450 52310
rect 25050 51798 26738 53222
rect 26802 51798 26822 53222
rect 27240 52390 27300 54020
rect 27220 52380 27300 52390
rect 27220 52320 27230 52380
rect 27290 52320 27300 52380
rect 27220 52310 27300 52320
rect 25050 51770 26822 51798
rect 25050 51512 26822 51540
rect 24390 50670 24470 50680
rect 24390 50610 24400 50670
rect 24460 50610 24470 50670
rect 24390 50600 24470 50610
rect 24390 48970 24450 50600
rect 25050 50088 26738 51512
rect 26802 50088 26822 51512
rect 27240 50680 27300 52310
rect 27220 50670 27300 50680
rect 27220 50610 27230 50670
rect 27290 50610 27300 50670
rect 27220 50600 27300 50610
rect 25050 50060 26822 50088
rect 25050 49802 26822 49830
rect 24390 48960 24470 48970
rect 24390 48900 24400 48960
rect 24460 48900 24470 48960
rect 24390 48890 24470 48900
rect 25050 48378 26738 49802
rect 26802 48378 26822 49802
rect 27240 48970 27300 50600
rect 27220 48960 27300 48970
rect 27220 48900 27230 48960
rect 27290 48900 27300 48960
rect 27220 48890 27300 48900
rect 25050 48350 26822 48378
rect 25050 48092 26822 48120
rect 24270 47250 24350 47260
rect 24270 47190 24280 47250
rect 24340 47190 24350 47250
rect 24270 47180 24350 47190
rect 25050 46668 26738 48092
rect 26802 46668 26822 48092
rect 27360 47260 27420 59150
rect 27340 47250 27420 47260
rect 27340 47190 27350 47250
rect 27410 47190 27420 47250
rect 27340 47180 27420 47190
rect 25050 46640 26822 46668
rect 25050 46382 26822 46410
rect 24150 45540 24230 45550
rect 24150 45480 24160 45540
rect 24220 45480 24230 45540
rect 24150 45470 24230 45480
rect 24150 43840 24210 45470
rect 25050 44958 26738 46382
rect 26802 44958 26822 46382
rect 27480 45550 27540 60850
rect 27460 45540 27540 45550
rect 27460 45480 27470 45540
rect 27530 45480 27540 45540
rect 27460 45470 27540 45480
rect 25050 44930 26822 44958
rect 25050 44672 26822 44700
rect 24150 43830 24230 43840
rect 24150 43770 24160 43830
rect 24220 43770 24230 43830
rect 24150 43760 24230 43770
rect 25050 43248 26738 44672
rect 26802 43248 26822 44672
rect 27480 43840 27540 45470
rect 27460 43830 27540 43840
rect 27460 43770 27470 43830
rect 27530 43770 27540 43830
rect 27460 43760 27540 43770
rect 25050 43220 26822 43248
rect 25050 42962 26822 42990
rect 24030 42120 24110 42130
rect 22590 42060 22600 42120
rect 22660 42060 22670 42120
rect 22590 42050 22670 42060
rect 20060 41510 21832 41538
rect 20060 41252 21832 41280
rect 19040 40410 19120 40420
rect 17600 40350 17610 40410
rect 17670 40350 17680 40410
rect 17600 40340 17680 40350
rect 19040 40350 19050 40410
rect 19110 40350 19120 40410
rect 19040 40340 19120 40350
rect 15070 39800 16842 39828
rect 20060 39828 21748 41252
rect 21812 39828 21832 41252
rect 22610 40420 22670 42050
rect 24030 42060 24040 42120
rect 24100 42060 24110 42120
rect 24030 42050 24110 42060
rect 22590 40410 22670 40420
rect 23200 40630 23340 40660
rect 23200 40560 23230 40630
rect 23310 40560 23340 40630
rect 23200 40520 23340 40560
rect 23200 40450 23230 40520
rect 23310 40450 23340 40520
rect 23200 40410 23340 40450
rect 24030 40420 24090 42050
rect 25050 41538 26738 42962
rect 26802 41538 26822 42962
rect 27600 42130 27660 64280
rect 29020 64290 29030 64350
rect 29090 64290 29100 64350
rect 29020 64280 29100 64290
rect 28190 62860 28330 62890
rect 28190 62790 28220 62860
rect 28300 62790 28330 62860
rect 28190 62750 28330 62790
rect 28190 62680 28220 62750
rect 28300 62680 28330 62750
rect 28190 62640 28330 62680
rect 28190 61150 28330 61180
rect 28190 61080 28220 61150
rect 28300 61080 28330 61150
rect 28190 61040 28330 61080
rect 28190 60970 28220 61040
rect 28300 60970 28330 61040
rect 28190 60930 28330 60970
rect 28190 59440 28330 59470
rect 28190 59370 28220 59440
rect 28300 59370 28330 59440
rect 28190 59330 28330 59370
rect 28190 59260 28220 59330
rect 28300 59260 28330 59330
rect 28190 59220 28330 59260
rect 28190 57730 28330 57760
rect 28190 57660 28220 57730
rect 28300 57660 28330 57730
rect 28190 57620 28330 57660
rect 28190 57550 28220 57620
rect 28300 57550 28330 57620
rect 28190 57510 28330 57550
rect 28190 56020 28330 56050
rect 28190 55950 28220 56020
rect 28300 55950 28330 56020
rect 28190 55910 28330 55950
rect 28190 55840 28220 55910
rect 28300 55840 28330 55910
rect 28190 55800 28330 55840
rect 28190 54310 28330 54340
rect 28190 54240 28220 54310
rect 28300 54240 28330 54310
rect 28190 54200 28330 54240
rect 28190 54130 28220 54200
rect 28300 54130 28330 54200
rect 28190 54090 28330 54130
rect 28190 52600 28330 52630
rect 28190 52530 28220 52600
rect 28300 52530 28330 52600
rect 28190 52490 28330 52530
rect 28190 52420 28220 52490
rect 28300 52420 28330 52490
rect 28190 52380 28330 52420
rect 28190 50890 28330 50920
rect 28190 50820 28220 50890
rect 28300 50820 28330 50890
rect 28190 50780 28330 50820
rect 28190 50710 28220 50780
rect 28300 50710 28330 50780
rect 28190 50670 28330 50710
rect 28190 49180 28330 49210
rect 28190 49110 28220 49180
rect 28300 49110 28330 49180
rect 28190 49070 28330 49110
rect 28190 49000 28220 49070
rect 28300 49000 28330 49070
rect 28190 48960 28330 49000
rect 28190 47470 28330 47500
rect 28190 47400 28220 47470
rect 28300 47400 28330 47470
rect 28190 47360 28330 47400
rect 28190 47290 28220 47360
rect 28300 47290 28330 47360
rect 28190 47250 28330 47290
rect 28190 45760 28330 45790
rect 28190 45690 28220 45760
rect 28300 45690 28330 45760
rect 28190 45650 28330 45690
rect 28190 45580 28220 45650
rect 28300 45580 28330 45650
rect 28190 45540 28330 45580
rect 28190 44050 28330 44080
rect 28190 43980 28220 44050
rect 28300 43980 28330 44050
rect 28190 43940 28330 43980
rect 28190 43870 28220 43940
rect 28300 43870 28330 43940
rect 28190 43830 28330 43870
rect 27580 42120 27660 42130
rect 28190 42340 28330 42370
rect 28190 42270 28220 42340
rect 28300 42270 28330 42340
rect 28190 42230 28330 42270
rect 28190 42160 28220 42230
rect 28300 42160 28330 42230
rect 28190 42120 28330 42160
rect 29020 42130 29080 64280
rect 30040 63768 31728 65192
rect 31792 63768 31812 65192
rect 32590 64360 32650 65990
rect 34010 66000 34020 66060
rect 34080 66000 34090 66060
rect 34010 65990 34090 66000
rect 32570 64350 32650 64360
rect 33180 64570 33320 64600
rect 33180 64500 33210 64570
rect 33290 64500 33320 64570
rect 33180 64460 33320 64500
rect 33180 64390 33210 64460
rect 33290 64390 33320 64460
rect 33180 64350 33320 64390
rect 34010 64360 34070 65990
rect 35030 65478 36718 66902
rect 36782 65478 36802 66902
rect 40020 66902 41792 66930
rect 37560 66590 37640 66600
rect 37560 66530 37570 66590
rect 37630 66530 37640 66590
rect 37560 66520 37640 66530
rect 37580 66080 37640 66520
rect 39000 66590 39080 66600
rect 39000 66530 39010 66590
rect 39070 66530 39080 66590
rect 39000 66520 39080 66530
rect 37560 66070 37640 66080
rect 37560 66010 37570 66070
rect 37630 66010 37640 66070
rect 38170 66280 38310 66310
rect 38170 66210 38200 66280
rect 38280 66210 38310 66280
rect 38170 66170 38310 66210
rect 38170 66100 38200 66170
rect 38280 66100 38310 66170
rect 38170 66060 38310 66100
rect 39000 66080 39060 66520
rect 39000 66070 39080 66080
rect 37560 66000 37640 66010
rect 35030 65450 36802 65478
rect 35030 65192 36802 65220
rect 34010 64350 34090 64360
rect 32570 64290 32580 64350
rect 32640 64290 32650 64350
rect 32570 64280 32650 64290
rect 30040 63740 31812 63768
rect 30040 63482 31812 63510
rect 29140 63160 29220 63170
rect 29140 63100 29150 63160
rect 29210 63100 29220 63160
rect 29140 63090 29220 63100
rect 29140 62650 29200 63090
rect 29140 62640 29220 62650
rect 29140 62580 29150 62640
rect 29210 62580 29220 62640
rect 29140 62570 29220 62580
rect 29140 60930 29200 62570
rect 30040 62058 31728 63482
rect 31792 62058 31812 63482
rect 32450 63160 32530 63170
rect 32450 63100 32460 63160
rect 32520 63100 32530 63160
rect 32450 63090 32530 63100
rect 32470 62650 32530 63090
rect 32450 62640 32530 62650
rect 32450 62580 32460 62640
rect 32520 62580 32530 62640
rect 32450 62570 32530 62580
rect 30040 62030 31812 62058
rect 30040 61772 31812 61800
rect 29140 60920 29220 60930
rect 29140 60860 29150 60920
rect 29210 60860 29220 60920
rect 29140 60850 29220 60860
rect 29140 45550 29200 60850
rect 30040 60348 31728 61772
rect 31792 60348 31812 61772
rect 32470 60940 32530 62570
rect 32450 60930 32530 60940
rect 32450 60870 32460 60930
rect 32520 60870 32530 60930
rect 32450 60860 32530 60870
rect 30040 60320 31812 60348
rect 30040 60062 31812 60090
rect 29260 59740 29340 59750
rect 29260 59680 29270 59740
rect 29330 59680 29340 59740
rect 29260 59670 29340 59680
rect 29260 59230 29320 59670
rect 29260 59220 29340 59230
rect 29260 59160 29270 59220
rect 29330 59160 29340 59220
rect 29260 59150 29340 59160
rect 29260 47260 29320 59150
rect 30040 58638 31728 60062
rect 31792 58638 31812 60062
rect 32330 59740 32410 59750
rect 32330 59680 32340 59740
rect 32400 59680 32410 59740
rect 32330 59670 32410 59680
rect 32350 59230 32410 59670
rect 32330 59220 32410 59230
rect 32330 59160 32340 59220
rect 32400 59160 32410 59220
rect 32330 59150 32410 59160
rect 30040 58610 31812 58638
rect 30040 58352 31812 58380
rect 29380 58030 29460 58040
rect 29380 57970 29390 58030
rect 29450 57970 29460 58030
rect 29380 57960 29460 57970
rect 29380 57520 29440 57960
rect 29380 57510 29460 57520
rect 29380 57450 29390 57510
rect 29450 57450 29460 57510
rect 29380 57440 29460 57450
rect 29380 55810 29440 57440
rect 30040 56928 31728 58352
rect 31792 56928 31812 58352
rect 32210 58030 32290 58040
rect 32210 57970 32220 58030
rect 32280 57970 32290 58030
rect 32210 57960 32290 57970
rect 32230 57520 32290 57960
rect 32210 57510 32290 57520
rect 32210 57450 32220 57510
rect 32280 57450 32290 57510
rect 32210 57440 32290 57450
rect 30040 56900 31812 56928
rect 30040 56642 31812 56670
rect 29380 55800 29460 55810
rect 29380 55740 29390 55800
rect 29450 55740 29460 55800
rect 29380 55730 29460 55740
rect 29380 54100 29440 55730
rect 30040 55218 31728 56642
rect 31792 55218 31812 56642
rect 32090 56320 32170 56330
rect 32090 56260 32100 56320
rect 32160 56260 32170 56320
rect 32090 56250 32170 56260
rect 32110 55810 32170 56250
rect 32090 55800 32170 55810
rect 32090 55740 32100 55800
rect 32160 55740 32170 55800
rect 32090 55730 32170 55740
rect 30040 55190 31812 55218
rect 30040 54932 31812 54960
rect 29380 54090 29460 54100
rect 29380 54030 29390 54090
rect 29450 54030 29460 54090
rect 29380 54020 29460 54030
rect 29380 52390 29440 54020
rect 30040 53508 31728 54932
rect 31792 53508 31812 54932
rect 31970 54610 32050 54620
rect 31970 54550 31980 54610
rect 32040 54550 32050 54610
rect 31970 54540 32050 54550
rect 31990 54100 32050 54540
rect 31970 54090 32050 54100
rect 31970 54030 31980 54090
rect 32040 54030 32050 54090
rect 31970 54020 32050 54030
rect 30040 53480 31812 53508
rect 30040 53222 31812 53250
rect 29380 52380 29460 52390
rect 29380 52320 29390 52380
rect 29450 52320 29460 52380
rect 29380 52310 29460 52320
rect 29380 50680 29440 52310
rect 30040 51798 31728 53222
rect 31792 51798 31812 53222
rect 31990 52390 32050 54020
rect 31970 52380 32050 52390
rect 31970 52320 31980 52380
rect 32040 52320 32050 52380
rect 31970 52310 32050 52320
rect 30040 51770 31812 51798
rect 30040 51512 31812 51540
rect 29380 50670 29460 50680
rect 29380 50610 29390 50670
rect 29450 50610 29460 50670
rect 29380 50600 29460 50610
rect 29380 48970 29440 50600
rect 30040 50088 31728 51512
rect 31792 50088 31812 51512
rect 32110 50680 32170 55730
rect 32090 50670 32170 50680
rect 32090 50610 32100 50670
rect 32160 50610 32170 50670
rect 32090 50600 32170 50610
rect 30040 50060 31812 50088
rect 30040 49802 31812 49830
rect 29380 48960 29460 48970
rect 29380 48900 29390 48960
rect 29450 48900 29460 48960
rect 29380 48890 29460 48900
rect 30040 48378 31728 49802
rect 31792 48378 31812 49802
rect 32230 48970 32290 57440
rect 32210 48960 32290 48970
rect 32210 48900 32220 48960
rect 32280 48900 32290 48960
rect 32210 48890 32290 48900
rect 30040 48350 31812 48378
rect 30040 48092 31812 48120
rect 29260 47250 29340 47260
rect 29260 47190 29270 47250
rect 29330 47190 29340 47250
rect 29260 47180 29340 47190
rect 30040 46668 31728 48092
rect 31792 46668 31812 48092
rect 32350 47260 32410 59150
rect 32330 47250 32410 47260
rect 32330 47190 32340 47250
rect 32400 47190 32410 47250
rect 32330 47180 32410 47190
rect 30040 46640 31812 46668
rect 30040 46382 31812 46410
rect 29140 45540 29220 45550
rect 29140 45480 29150 45540
rect 29210 45480 29220 45540
rect 29140 45470 29220 45480
rect 29140 43840 29200 45470
rect 30040 44958 31728 46382
rect 31792 44958 31812 46382
rect 32470 45550 32530 60860
rect 32450 45540 32530 45550
rect 32450 45480 32460 45540
rect 32520 45480 32530 45540
rect 32450 45470 32530 45480
rect 30040 44930 31812 44958
rect 30040 44672 31812 44700
rect 29140 43830 29220 43840
rect 29140 43770 29150 43830
rect 29210 43770 29220 43830
rect 29140 43760 29220 43770
rect 30040 43248 31728 44672
rect 31792 43248 31812 44672
rect 32470 43840 32530 45470
rect 32450 43830 32530 43840
rect 32450 43770 32460 43830
rect 32520 43770 32530 43830
rect 32450 43760 32530 43770
rect 30040 43220 31812 43248
rect 30040 42962 31812 42990
rect 29020 42120 29100 42130
rect 27580 42060 27590 42120
rect 27650 42060 27660 42120
rect 27580 42050 27660 42060
rect 25050 41510 26822 41538
rect 25050 41252 26822 41280
rect 24030 40410 24110 40420
rect 22590 40350 22600 40410
rect 22660 40350 22670 40410
rect 22590 40340 22670 40350
rect 24030 40350 24040 40410
rect 24100 40350 24110 40410
rect 24030 40340 24110 40350
rect 20060 39800 21832 39828
rect 25050 39828 26738 41252
rect 26802 39828 26822 41252
rect 27600 40420 27660 42050
rect 29020 42060 29030 42120
rect 29090 42060 29100 42120
rect 29020 42050 29100 42060
rect 27580 40410 27660 40420
rect 28190 40630 28330 40660
rect 28190 40560 28220 40630
rect 28300 40560 28330 40630
rect 28190 40520 28330 40560
rect 28190 40450 28220 40520
rect 28300 40450 28330 40520
rect 28190 40410 28330 40450
rect 29020 40420 29080 42050
rect 30040 41538 31728 42962
rect 31792 41538 31812 42962
rect 32590 42130 32650 64280
rect 34010 64290 34020 64350
rect 34080 64290 34090 64350
rect 34010 64280 34090 64290
rect 33180 62860 33320 62890
rect 33180 62790 33210 62860
rect 33290 62790 33320 62860
rect 33180 62750 33320 62790
rect 33180 62680 33210 62750
rect 33290 62680 33320 62750
rect 33180 62640 33320 62680
rect 33180 61150 33320 61180
rect 33180 61080 33210 61150
rect 33290 61080 33320 61150
rect 33180 61040 33320 61080
rect 33180 60970 33210 61040
rect 33290 60970 33320 61040
rect 33180 60930 33320 60970
rect 33180 59440 33320 59470
rect 33180 59370 33210 59440
rect 33290 59370 33320 59440
rect 33180 59330 33320 59370
rect 33180 59260 33210 59330
rect 33290 59260 33320 59330
rect 33180 59220 33320 59260
rect 33180 57730 33320 57760
rect 33180 57660 33210 57730
rect 33290 57660 33320 57730
rect 33180 57620 33320 57660
rect 33180 57550 33210 57620
rect 33290 57550 33320 57620
rect 33180 57510 33320 57550
rect 33180 56020 33320 56050
rect 33180 55950 33210 56020
rect 33290 55950 33320 56020
rect 33180 55910 33320 55950
rect 33180 55840 33210 55910
rect 33290 55840 33320 55910
rect 33180 55800 33320 55840
rect 33180 54310 33320 54340
rect 33180 54240 33210 54310
rect 33290 54240 33320 54310
rect 33180 54200 33320 54240
rect 33180 54130 33210 54200
rect 33290 54130 33320 54200
rect 33180 54090 33320 54130
rect 33180 52600 33320 52630
rect 33180 52530 33210 52600
rect 33290 52530 33320 52600
rect 33180 52490 33320 52530
rect 33180 52420 33210 52490
rect 33290 52420 33320 52490
rect 33180 52380 33320 52420
rect 33180 50890 33320 50920
rect 33180 50820 33210 50890
rect 33290 50820 33320 50890
rect 33180 50780 33320 50820
rect 33180 50710 33210 50780
rect 33290 50710 33320 50780
rect 33180 50670 33320 50710
rect 33180 49180 33320 49210
rect 33180 49110 33210 49180
rect 33290 49110 33320 49180
rect 33180 49070 33320 49110
rect 33180 49000 33210 49070
rect 33290 49000 33320 49070
rect 33180 48960 33320 49000
rect 33180 47470 33320 47500
rect 33180 47400 33210 47470
rect 33290 47400 33320 47470
rect 33180 47360 33320 47400
rect 33180 47290 33210 47360
rect 33290 47290 33320 47360
rect 33180 47250 33320 47290
rect 33180 45760 33320 45790
rect 33180 45690 33210 45760
rect 33290 45690 33320 45760
rect 33180 45650 33320 45690
rect 33180 45580 33210 45650
rect 33290 45580 33320 45650
rect 33180 45540 33320 45580
rect 33180 44050 33320 44080
rect 33180 43980 33210 44050
rect 33290 43980 33320 44050
rect 33180 43940 33320 43980
rect 33180 43870 33210 43940
rect 33290 43870 33320 43940
rect 33180 43830 33320 43870
rect 32570 42120 32650 42130
rect 33180 42340 33320 42370
rect 33180 42270 33210 42340
rect 33290 42270 33320 42340
rect 33180 42230 33320 42270
rect 33180 42160 33210 42230
rect 33290 42160 33320 42230
rect 33180 42120 33320 42160
rect 34010 42130 34070 64280
rect 35030 63768 36718 65192
rect 36782 63768 36802 65192
rect 37580 64370 37640 66000
rect 39000 66010 39010 66070
rect 39070 66010 39080 66070
rect 39000 66000 39080 66010
rect 37560 64360 37640 64370
rect 37560 64300 37570 64360
rect 37630 64300 37640 64360
rect 38170 64570 38310 64600
rect 38170 64500 38200 64570
rect 38280 64500 38310 64570
rect 38170 64460 38310 64500
rect 38170 64390 38200 64460
rect 38280 64390 38310 64460
rect 38170 64350 38310 64390
rect 39000 64370 39060 66000
rect 40020 65478 41708 66902
rect 41772 65478 41792 66902
rect 45010 66902 46782 66930
rect 42550 66590 42630 66600
rect 42550 66530 42560 66590
rect 42620 66530 42630 66590
rect 42550 66520 42630 66530
rect 42570 66080 42630 66520
rect 43990 66590 44070 66600
rect 43990 66530 44000 66590
rect 44060 66530 44070 66590
rect 43990 66520 44070 66530
rect 42550 66070 42630 66080
rect 42550 66010 42560 66070
rect 42620 66010 42630 66070
rect 43160 66280 43300 66310
rect 43160 66210 43190 66280
rect 43270 66210 43300 66280
rect 43160 66170 43300 66210
rect 43160 66100 43190 66170
rect 43270 66100 43300 66170
rect 43160 66060 43300 66100
rect 43990 66080 44050 66520
rect 43990 66070 44070 66080
rect 42550 66000 42630 66010
rect 40020 65450 41792 65478
rect 40020 65192 41792 65220
rect 39000 64360 39080 64370
rect 37560 64290 37640 64300
rect 35030 63740 36802 63768
rect 35030 63482 36802 63510
rect 34130 63160 34210 63170
rect 34130 63100 34140 63160
rect 34200 63100 34210 63160
rect 34130 63090 34210 63100
rect 34130 62650 34190 63090
rect 34130 62640 34210 62650
rect 34130 62580 34140 62640
rect 34200 62580 34210 62640
rect 34130 62570 34210 62580
rect 34130 60940 34190 62570
rect 35030 62058 36718 63482
rect 36782 62058 36802 63482
rect 37440 63170 37520 63180
rect 37440 63110 37450 63170
rect 37510 63110 37520 63170
rect 37440 63100 37520 63110
rect 37460 62660 37520 63100
rect 37440 62650 37520 62660
rect 37440 62590 37450 62650
rect 37510 62590 37520 62650
rect 37440 62580 37520 62590
rect 35030 62030 36802 62058
rect 35030 61772 36802 61800
rect 34130 60930 34210 60940
rect 34130 60870 34140 60930
rect 34200 60870 34210 60930
rect 34130 60860 34210 60870
rect 34130 45550 34190 60860
rect 35030 60348 36718 61772
rect 36782 60348 36802 61772
rect 37460 60950 37520 62580
rect 37440 60940 37520 60950
rect 37440 60880 37450 60940
rect 37510 60880 37520 60940
rect 37440 60870 37520 60880
rect 35030 60320 36802 60348
rect 35030 60062 36802 60090
rect 34250 59740 34330 59750
rect 34250 59680 34260 59740
rect 34320 59680 34330 59740
rect 34250 59670 34330 59680
rect 34250 59230 34310 59670
rect 34250 59220 34330 59230
rect 34250 59160 34260 59220
rect 34320 59160 34330 59220
rect 34250 59150 34330 59160
rect 34250 47260 34310 59150
rect 35030 58638 36718 60062
rect 36782 58638 36802 60062
rect 37320 59750 37400 59760
rect 37320 59690 37330 59750
rect 37390 59690 37400 59750
rect 37320 59680 37400 59690
rect 37340 59240 37400 59680
rect 37320 59230 37400 59240
rect 37320 59170 37330 59230
rect 37390 59170 37400 59230
rect 37320 59160 37400 59170
rect 35030 58610 36802 58638
rect 35030 58352 36802 58380
rect 34370 58030 34450 58040
rect 34370 57970 34380 58030
rect 34440 57970 34450 58030
rect 34370 57960 34450 57970
rect 34370 57520 34430 57960
rect 34370 57510 34450 57520
rect 34370 57450 34380 57510
rect 34440 57450 34450 57510
rect 34370 57440 34450 57450
rect 34370 48970 34430 57440
rect 35030 56928 36718 58352
rect 36782 56928 36802 58352
rect 37200 58040 37280 58050
rect 37200 57980 37210 58040
rect 37270 57980 37280 58040
rect 37200 57970 37280 57980
rect 37220 57530 37280 57970
rect 37200 57520 37280 57530
rect 37200 57460 37210 57520
rect 37270 57460 37280 57520
rect 37200 57450 37280 57460
rect 35030 56900 36802 56928
rect 35030 56642 36802 56670
rect 34490 56320 34570 56330
rect 34490 56260 34500 56320
rect 34560 56260 34570 56320
rect 34490 56250 34570 56260
rect 34490 55810 34550 56250
rect 34490 55800 34570 55810
rect 34490 55740 34500 55800
rect 34560 55740 34570 55800
rect 34490 55730 34570 55740
rect 34490 50680 34550 55730
rect 35030 55218 36718 56642
rect 36782 55218 36802 56642
rect 37080 56330 37160 56340
rect 37080 56270 37090 56330
rect 37150 56270 37160 56330
rect 37080 56260 37160 56270
rect 37100 55820 37160 56260
rect 37080 55810 37160 55820
rect 37080 55750 37090 55810
rect 37150 55750 37160 55810
rect 37080 55740 37160 55750
rect 35030 55190 36802 55218
rect 35030 54932 36802 54960
rect 34610 54610 34690 54620
rect 34610 54550 34620 54610
rect 34680 54550 34690 54610
rect 34610 54540 34690 54550
rect 34610 54100 34670 54540
rect 34610 54090 34690 54100
rect 34610 54030 34620 54090
rect 34680 54030 34690 54090
rect 34610 54020 34690 54030
rect 34610 52390 34670 54020
rect 35030 53508 36718 54932
rect 36782 53508 36802 54932
rect 36960 54610 37040 54620
rect 36960 54550 36970 54610
rect 37030 54550 37040 54610
rect 36960 54540 37040 54550
rect 35030 53480 36802 53508
rect 35030 53222 36802 53250
rect 34610 52380 34690 52390
rect 34610 52320 34620 52380
rect 34680 52320 34690 52380
rect 34610 52310 34690 52320
rect 35030 51798 36718 53222
rect 36782 51798 36802 53222
rect 36980 52400 37040 54540
rect 36960 52390 37040 52400
rect 36960 52330 36970 52390
rect 37030 52330 37040 52390
rect 36960 52320 37040 52330
rect 35030 51770 36802 51798
rect 35030 51512 36802 51540
rect 34490 50670 34570 50680
rect 34490 50610 34500 50670
rect 34560 50610 34570 50670
rect 34490 50600 34570 50610
rect 35030 50088 36718 51512
rect 36782 50088 36802 51512
rect 37100 50690 37160 55740
rect 37080 50680 37160 50690
rect 37080 50620 37090 50680
rect 37150 50620 37160 50680
rect 37080 50610 37160 50620
rect 35030 50060 36802 50088
rect 35030 49802 36802 49830
rect 34370 48960 34450 48970
rect 34370 48900 34380 48960
rect 34440 48900 34450 48960
rect 34370 48890 34450 48900
rect 35030 48378 36718 49802
rect 36782 48378 36802 49802
rect 37220 48980 37280 57450
rect 37200 48970 37280 48980
rect 37200 48910 37210 48970
rect 37270 48910 37280 48970
rect 37200 48900 37280 48910
rect 35030 48350 36802 48378
rect 35030 48092 36802 48120
rect 34250 47250 34330 47260
rect 34250 47190 34260 47250
rect 34320 47190 34330 47250
rect 34250 47180 34330 47190
rect 35030 46668 36718 48092
rect 36782 46668 36802 48092
rect 37340 47270 37400 59160
rect 37320 47260 37400 47270
rect 37320 47200 37330 47260
rect 37390 47200 37400 47260
rect 37320 47190 37400 47200
rect 35030 46640 36802 46668
rect 35030 46382 36802 46410
rect 34130 45540 34210 45550
rect 34130 45480 34140 45540
rect 34200 45480 34210 45540
rect 34130 45470 34210 45480
rect 34130 43840 34190 45470
rect 35030 44958 36718 46382
rect 36782 44958 36802 46382
rect 37460 45560 37520 60870
rect 37440 45550 37520 45560
rect 37440 45490 37450 45550
rect 37510 45490 37520 45550
rect 37440 45480 37520 45490
rect 35030 44930 36802 44958
rect 35030 44672 36802 44700
rect 34130 43830 34210 43840
rect 34130 43770 34140 43830
rect 34200 43770 34210 43830
rect 34130 43760 34210 43770
rect 35030 43248 36718 44672
rect 36782 43248 36802 44672
rect 37460 43850 37520 45480
rect 37440 43840 37520 43850
rect 37440 43780 37450 43840
rect 37510 43780 37520 43840
rect 37440 43770 37520 43780
rect 35030 43220 36802 43248
rect 35030 42962 36802 42990
rect 34010 42120 34090 42130
rect 32570 42060 32580 42120
rect 32640 42060 32650 42120
rect 32570 42050 32650 42060
rect 30040 41510 31812 41538
rect 30040 41252 31812 41280
rect 29020 40410 29100 40420
rect 27580 40350 27590 40410
rect 27650 40350 27660 40410
rect 27580 40340 27660 40350
rect 29020 40350 29030 40410
rect 29090 40350 29100 40410
rect 29020 40340 29100 40350
rect 25050 39800 26822 39828
rect 30040 39828 31728 41252
rect 31792 39828 31812 41252
rect 32590 40420 32650 42050
rect 34010 42060 34020 42120
rect 34080 42060 34090 42120
rect 34010 42050 34090 42060
rect 32570 40410 32650 40420
rect 33180 40630 33320 40660
rect 33180 40560 33210 40630
rect 33290 40560 33320 40630
rect 33180 40520 33320 40560
rect 33180 40450 33210 40520
rect 33290 40450 33320 40520
rect 33180 40410 33320 40450
rect 34010 40420 34070 42050
rect 35030 41538 36718 42962
rect 36782 41538 36802 42962
rect 37580 42140 37640 64290
rect 39000 64300 39010 64360
rect 39070 64300 39080 64360
rect 39000 64290 39080 64300
rect 38170 62860 38310 62890
rect 38170 62790 38200 62860
rect 38280 62790 38310 62860
rect 38170 62750 38310 62790
rect 38170 62680 38200 62750
rect 38280 62680 38310 62750
rect 38170 62640 38310 62680
rect 38170 61150 38310 61180
rect 38170 61080 38200 61150
rect 38280 61080 38310 61150
rect 38170 61040 38310 61080
rect 38170 60970 38200 61040
rect 38280 60970 38310 61040
rect 38170 60930 38310 60970
rect 38170 59440 38310 59470
rect 38170 59370 38200 59440
rect 38280 59370 38310 59440
rect 38170 59330 38310 59370
rect 38170 59260 38200 59330
rect 38280 59260 38310 59330
rect 38170 59220 38310 59260
rect 38170 57730 38310 57760
rect 38170 57660 38200 57730
rect 38280 57660 38310 57730
rect 38170 57620 38310 57660
rect 38170 57550 38200 57620
rect 38280 57550 38310 57620
rect 38170 57510 38310 57550
rect 38170 56020 38310 56050
rect 38170 55950 38200 56020
rect 38280 55950 38310 56020
rect 38170 55910 38310 55950
rect 38170 55840 38200 55910
rect 38280 55840 38310 55910
rect 38170 55800 38310 55840
rect 38170 54310 38310 54340
rect 38170 54240 38200 54310
rect 38280 54240 38310 54310
rect 38170 54200 38310 54240
rect 38170 54130 38200 54200
rect 38280 54130 38310 54200
rect 38170 54090 38310 54130
rect 38170 52600 38310 52630
rect 38170 52530 38200 52600
rect 38280 52530 38310 52600
rect 38170 52490 38310 52530
rect 38170 52420 38200 52490
rect 38280 52420 38310 52490
rect 38170 52380 38310 52420
rect 38170 50890 38310 50920
rect 38170 50820 38200 50890
rect 38280 50820 38310 50890
rect 38170 50780 38310 50820
rect 38170 50710 38200 50780
rect 38280 50710 38310 50780
rect 38170 50670 38310 50710
rect 38170 49180 38310 49210
rect 38170 49110 38200 49180
rect 38280 49110 38310 49180
rect 38170 49070 38310 49110
rect 38170 49000 38200 49070
rect 38280 49000 38310 49070
rect 38170 48960 38310 49000
rect 38170 47470 38310 47500
rect 38170 47400 38200 47470
rect 38280 47400 38310 47470
rect 38170 47360 38310 47400
rect 38170 47290 38200 47360
rect 38280 47290 38310 47360
rect 38170 47250 38310 47290
rect 38170 45760 38310 45790
rect 38170 45690 38200 45760
rect 38280 45690 38310 45760
rect 38170 45650 38310 45690
rect 38170 45580 38200 45650
rect 38280 45580 38310 45650
rect 38170 45540 38310 45580
rect 38170 44050 38310 44080
rect 38170 43980 38200 44050
rect 38280 43980 38310 44050
rect 38170 43940 38310 43980
rect 38170 43870 38200 43940
rect 38280 43870 38310 43940
rect 38170 43830 38310 43870
rect 37560 42130 37640 42140
rect 37560 42070 37570 42130
rect 37630 42070 37640 42130
rect 38170 42340 38310 42370
rect 38170 42270 38200 42340
rect 38280 42270 38310 42340
rect 38170 42230 38310 42270
rect 38170 42160 38200 42230
rect 38280 42160 38310 42230
rect 38170 42120 38310 42160
rect 39000 42130 39060 64290
rect 40020 63768 41708 65192
rect 41772 63768 41792 65192
rect 42570 64370 42630 66000
rect 43990 66010 44000 66070
rect 44060 66010 44070 66070
rect 43990 66000 44070 66010
rect 42550 64360 42630 64370
rect 42550 64300 42560 64360
rect 42620 64300 42630 64360
rect 43160 64570 43300 64600
rect 43160 64500 43190 64570
rect 43270 64500 43300 64570
rect 43160 64460 43300 64500
rect 43160 64390 43190 64460
rect 43270 64390 43300 64460
rect 43160 64350 43300 64390
rect 43990 64370 44050 66000
rect 45010 65478 46698 66902
rect 46762 65478 46782 66902
rect 50000 66902 51772 66930
rect 47540 66580 47620 66590
rect 47540 66520 47550 66580
rect 47610 66520 47620 66580
rect 47540 66510 47620 66520
rect 47560 66070 47620 66510
rect 48980 66580 49060 66590
rect 48980 66520 48990 66580
rect 49050 66520 49060 66580
rect 48980 66510 49060 66520
rect 47540 66060 47620 66070
rect 48150 66280 48290 66310
rect 48150 66210 48180 66280
rect 48260 66210 48290 66280
rect 48150 66170 48290 66210
rect 48150 66100 48180 66170
rect 48260 66100 48290 66170
rect 48150 66060 48290 66100
rect 48980 66070 49040 66510
rect 48980 66060 49060 66070
rect 47540 66000 47550 66060
rect 47610 66000 47620 66060
rect 47540 65990 47620 66000
rect 45010 65450 46782 65478
rect 45010 65192 46782 65220
rect 43990 64360 44070 64370
rect 42550 64290 42630 64300
rect 40020 63740 41792 63768
rect 40020 63482 41792 63510
rect 39120 63170 39200 63180
rect 39120 63110 39130 63170
rect 39190 63110 39200 63170
rect 39120 63100 39200 63110
rect 39120 62660 39180 63100
rect 39120 62650 39200 62660
rect 39120 62590 39130 62650
rect 39190 62590 39200 62650
rect 39120 62580 39200 62590
rect 39120 60950 39180 62580
rect 40020 62058 41708 63482
rect 41772 62058 41792 63482
rect 42430 63170 42510 63180
rect 42430 63110 42440 63170
rect 42500 63110 42510 63170
rect 42430 63100 42510 63110
rect 42450 62660 42510 63100
rect 42430 62650 42510 62660
rect 42430 62590 42440 62650
rect 42500 62590 42510 62650
rect 42430 62580 42510 62590
rect 40020 62030 41792 62058
rect 40020 61772 41792 61800
rect 39120 60940 39200 60950
rect 39120 60880 39130 60940
rect 39190 60880 39200 60940
rect 39120 60870 39200 60880
rect 39120 45560 39180 60870
rect 40020 60348 41708 61772
rect 41772 60348 41792 61772
rect 42450 60950 42510 62580
rect 42430 60940 42510 60950
rect 42430 60880 42440 60940
rect 42500 60880 42510 60940
rect 42430 60870 42510 60880
rect 40020 60320 41792 60348
rect 40020 60062 41792 60090
rect 39240 59750 39320 59760
rect 39240 59690 39250 59750
rect 39310 59690 39320 59750
rect 39240 59680 39320 59690
rect 39240 59240 39300 59680
rect 39240 59230 39320 59240
rect 39240 59170 39250 59230
rect 39310 59170 39320 59230
rect 39240 59160 39320 59170
rect 39240 47270 39300 59160
rect 40020 58638 41708 60062
rect 41772 58638 41792 60062
rect 42310 59750 42390 59760
rect 42310 59690 42320 59750
rect 42380 59690 42390 59750
rect 42310 59680 42390 59690
rect 42330 59240 42390 59680
rect 42310 59230 42390 59240
rect 42310 59170 42320 59230
rect 42380 59170 42390 59230
rect 42310 59160 42390 59170
rect 40020 58610 41792 58638
rect 40020 58352 41792 58380
rect 39360 58040 39440 58050
rect 39360 57980 39370 58040
rect 39430 57980 39440 58040
rect 39360 57970 39440 57980
rect 39360 57530 39420 57970
rect 39360 57520 39440 57530
rect 39360 57460 39370 57520
rect 39430 57460 39440 57520
rect 39360 57450 39440 57460
rect 39360 48980 39420 57450
rect 40020 56928 41708 58352
rect 41772 56928 41792 58352
rect 42190 58040 42270 58050
rect 42190 57980 42200 58040
rect 42260 57980 42270 58040
rect 42190 57970 42270 57980
rect 42210 57530 42270 57970
rect 42190 57520 42270 57530
rect 42190 57460 42200 57520
rect 42260 57460 42270 57520
rect 42190 57450 42270 57460
rect 40020 56900 41792 56928
rect 40020 56642 41792 56670
rect 39480 56330 39560 56340
rect 39480 56270 39490 56330
rect 39550 56270 39560 56330
rect 39480 56260 39560 56270
rect 39480 55820 39540 56260
rect 39480 55810 39560 55820
rect 39480 55750 39490 55810
rect 39550 55750 39560 55810
rect 39480 55740 39560 55750
rect 39480 50690 39540 55740
rect 40020 55218 41708 56642
rect 41772 55218 41792 56642
rect 42070 56330 42150 56340
rect 42070 56270 42080 56330
rect 42140 56270 42150 56330
rect 42070 56260 42150 56270
rect 42090 55820 42150 56260
rect 42070 55810 42150 55820
rect 42070 55750 42080 55810
rect 42140 55750 42150 55810
rect 42070 55740 42150 55750
rect 40020 55190 41792 55218
rect 40020 54932 41792 54960
rect 39600 54660 39680 54670
rect 39600 54600 39610 54660
rect 39670 54600 39680 54660
rect 39600 54590 39680 54600
rect 39600 52400 39660 54590
rect 40020 53508 41708 54932
rect 41772 53508 41792 54932
rect 41950 54610 42030 54620
rect 41950 54550 41960 54610
rect 42020 54550 42030 54610
rect 41950 54540 42030 54550
rect 40020 53480 41792 53508
rect 40020 53222 41792 53250
rect 39600 52390 39680 52400
rect 39600 52330 39610 52390
rect 39670 52330 39680 52390
rect 39600 52320 39680 52330
rect 40020 51798 41708 53222
rect 41772 51798 41792 53222
rect 41970 52400 42030 54540
rect 41950 52390 42030 52400
rect 41950 52330 41960 52390
rect 42020 52330 42030 52390
rect 41950 52320 42030 52330
rect 40020 51770 41792 51798
rect 40020 51512 41792 51540
rect 39480 50680 39560 50690
rect 39480 50620 39490 50680
rect 39550 50620 39560 50680
rect 39480 50610 39560 50620
rect 40020 50088 41708 51512
rect 41772 50088 41792 51512
rect 42090 50690 42150 55740
rect 42070 50680 42150 50690
rect 42070 50620 42080 50680
rect 42140 50620 42150 50680
rect 42070 50610 42150 50620
rect 40020 50060 41792 50088
rect 40020 49802 41792 49830
rect 39360 48970 39440 48980
rect 39360 48910 39370 48970
rect 39430 48910 39440 48970
rect 39360 48900 39440 48910
rect 40020 48378 41708 49802
rect 41772 48378 41792 49802
rect 42210 48980 42270 57450
rect 42190 48970 42270 48980
rect 42190 48910 42200 48970
rect 42260 48910 42270 48970
rect 42190 48900 42270 48910
rect 40020 48350 41792 48378
rect 40020 48092 41792 48120
rect 39240 47260 39320 47270
rect 39240 47200 39250 47260
rect 39310 47200 39320 47260
rect 39240 47190 39320 47200
rect 40020 46668 41708 48092
rect 41772 46668 41792 48092
rect 42330 47270 42390 59160
rect 42310 47260 42390 47270
rect 42310 47200 42320 47260
rect 42380 47200 42390 47260
rect 42310 47190 42390 47200
rect 40020 46640 41792 46668
rect 40020 46382 41792 46410
rect 39120 45550 39200 45560
rect 39120 45490 39130 45550
rect 39190 45490 39200 45550
rect 39120 45480 39200 45490
rect 39120 43840 39180 45480
rect 40020 44958 41708 46382
rect 41772 44958 41792 46382
rect 42450 45560 42510 60870
rect 42430 45550 42510 45560
rect 42430 45490 42440 45550
rect 42500 45490 42510 45550
rect 42430 45480 42510 45490
rect 40020 44930 41792 44958
rect 40020 44672 41792 44700
rect 39120 43830 39200 43840
rect 39120 43770 39130 43830
rect 39190 43770 39200 43830
rect 39120 43760 39200 43770
rect 40020 43248 41708 44672
rect 41772 43248 41792 44672
rect 42450 43850 42510 45480
rect 42430 43840 42510 43850
rect 42430 43780 42440 43840
rect 42500 43780 42510 43840
rect 42430 43770 42510 43780
rect 40020 43220 41792 43248
rect 40020 42962 41792 42990
rect 39000 42120 39080 42130
rect 37560 42060 37640 42070
rect 35030 41510 36802 41538
rect 35030 41252 36802 41280
rect 34010 40410 34090 40420
rect 32570 40350 32580 40410
rect 32640 40350 32650 40410
rect 32570 40340 32650 40350
rect 34010 40350 34020 40410
rect 34080 40350 34090 40410
rect 34010 40340 34090 40350
rect 30040 39800 31812 39828
rect 35030 39828 36718 41252
rect 36782 39828 36802 41252
rect 37580 40430 37640 42060
rect 39000 42060 39010 42120
rect 39070 42060 39080 42120
rect 39000 42050 39080 42060
rect 37560 40420 37640 40430
rect 37560 40360 37570 40420
rect 37630 40360 37640 40420
rect 38170 40630 38310 40660
rect 38170 40560 38200 40630
rect 38280 40560 38310 40630
rect 38170 40520 38310 40560
rect 38170 40450 38200 40520
rect 38280 40450 38310 40520
rect 38170 40410 38310 40450
rect 39000 40430 39060 42050
rect 40020 41538 41708 42962
rect 41772 41538 41792 42962
rect 42570 42140 42630 64290
rect 43990 64300 44000 64360
rect 44060 64300 44070 64360
rect 43990 64290 44070 64300
rect 43160 62860 43300 62890
rect 43160 62790 43190 62860
rect 43270 62790 43300 62860
rect 43160 62750 43300 62790
rect 43160 62680 43190 62750
rect 43270 62680 43300 62750
rect 43160 62640 43300 62680
rect 43160 61150 43300 61180
rect 43160 61080 43190 61150
rect 43270 61080 43300 61150
rect 43160 61040 43300 61080
rect 43160 60970 43190 61040
rect 43270 60970 43300 61040
rect 43160 60930 43300 60970
rect 43160 59440 43300 59470
rect 43160 59370 43190 59440
rect 43270 59370 43300 59440
rect 43160 59330 43300 59370
rect 43160 59260 43190 59330
rect 43270 59260 43300 59330
rect 43160 59220 43300 59260
rect 43160 57730 43300 57760
rect 43160 57660 43190 57730
rect 43270 57660 43300 57730
rect 43160 57620 43300 57660
rect 43160 57550 43190 57620
rect 43270 57550 43300 57620
rect 43160 57510 43300 57550
rect 43160 56020 43300 56050
rect 43160 55950 43190 56020
rect 43270 55950 43300 56020
rect 43160 55910 43300 55950
rect 43160 55840 43190 55910
rect 43270 55840 43300 55910
rect 43160 55800 43300 55840
rect 43160 54310 43300 54340
rect 43160 54240 43190 54310
rect 43270 54240 43300 54310
rect 43160 54200 43300 54240
rect 43160 54130 43190 54200
rect 43270 54130 43300 54200
rect 43160 54090 43300 54130
rect 43160 52600 43300 52630
rect 43160 52530 43190 52600
rect 43270 52530 43300 52600
rect 43160 52490 43300 52530
rect 43160 52420 43190 52490
rect 43270 52420 43300 52490
rect 43160 52380 43300 52420
rect 43160 50890 43300 50920
rect 43160 50820 43190 50890
rect 43270 50820 43300 50890
rect 43160 50780 43300 50820
rect 43160 50710 43190 50780
rect 43270 50710 43300 50780
rect 43160 50670 43300 50710
rect 43160 49180 43300 49210
rect 43160 49110 43190 49180
rect 43270 49110 43300 49180
rect 43160 49070 43300 49110
rect 43160 49000 43190 49070
rect 43270 49000 43300 49070
rect 43160 48960 43300 49000
rect 43160 47470 43300 47500
rect 43160 47400 43190 47470
rect 43270 47400 43300 47470
rect 43160 47360 43300 47400
rect 43160 47290 43190 47360
rect 43270 47290 43300 47360
rect 43160 47250 43300 47290
rect 43160 45760 43300 45790
rect 43160 45690 43190 45760
rect 43270 45690 43300 45760
rect 43160 45650 43300 45690
rect 43160 45580 43190 45650
rect 43270 45580 43300 45650
rect 43160 45540 43300 45580
rect 43160 44050 43300 44080
rect 43160 43980 43190 44050
rect 43270 43980 43300 44050
rect 43160 43940 43300 43980
rect 43160 43870 43190 43940
rect 43270 43870 43300 43940
rect 43160 43830 43300 43870
rect 42550 42130 42630 42140
rect 42550 42070 42560 42130
rect 42620 42070 42630 42130
rect 43160 42340 43300 42370
rect 43160 42270 43190 42340
rect 43270 42270 43300 42340
rect 43160 42230 43300 42270
rect 43160 42160 43190 42230
rect 43270 42160 43300 42230
rect 43160 42120 43300 42160
rect 43990 42130 44050 64290
rect 45010 63768 46698 65192
rect 46762 63768 46782 65192
rect 47560 64360 47620 65990
rect 48980 66000 48990 66060
rect 49050 66000 49060 66060
rect 48980 65990 49060 66000
rect 47540 64350 47620 64360
rect 48150 64570 48290 64600
rect 48150 64500 48180 64570
rect 48260 64500 48290 64570
rect 48150 64460 48290 64500
rect 48150 64390 48180 64460
rect 48260 64390 48290 64460
rect 48150 64350 48290 64390
rect 48980 64360 49040 65990
rect 50000 65478 51688 66902
rect 51752 65478 51772 66902
rect 54990 66902 56762 66930
rect 52530 66580 52610 66590
rect 52530 66520 52540 66580
rect 52600 66520 52610 66580
rect 52530 66510 52610 66520
rect 52550 66070 52610 66510
rect 53970 66580 54050 66590
rect 53970 66520 53980 66580
rect 54040 66520 54050 66580
rect 53970 66510 54050 66520
rect 52530 66060 52610 66070
rect 53140 66280 53280 66310
rect 53140 66210 53170 66280
rect 53250 66210 53280 66280
rect 53140 66170 53280 66210
rect 53140 66100 53170 66170
rect 53250 66100 53280 66170
rect 53140 66060 53280 66100
rect 53970 66070 54030 66510
rect 53970 66060 54050 66070
rect 52530 66000 52540 66060
rect 52600 66000 52610 66060
rect 52530 65990 52610 66000
rect 50000 65450 51772 65478
rect 50000 65192 51772 65220
rect 48980 64350 49060 64360
rect 47540 64290 47550 64350
rect 47610 64290 47620 64350
rect 47540 64280 47620 64290
rect 45010 63740 46782 63768
rect 45010 63482 46782 63510
rect 44110 63170 44190 63180
rect 44110 63110 44120 63170
rect 44180 63110 44190 63170
rect 44110 63100 44190 63110
rect 44110 62660 44170 63100
rect 44110 62650 44190 62660
rect 44110 62590 44120 62650
rect 44180 62590 44190 62650
rect 44110 62580 44190 62590
rect 44110 60950 44170 62580
rect 45010 62058 46698 63482
rect 46762 62058 46782 63482
rect 47420 63160 47500 63170
rect 47420 63100 47430 63160
rect 47490 63100 47500 63160
rect 47420 63090 47500 63100
rect 47440 62650 47500 63090
rect 47420 62640 47500 62650
rect 47420 62580 47430 62640
rect 47490 62580 47500 62640
rect 47420 62570 47500 62580
rect 45010 62030 46782 62058
rect 45010 61772 46782 61800
rect 44110 60940 44190 60950
rect 44110 60880 44120 60940
rect 44180 60880 44190 60940
rect 44110 60870 44190 60880
rect 44110 45560 44170 60870
rect 45010 60348 46698 61772
rect 46762 60348 46782 61772
rect 47440 60940 47500 62570
rect 47420 60930 47500 60940
rect 47420 60870 47430 60930
rect 47490 60870 47500 60930
rect 47420 60860 47500 60870
rect 45010 60320 46782 60348
rect 45010 60062 46782 60090
rect 44230 59750 44310 59760
rect 44230 59690 44240 59750
rect 44300 59690 44310 59750
rect 44230 59680 44310 59690
rect 44230 59240 44290 59680
rect 44230 59230 44310 59240
rect 44230 59170 44240 59230
rect 44300 59170 44310 59230
rect 44230 59160 44310 59170
rect 44230 47270 44290 59160
rect 45010 58638 46698 60062
rect 46762 58638 46782 60062
rect 47300 59740 47380 59750
rect 47300 59680 47310 59740
rect 47370 59680 47380 59740
rect 47300 59670 47380 59680
rect 47320 59230 47380 59670
rect 47300 59220 47380 59230
rect 47300 59160 47310 59220
rect 47370 59160 47380 59220
rect 47300 59150 47380 59160
rect 45010 58610 46782 58638
rect 45010 58352 46782 58380
rect 44350 58040 44430 58050
rect 44350 57980 44360 58040
rect 44420 57980 44430 58040
rect 44350 57970 44430 57980
rect 44350 57530 44410 57970
rect 44350 57520 44430 57530
rect 44350 57460 44360 57520
rect 44420 57460 44430 57520
rect 44350 57450 44430 57460
rect 44350 48980 44410 57450
rect 45010 56928 46698 58352
rect 46762 56928 46782 58352
rect 47180 58030 47260 58040
rect 47180 57970 47190 58030
rect 47250 57970 47260 58030
rect 47180 57960 47260 57970
rect 47200 57520 47260 57960
rect 47180 57510 47260 57520
rect 47180 57450 47190 57510
rect 47250 57450 47260 57510
rect 47180 57440 47260 57450
rect 45010 56900 46782 56928
rect 45010 56642 46782 56670
rect 44470 56330 44550 56340
rect 44470 56270 44480 56330
rect 44540 56270 44550 56330
rect 44470 56260 44550 56270
rect 44470 55820 44530 56260
rect 44470 55810 44550 55820
rect 44470 55750 44480 55810
rect 44540 55750 44550 55810
rect 44470 55740 44550 55750
rect 44470 50690 44530 55740
rect 45010 55218 46698 56642
rect 46762 55218 46782 56642
rect 47060 56320 47140 56330
rect 47060 56260 47070 56320
rect 47130 56260 47140 56320
rect 47060 56250 47140 56260
rect 47080 55810 47140 56250
rect 47060 55800 47140 55810
rect 47060 55740 47070 55800
rect 47130 55740 47140 55800
rect 47060 55730 47140 55740
rect 45010 55190 46782 55218
rect 45010 54932 46782 54960
rect 44590 54660 44670 54670
rect 44590 54600 44600 54660
rect 44660 54600 44670 54660
rect 44590 54590 44670 54600
rect 44590 52400 44650 54590
rect 45010 53508 46698 54932
rect 46762 53508 46782 54932
rect 46940 54610 47020 54620
rect 46940 54550 46950 54610
rect 47010 54550 47020 54610
rect 46940 54540 47020 54550
rect 46960 54100 47020 54540
rect 46940 54090 47020 54100
rect 46940 54030 46950 54090
rect 47010 54030 47020 54090
rect 46940 54020 47020 54030
rect 45010 53480 46782 53508
rect 45010 53222 46782 53250
rect 44590 52390 44670 52400
rect 44590 52330 44600 52390
rect 44660 52330 44670 52390
rect 44590 52320 44670 52330
rect 45010 51798 46698 53222
rect 46762 51798 46782 53222
rect 46960 52390 47020 54020
rect 46940 52380 47020 52390
rect 46940 52320 46950 52380
rect 47010 52320 47020 52380
rect 46940 52310 47020 52320
rect 45010 51770 46782 51798
rect 45010 51512 46782 51540
rect 44470 50680 44550 50690
rect 44470 50620 44480 50680
rect 44540 50620 44550 50680
rect 44470 50610 44550 50620
rect 45010 50088 46698 51512
rect 46762 50088 46782 51512
rect 47080 50680 47140 55730
rect 47060 50670 47140 50680
rect 47060 50610 47070 50670
rect 47130 50610 47140 50670
rect 47060 50600 47140 50610
rect 45010 50060 46782 50088
rect 45010 49802 46782 49830
rect 44350 48970 44430 48980
rect 44350 48910 44360 48970
rect 44420 48910 44430 48970
rect 44350 48900 44430 48910
rect 45010 48378 46698 49802
rect 46762 48378 46782 49802
rect 47200 48970 47260 57440
rect 47180 48960 47260 48970
rect 47180 48900 47190 48960
rect 47250 48900 47260 48960
rect 47180 48890 47260 48900
rect 45010 48350 46782 48378
rect 45010 48092 46782 48120
rect 44230 47260 44310 47270
rect 44230 47200 44240 47260
rect 44300 47200 44310 47260
rect 44230 47190 44310 47200
rect 45010 46668 46698 48092
rect 46762 46668 46782 48092
rect 47320 47260 47380 59150
rect 47300 47250 47380 47260
rect 47300 47190 47310 47250
rect 47370 47190 47380 47250
rect 47300 47180 47380 47190
rect 45010 46640 46782 46668
rect 45010 46382 46782 46410
rect 44110 45550 44190 45560
rect 44110 45490 44120 45550
rect 44180 45490 44190 45550
rect 44110 45480 44190 45490
rect 44110 43840 44170 45480
rect 45010 44958 46698 46382
rect 46762 44958 46782 46382
rect 47440 45550 47500 60860
rect 47420 45540 47500 45550
rect 47420 45480 47430 45540
rect 47490 45480 47500 45540
rect 47420 45470 47500 45480
rect 45010 44930 46782 44958
rect 45010 44672 46782 44700
rect 44110 43830 44190 43840
rect 44110 43770 44120 43830
rect 44180 43770 44190 43830
rect 44110 43760 44190 43770
rect 45010 43248 46698 44672
rect 46762 43248 46782 44672
rect 47440 43840 47500 45470
rect 47420 43830 47500 43840
rect 47420 43770 47430 43830
rect 47490 43770 47500 43830
rect 47420 43760 47500 43770
rect 45010 43220 46782 43248
rect 45010 42962 46782 42990
rect 43990 42120 44070 42130
rect 42550 42060 42630 42070
rect 40020 41510 41792 41538
rect 40020 41252 41792 41280
rect 39000 40420 39080 40430
rect 37560 40350 37640 40360
rect 39000 40360 39010 40420
rect 39070 40360 39080 40420
rect 39000 40350 39080 40360
rect 39000 40220 39060 40350
rect 39000 40210 39080 40220
rect 39000 40150 39010 40210
rect 39070 40150 39080 40210
rect 39000 40140 39080 40150
rect 35030 39800 36802 39828
rect 40020 39828 41708 41252
rect 41772 39828 41792 41252
rect 42570 40430 42630 42060
rect 43990 42060 44000 42120
rect 44060 42060 44070 42120
rect 43990 42050 44070 42060
rect 42550 40420 42630 40430
rect 42550 40360 42560 40420
rect 42620 40360 42630 40420
rect 43160 40630 43300 40660
rect 43160 40560 43190 40630
rect 43270 40560 43300 40630
rect 43160 40520 43300 40560
rect 43160 40450 43190 40520
rect 43270 40450 43300 40520
rect 43160 40410 43300 40450
rect 43990 40430 44050 42050
rect 45010 41538 46698 42962
rect 46762 41538 46782 42962
rect 47560 42130 47620 64280
rect 48980 64290 48990 64350
rect 49050 64290 49060 64350
rect 48980 64280 49060 64290
rect 48150 62860 48290 62890
rect 48150 62790 48180 62860
rect 48260 62790 48290 62860
rect 48150 62750 48290 62790
rect 48150 62680 48180 62750
rect 48260 62680 48290 62750
rect 48150 62640 48290 62680
rect 48150 61150 48290 61180
rect 48150 61080 48180 61150
rect 48260 61080 48290 61150
rect 48150 61040 48290 61080
rect 48150 60970 48180 61040
rect 48260 60970 48290 61040
rect 48150 60930 48290 60970
rect 48150 59440 48290 59470
rect 48150 59370 48180 59440
rect 48260 59370 48290 59440
rect 48150 59330 48290 59370
rect 48150 59260 48180 59330
rect 48260 59260 48290 59330
rect 48150 59220 48290 59260
rect 48150 57730 48290 57760
rect 48150 57660 48180 57730
rect 48260 57660 48290 57730
rect 48150 57620 48290 57660
rect 48150 57550 48180 57620
rect 48260 57550 48290 57620
rect 48150 57510 48290 57550
rect 48150 56020 48290 56050
rect 48150 55950 48180 56020
rect 48260 55950 48290 56020
rect 48150 55910 48290 55950
rect 48150 55840 48180 55910
rect 48260 55840 48290 55910
rect 48150 55800 48290 55840
rect 48150 54310 48290 54340
rect 48150 54240 48180 54310
rect 48260 54240 48290 54310
rect 48150 54200 48290 54240
rect 48150 54130 48180 54200
rect 48260 54130 48290 54200
rect 48150 54090 48290 54130
rect 48150 52600 48290 52630
rect 48150 52530 48180 52600
rect 48260 52530 48290 52600
rect 48150 52490 48290 52530
rect 48150 52420 48180 52490
rect 48260 52420 48290 52490
rect 48150 52380 48290 52420
rect 48150 50890 48290 50920
rect 48150 50820 48180 50890
rect 48260 50820 48290 50890
rect 48150 50780 48290 50820
rect 48150 50710 48180 50780
rect 48260 50710 48290 50780
rect 48150 50670 48290 50710
rect 48150 49180 48290 49210
rect 48150 49110 48180 49180
rect 48260 49110 48290 49180
rect 48150 49070 48290 49110
rect 48150 49000 48180 49070
rect 48260 49000 48290 49070
rect 48150 48960 48290 49000
rect 48150 47470 48290 47500
rect 48150 47400 48180 47470
rect 48260 47400 48290 47470
rect 48150 47360 48290 47400
rect 48150 47290 48180 47360
rect 48260 47290 48290 47360
rect 48150 47250 48290 47290
rect 48150 45760 48290 45790
rect 48150 45690 48180 45760
rect 48260 45690 48290 45760
rect 48150 45650 48290 45690
rect 48150 45580 48180 45650
rect 48260 45580 48290 45650
rect 48150 45540 48290 45580
rect 48150 44050 48290 44080
rect 48150 43980 48180 44050
rect 48260 43980 48290 44050
rect 48150 43940 48290 43980
rect 48150 43870 48180 43940
rect 48260 43870 48290 43940
rect 48150 43830 48290 43870
rect 47540 42120 47620 42130
rect 48150 42340 48290 42370
rect 48150 42270 48180 42340
rect 48260 42270 48290 42340
rect 48150 42230 48290 42270
rect 48150 42160 48180 42230
rect 48260 42160 48290 42230
rect 48150 42120 48290 42160
rect 48980 42130 49040 64280
rect 50000 63768 51688 65192
rect 51752 63768 51772 65192
rect 52550 64360 52610 65990
rect 53970 66000 53980 66060
rect 54040 66000 54050 66060
rect 53970 65990 54050 66000
rect 52530 64350 52610 64360
rect 53140 64570 53280 64600
rect 53140 64500 53170 64570
rect 53250 64500 53280 64570
rect 53140 64460 53280 64500
rect 53140 64390 53170 64460
rect 53250 64390 53280 64460
rect 53140 64350 53280 64390
rect 53970 64360 54030 65990
rect 54990 65478 56678 66902
rect 56742 65478 56762 66902
rect 59980 66902 61752 66930
rect 57520 66580 57600 66590
rect 57520 66520 57530 66580
rect 57590 66520 57600 66580
rect 57520 66510 57600 66520
rect 57540 66070 57600 66510
rect 58960 66580 59040 66590
rect 58960 66520 58970 66580
rect 59030 66520 59040 66580
rect 58960 66510 59040 66520
rect 57520 66060 57600 66070
rect 58130 66280 58270 66310
rect 58130 66210 58160 66280
rect 58240 66210 58270 66280
rect 58130 66170 58270 66210
rect 58130 66100 58160 66170
rect 58240 66100 58270 66170
rect 58130 66060 58270 66100
rect 58960 66070 59020 66510
rect 58960 66060 59040 66070
rect 57520 66000 57530 66060
rect 57590 66000 57600 66060
rect 57520 65990 57600 66000
rect 54990 65450 56762 65478
rect 54990 65192 56762 65220
rect 53970 64350 54050 64360
rect 52530 64290 52540 64350
rect 52600 64290 52610 64350
rect 52530 64280 52610 64290
rect 50000 63740 51772 63768
rect 50000 63482 51772 63510
rect 49100 63160 49180 63170
rect 49100 63100 49110 63160
rect 49170 63100 49180 63160
rect 49100 63090 49180 63100
rect 49100 62650 49160 63090
rect 49100 62640 49180 62650
rect 49100 62580 49110 62640
rect 49170 62580 49180 62640
rect 49100 62570 49180 62580
rect 49100 60940 49160 62570
rect 50000 62058 51688 63482
rect 51752 62058 51772 63482
rect 52410 63160 52490 63170
rect 52410 63100 52420 63160
rect 52480 63100 52490 63160
rect 52410 63090 52490 63100
rect 52430 62650 52490 63090
rect 52410 62640 52490 62650
rect 52410 62580 52420 62640
rect 52480 62580 52490 62640
rect 52410 62570 52490 62580
rect 50000 62030 51772 62058
rect 50000 61772 51772 61800
rect 49100 60930 49180 60940
rect 49100 60870 49110 60930
rect 49170 60870 49180 60930
rect 49100 60860 49180 60870
rect 49100 45550 49160 60860
rect 50000 60348 51688 61772
rect 51752 60348 51772 61772
rect 52430 60930 52490 62570
rect 52410 60920 52490 60930
rect 52410 60860 52420 60920
rect 52480 60860 52490 60920
rect 52410 60850 52490 60860
rect 50000 60320 51772 60348
rect 50000 60062 51772 60090
rect 49220 59740 49300 59750
rect 49220 59680 49230 59740
rect 49290 59680 49300 59740
rect 49220 59670 49300 59680
rect 49220 59230 49280 59670
rect 49220 59220 49300 59230
rect 49220 59160 49230 59220
rect 49290 59160 49300 59220
rect 49220 59150 49300 59160
rect 49220 47260 49280 59150
rect 50000 58638 51688 60062
rect 51752 58638 51772 60062
rect 52290 59740 52370 59750
rect 52290 59680 52300 59740
rect 52360 59680 52370 59740
rect 52290 59670 52370 59680
rect 52310 59230 52370 59670
rect 52290 59220 52370 59230
rect 52290 59160 52300 59220
rect 52360 59160 52370 59220
rect 52290 59150 52370 59160
rect 50000 58610 51772 58638
rect 50000 58352 51772 58380
rect 49340 58030 49420 58040
rect 49340 57970 49350 58030
rect 49410 57970 49420 58030
rect 49340 57960 49420 57970
rect 49340 57520 49400 57960
rect 49340 57510 49420 57520
rect 49340 57450 49350 57510
rect 49410 57450 49420 57510
rect 49340 57440 49420 57450
rect 49340 48970 49400 57440
rect 50000 56928 51688 58352
rect 51752 56928 51772 58352
rect 52170 58030 52250 58040
rect 52170 57970 52180 58030
rect 52240 57970 52250 58030
rect 52170 57960 52250 57970
rect 52190 57520 52250 57960
rect 52170 57510 52250 57520
rect 52170 57450 52180 57510
rect 52240 57450 52250 57510
rect 52170 57440 52250 57450
rect 50000 56900 51772 56928
rect 50000 56642 51772 56670
rect 49460 56320 49540 56330
rect 49460 56260 49470 56320
rect 49530 56260 49540 56320
rect 49460 56250 49540 56260
rect 49460 55810 49520 56250
rect 49460 55800 49540 55810
rect 49460 55740 49470 55800
rect 49530 55740 49540 55800
rect 49460 55730 49540 55740
rect 49460 50680 49520 55730
rect 50000 55218 51688 56642
rect 51752 55218 51772 56642
rect 52190 55810 52250 57440
rect 52170 55800 52250 55810
rect 52170 55740 52180 55800
rect 52240 55740 52250 55800
rect 52170 55730 52250 55740
rect 50000 55190 51772 55218
rect 50000 54932 51772 54960
rect 49580 54610 49660 54620
rect 49580 54550 49590 54610
rect 49650 54550 49660 54610
rect 49580 54540 49660 54550
rect 49580 54100 49640 54540
rect 49580 54090 49660 54100
rect 49580 54030 49590 54090
rect 49650 54030 49660 54090
rect 49580 54020 49660 54030
rect 49580 52390 49640 54020
rect 50000 53508 51688 54932
rect 51752 53508 51772 54932
rect 52190 54100 52250 55730
rect 52170 54090 52250 54100
rect 52170 54030 52180 54090
rect 52240 54030 52250 54090
rect 52170 54020 52250 54030
rect 50000 53480 51772 53508
rect 50000 53222 51772 53250
rect 49580 52380 49660 52390
rect 49580 52320 49590 52380
rect 49650 52320 49660 52380
rect 49580 52310 49660 52320
rect 50000 51798 51688 53222
rect 51752 51798 51772 53222
rect 52190 52390 52250 54020
rect 52170 52380 52250 52390
rect 52170 52320 52180 52380
rect 52240 52320 52250 52380
rect 52170 52310 52250 52320
rect 50000 51770 51772 51798
rect 50000 51512 51772 51540
rect 49460 50670 49540 50680
rect 49460 50610 49470 50670
rect 49530 50610 49540 50670
rect 49460 50600 49540 50610
rect 50000 50088 51688 51512
rect 51752 50088 51772 51512
rect 52190 50680 52250 52310
rect 52170 50670 52250 50680
rect 52170 50610 52180 50670
rect 52240 50610 52250 50670
rect 52170 50600 52250 50610
rect 50000 50060 51772 50088
rect 50000 49802 51772 49830
rect 49340 48960 49420 48970
rect 49340 48900 49350 48960
rect 49410 48900 49420 48960
rect 49340 48890 49420 48900
rect 50000 48378 51688 49802
rect 51752 48378 51772 49802
rect 52190 48970 52250 50600
rect 52170 48960 52250 48970
rect 52170 48900 52180 48960
rect 52240 48900 52250 48960
rect 52170 48890 52250 48900
rect 50000 48350 51772 48378
rect 50000 48092 51772 48120
rect 49220 47250 49300 47260
rect 49220 47190 49230 47250
rect 49290 47190 49300 47250
rect 49220 47180 49300 47190
rect 50000 46668 51688 48092
rect 51752 46668 51772 48092
rect 52310 47260 52370 59150
rect 52290 47250 52370 47260
rect 52290 47190 52300 47250
rect 52360 47190 52370 47250
rect 52290 47180 52370 47190
rect 50000 46640 51772 46668
rect 50000 46382 51772 46410
rect 49100 45540 49180 45550
rect 49100 45480 49110 45540
rect 49170 45480 49180 45540
rect 49100 45470 49180 45480
rect 49100 43840 49160 45470
rect 50000 44958 51688 46382
rect 51752 44958 51772 46382
rect 52430 45550 52490 60850
rect 52410 45540 52490 45550
rect 52410 45480 52420 45540
rect 52480 45480 52490 45540
rect 52410 45470 52490 45480
rect 50000 44930 51772 44958
rect 50000 44672 51772 44700
rect 49100 43830 49180 43840
rect 49100 43770 49110 43830
rect 49170 43770 49180 43830
rect 49100 43760 49180 43770
rect 50000 43248 51688 44672
rect 51752 43248 51772 44672
rect 52430 43840 52490 45470
rect 52410 43830 52490 43840
rect 52410 43770 52420 43830
rect 52480 43770 52490 43830
rect 52410 43760 52490 43770
rect 50000 43220 51772 43248
rect 50000 42962 51772 42990
rect 48980 42120 49060 42130
rect 47540 42060 47550 42120
rect 47610 42060 47620 42120
rect 47540 42050 47620 42060
rect 45010 41510 46782 41538
rect 45010 41252 46782 41280
rect 43990 40420 44070 40430
rect 42550 40350 42630 40360
rect 43990 40360 44000 40420
rect 44060 40360 44070 40420
rect 43990 40350 44070 40360
rect 43990 40220 44050 40350
rect 43990 40210 44070 40220
rect 43990 40150 44000 40210
rect 44060 40150 44070 40210
rect 43990 40140 44070 40150
rect 40020 39800 41792 39828
rect 45010 39828 46698 41252
rect 46762 39828 46782 41252
rect 47560 40420 47620 42050
rect 48980 42060 48990 42120
rect 49050 42060 49060 42120
rect 48980 42050 49060 42060
rect 47540 40410 47620 40420
rect 48150 40630 48290 40660
rect 48150 40560 48180 40630
rect 48260 40560 48290 40630
rect 48150 40520 48290 40560
rect 48150 40450 48180 40520
rect 48260 40450 48290 40520
rect 48150 40410 48290 40450
rect 48980 40420 49040 42050
rect 50000 41538 51688 42962
rect 51752 41538 51772 42962
rect 52550 42130 52610 64280
rect 53970 64290 53980 64350
rect 54040 64290 54050 64350
rect 53970 64280 54050 64290
rect 53140 62860 53280 62890
rect 53140 62790 53170 62860
rect 53250 62790 53280 62860
rect 53140 62750 53280 62790
rect 53140 62680 53170 62750
rect 53250 62680 53280 62750
rect 53140 62640 53280 62680
rect 53140 61150 53280 61180
rect 53140 61080 53170 61150
rect 53250 61080 53280 61150
rect 53140 61040 53280 61080
rect 53140 60970 53170 61040
rect 53250 60970 53280 61040
rect 53140 60930 53280 60970
rect 53140 59440 53280 59470
rect 53140 59370 53170 59440
rect 53250 59370 53280 59440
rect 53140 59330 53280 59370
rect 53140 59260 53170 59330
rect 53250 59260 53280 59330
rect 53140 59220 53280 59260
rect 53140 57730 53280 57760
rect 53140 57660 53170 57730
rect 53250 57660 53280 57730
rect 53140 57620 53280 57660
rect 53140 57550 53170 57620
rect 53250 57550 53280 57620
rect 53140 57510 53280 57550
rect 53140 56020 53280 56050
rect 53140 55950 53170 56020
rect 53250 55950 53280 56020
rect 53140 55910 53280 55950
rect 53140 55840 53170 55910
rect 53250 55840 53280 55910
rect 53140 55800 53280 55840
rect 53140 54310 53280 54340
rect 53140 54240 53170 54310
rect 53250 54240 53280 54310
rect 53140 54200 53280 54240
rect 53140 54130 53170 54200
rect 53250 54130 53280 54200
rect 53140 54090 53280 54130
rect 53140 52600 53280 52630
rect 53140 52530 53170 52600
rect 53250 52530 53280 52600
rect 53140 52490 53280 52530
rect 53140 52420 53170 52490
rect 53250 52420 53280 52490
rect 53140 52380 53280 52420
rect 53140 50890 53280 50920
rect 53140 50820 53170 50890
rect 53250 50820 53280 50890
rect 53140 50780 53280 50820
rect 53140 50710 53170 50780
rect 53250 50710 53280 50780
rect 53140 50670 53280 50710
rect 53140 49180 53280 49210
rect 53140 49110 53170 49180
rect 53250 49110 53280 49180
rect 53140 49070 53280 49110
rect 53140 49000 53170 49070
rect 53250 49000 53280 49070
rect 53140 48960 53280 49000
rect 53140 47470 53280 47500
rect 53140 47400 53170 47470
rect 53250 47400 53280 47470
rect 53140 47360 53280 47400
rect 53140 47290 53170 47360
rect 53250 47290 53280 47360
rect 53140 47250 53280 47290
rect 53140 45760 53280 45790
rect 53140 45690 53170 45760
rect 53250 45690 53280 45760
rect 53140 45650 53280 45690
rect 53140 45580 53170 45650
rect 53250 45580 53280 45650
rect 53140 45540 53280 45580
rect 53140 44050 53280 44080
rect 53140 43980 53170 44050
rect 53250 43980 53280 44050
rect 53140 43940 53280 43980
rect 53140 43870 53170 43940
rect 53250 43870 53280 43940
rect 53140 43830 53280 43870
rect 52530 42120 52610 42130
rect 53140 42340 53280 42370
rect 53140 42270 53170 42340
rect 53250 42270 53280 42340
rect 53140 42230 53280 42270
rect 53140 42160 53170 42230
rect 53250 42160 53280 42230
rect 53140 42120 53280 42160
rect 53970 42130 54030 64280
rect 54990 63768 56678 65192
rect 56742 63768 56762 65192
rect 57540 64360 57600 65990
rect 58960 66000 58970 66060
rect 59030 66000 59040 66060
rect 58960 65990 59040 66000
rect 57520 64350 57600 64360
rect 58130 64570 58270 64600
rect 58130 64500 58160 64570
rect 58240 64500 58270 64570
rect 58130 64460 58270 64500
rect 58130 64390 58160 64460
rect 58240 64390 58270 64460
rect 58130 64350 58270 64390
rect 58960 64360 59020 65990
rect 59980 65478 61668 66902
rect 61732 65478 61752 66902
rect 64970 66902 66742 66930
rect 62510 66580 62590 66590
rect 62510 66520 62520 66580
rect 62580 66520 62590 66580
rect 62510 66510 62590 66520
rect 62530 66070 62590 66510
rect 63950 66580 64030 66590
rect 63950 66520 63960 66580
rect 64020 66520 64030 66580
rect 63950 66510 64030 66520
rect 62510 66060 62590 66070
rect 63120 66280 63260 66310
rect 63120 66210 63150 66280
rect 63230 66210 63260 66280
rect 63120 66170 63260 66210
rect 63120 66100 63150 66170
rect 63230 66100 63260 66170
rect 63120 66060 63260 66100
rect 63950 66070 64010 66510
rect 63950 66060 64030 66070
rect 62510 66000 62520 66060
rect 62580 66000 62590 66060
rect 62510 65990 62590 66000
rect 59980 65450 61752 65478
rect 59980 65192 61752 65220
rect 58960 64350 59040 64360
rect 57520 64290 57530 64350
rect 57590 64290 57600 64350
rect 57520 64280 57600 64290
rect 54990 63740 56762 63768
rect 54990 63482 56762 63510
rect 54090 63160 54170 63170
rect 54090 63100 54100 63160
rect 54160 63100 54170 63160
rect 54090 63090 54170 63100
rect 54090 62650 54150 63090
rect 54090 62640 54170 62650
rect 54090 62580 54100 62640
rect 54160 62580 54170 62640
rect 54090 62570 54170 62580
rect 54090 60930 54150 62570
rect 54990 62058 56678 63482
rect 56742 62058 56762 63482
rect 57400 63160 57480 63170
rect 57400 63100 57410 63160
rect 57470 63100 57480 63160
rect 57400 63090 57480 63100
rect 57420 62650 57480 63090
rect 57400 62640 57480 62650
rect 57400 62580 57410 62640
rect 57470 62580 57480 62640
rect 57400 62570 57480 62580
rect 54990 62030 56762 62058
rect 54990 61772 56762 61800
rect 54090 60920 54170 60930
rect 54090 60860 54100 60920
rect 54160 60860 54170 60920
rect 54090 60850 54170 60860
rect 54090 45550 54150 60850
rect 54990 60348 56678 61772
rect 56742 60348 56762 61772
rect 57420 60930 57480 62570
rect 57400 60920 57480 60930
rect 57400 60860 57410 60920
rect 57470 60860 57480 60920
rect 57400 60850 57480 60860
rect 54990 60320 56762 60348
rect 54990 60062 56762 60090
rect 54210 59740 54290 59750
rect 54210 59680 54220 59740
rect 54280 59680 54290 59740
rect 54210 59670 54290 59680
rect 54210 59230 54270 59670
rect 54210 59220 54290 59230
rect 54210 59160 54220 59220
rect 54280 59160 54290 59220
rect 54210 59150 54290 59160
rect 54210 47260 54270 59150
rect 54990 58638 56678 60062
rect 56742 58638 56762 60062
rect 57280 59740 57360 59750
rect 57280 59680 57290 59740
rect 57350 59680 57360 59740
rect 57280 59670 57360 59680
rect 57300 59230 57360 59670
rect 57280 59220 57360 59230
rect 57280 59160 57290 59220
rect 57350 59160 57360 59220
rect 57280 59150 57360 59160
rect 54990 58610 56762 58638
rect 54990 58352 56762 58380
rect 54330 58030 54410 58040
rect 54330 57970 54340 58030
rect 54400 57970 54410 58030
rect 54330 57960 54410 57970
rect 54330 57520 54390 57960
rect 54330 57510 54410 57520
rect 54330 57450 54340 57510
rect 54400 57450 54410 57510
rect 54330 57440 54410 57450
rect 54330 55810 54390 57440
rect 54990 56928 56678 58352
rect 56742 56928 56762 58352
rect 57160 58030 57240 58040
rect 57160 57970 57170 58030
rect 57230 57970 57240 58030
rect 57160 57960 57240 57970
rect 57180 57520 57240 57960
rect 57160 57510 57240 57520
rect 57160 57450 57170 57510
rect 57230 57450 57240 57510
rect 57160 57440 57240 57450
rect 54990 56900 56762 56928
rect 54990 56642 56762 56670
rect 54330 55800 54410 55810
rect 54330 55740 54340 55800
rect 54400 55740 54410 55800
rect 54330 55730 54410 55740
rect 54330 54100 54390 55730
rect 54990 55218 56678 56642
rect 56742 55218 56762 56642
rect 57180 55810 57240 57440
rect 57160 55800 57240 55810
rect 57160 55740 57170 55800
rect 57230 55740 57240 55800
rect 57160 55730 57240 55740
rect 54990 55190 56762 55218
rect 54990 54932 56762 54960
rect 54330 54090 54410 54100
rect 54330 54030 54340 54090
rect 54400 54030 54410 54090
rect 54330 54020 54410 54030
rect 54330 52390 54390 54020
rect 54990 53508 56678 54932
rect 56742 53508 56762 54932
rect 57180 54100 57240 55730
rect 57160 54090 57240 54100
rect 57160 54030 57170 54090
rect 57230 54030 57240 54090
rect 57160 54020 57240 54030
rect 54990 53480 56762 53508
rect 54990 53222 56762 53250
rect 54330 52380 54410 52390
rect 54330 52320 54340 52380
rect 54400 52320 54410 52380
rect 54330 52310 54410 52320
rect 54330 50680 54390 52310
rect 54990 51798 56678 53222
rect 56742 51798 56762 53222
rect 57180 52390 57240 54020
rect 57160 52380 57240 52390
rect 57160 52320 57170 52380
rect 57230 52320 57240 52380
rect 57160 52310 57240 52320
rect 54990 51770 56762 51798
rect 54990 51512 56762 51540
rect 54330 50670 54410 50680
rect 54330 50610 54340 50670
rect 54400 50610 54410 50670
rect 54330 50600 54410 50610
rect 54330 48970 54390 50600
rect 54990 50088 56678 51512
rect 56742 50088 56762 51512
rect 57180 50680 57240 52310
rect 57160 50670 57240 50680
rect 57160 50610 57170 50670
rect 57230 50610 57240 50670
rect 57160 50600 57240 50610
rect 54990 50060 56762 50088
rect 54990 49802 56762 49830
rect 54330 48960 54410 48970
rect 54330 48900 54340 48960
rect 54400 48900 54410 48960
rect 54330 48890 54410 48900
rect 54990 48378 56678 49802
rect 56742 48378 56762 49802
rect 57180 48970 57240 50600
rect 57160 48960 57240 48970
rect 57160 48900 57170 48960
rect 57230 48900 57240 48960
rect 57160 48890 57240 48900
rect 54990 48350 56762 48378
rect 54990 48092 56762 48120
rect 54210 47250 54290 47260
rect 54210 47190 54220 47250
rect 54280 47190 54290 47250
rect 54210 47180 54290 47190
rect 54990 46668 56678 48092
rect 56742 46668 56762 48092
rect 57300 47260 57360 59150
rect 57280 47250 57360 47260
rect 57280 47190 57290 47250
rect 57350 47190 57360 47250
rect 57280 47180 57360 47190
rect 54990 46640 56762 46668
rect 54990 46382 56762 46410
rect 54090 45540 54170 45550
rect 54090 45480 54100 45540
rect 54160 45480 54170 45540
rect 54090 45470 54170 45480
rect 54090 43840 54150 45470
rect 54990 44958 56678 46382
rect 56742 44958 56762 46382
rect 57420 45550 57480 60850
rect 57400 45540 57480 45550
rect 57400 45480 57410 45540
rect 57470 45480 57480 45540
rect 57400 45470 57480 45480
rect 54990 44930 56762 44958
rect 54990 44672 56762 44700
rect 54090 43830 54170 43840
rect 54090 43770 54100 43830
rect 54160 43770 54170 43830
rect 54090 43760 54170 43770
rect 54990 43248 56678 44672
rect 56742 43248 56762 44672
rect 57420 43840 57480 45470
rect 57400 43830 57480 43840
rect 57400 43770 57410 43830
rect 57470 43770 57480 43830
rect 57400 43760 57480 43770
rect 54990 43220 56762 43248
rect 54990 42962 56762 42990
rect 53970 42120 54050 42130
rect 52530 42060 52540 42120
rect 52600 42060 52610 42120
rect 52530 42050 52610 42060
rect 50000 41510 51772 41538
rect 50000 41252 51772 41280
rect 48980 40410 49060 40420
rect 47540 40350 47550 40410
rect 47610 40350 47620 40410
rect 47540 40340 47620 40350
rect 48980 40350 48990 40410
rect 49050 40350 49060 40410
rect 48980 40340 49060 40350
rect 45010 39800 46782 39828
rect 50000 39828 51688 41252
rect 51752 39828 51772 41252
rect 52550 40420 52610 42050
rect 53970 42060 53980 42120
rect 54040 42060 54050 42120
rect 53970 42050 54050 42060
rect 52530 40410 52610 40420
rect 53140 40630 53280 40660
rect 53140 40560 53170 40630
rect 53250 40560 53280 40630
rect 53140 40520 53280 40560
rect 53140 40450 53170 40520
rect 53250 40450 53280 40520
rect 53140 40410 53280 40450
rect 53970 40420 54030 42050
rect 54990 41538 56678 42962
rect 56742 41538 56762 42962
rect 57540 42130 57600 64280
rect 58960 64290 58970 64350
rect 59030 64290 59040 64350
rect 58960 64280 59040 64290
rect 58130 62860 58270 62890
rect 58130 62790 58160 62860
rect 58240 62790 58270 62860
rect 58130 62750 58270 62790
rect 58130 62680 58160 62750
rect 58240 62680 58270 62750
rect 58130 62640 58270 62680
rect 58130 61150 58270 61180
rect 58130 61080 58160 61150
rect 58240 61080 58270 61150
rect 58130 61040 58270 61080
rect 58130 60970 58160 61040
rect 58240 60970 58270 61040
rect 58130 60930 58270 60970
rect 58130 59440 58270 59470
rect 58130 59370 58160 59440
rect 58240 59370 58270 59440
rect 58130 59330 58270 59370
rect 58130 59260 58160 59330
rect 58240 59260 58270 59330
rect 58130 59220 58270 59260
rect 58130 57730 58270 57760
rect 58130 57660 58160 57730
rect 58240 57660 58270 57730
rect 58130 57620 58270 57660
rect 58130 57550 58160 57620
rect 58240 57550 58270 57620
rect 58130 57510 58270 57550
rect 58130 56020 58270 56050
rect 58130 55950 58160 56020
rect 58240 55950 58270 56020
rect 58130 55910 58270 55950
rect 58130 55840 58160 55910
rect 58240 55840 58270 55910
rect 58130 55800 58270 55840
rect 58130 54310 58270 54340
rect 58130 54240 58160 54310
rect 58240 54240 58270 54310
rect 58130 54200 58270 54240
rect 58130 54130 58160 54200
rect 58240 54130 58270 54200
rect 58130 54090 58270 54130
rect 58130 52600 58270 52630
rect 58130 52530 58160 52600
rect 58240 52530 58270 52600
rect 58130 52490 58270 52530
rect 58130 52420 58160 52490
rect 58240 52420 58270 52490
rect 58130 52380 58270 52420
rect 58130 50890 58270 50920
rect 58130 50820 58160 50890
rect 58240 50820 58270 50890
rect 58130 50780 58270 50820
rect 58130 50710 58160 50780
rect 58240 50710 58270 50780
rect 58130 50670 58270 50710
rect 58130 49180 58270 49210
rect 58130 49110 58160 49180
rect 58240 49110 58270 49180
rect 58130 49070 58270 49110
rect 58130 49000 58160 49070
rect 58240 49000 58270 49070
rect 58130 48960 58270 49000
rect 58130 47470 58270 47500
rect 58130 47400 58160 47470
rect 58240 47400 58270 47470
rect 58130 47360 58270 47400
rect 58130 47290 58160 47360
rect 58240 47290 58270 47360
rect 58130 47250 58270 47290
rect 58130 45760 58270 45790
rect 58130 45690 58160 45760
rect 58240 45690 58270 45760
rect 58130 45650 58270 45690
rect 58130 45580 58160 45650
rect 58240 45580 58270 45650
rect 58130 45540 58270 45580
rect 58130 44050 58270 44080
rect 58130 43980 58160 44050
rect 58240 43980 58270 44050
rect 58130 43940 58270 43980
rect 58130 43870 58160 43940
rect 58240 43870 58270 43940
rect 58130 43830 58270 43870
rect 57520 42120 57600 42130
rect 58130 42340 58270 42370
rect 58130 42270 58160 42340
rect 58240 42270 58270 42340
rect 58130 42230 58270 42270
rect 58130 42160 58160 42230
rect 58240 42160 58270 42230
rect 58130 42120 58270 42160
rect 58960 42130 59020 64280
rect 59980 63768 61668 65192
rect 61732 63768 61752 65192
rect 62530 64360 62590 65990
rect 63950 66000 63960 66060
rect 64020 66000 64030 66060
rect 63950 65990 64030 66000
rect 62510 64350 62590 64360
rect 63120 64570 63260 64600
rect 63120 64500 63150 64570
rect 63230 64500 63260 64570
rect 63120 64460 63260 64500
rect 63120 64390 63150 64460
rect 63230 64390 63260 64460
rect 63120 64350 63260 64390
rect 63950 64360 64010 65990
rect 64970 65478 66658 66902
rect 66722 65478 66742 66902
rect 69960 66902 71732 66930
rect 67500 66580 67580 66590
rect 67500 66520 67510 66580
rect 67570 66520 67580 66580
rect 67500 66510 67580 66520
rect 67520 66070 67580 66510
rect 68940 66580 69020 66590
rect 68940 66520 68950 66580
rect 69010 66520 69020 66580
rect 68940 66510 69020 66520
rect 67500 66060 67580 66070
rect 68110 66280 68250 66310
rect 68110 66210 68140 66280
rect 68220 66210 68250 66280
rect 68110 66170 68250 66210
rect 68110 66100 68140 66170
rect 68220 66100 68250 66170
rect 68110 66060 68250 66100
rect 68940 66070 69000 66510
rect 68940 66060 69020 66070
rect 67500 66000 67510 66060
rect 67570 66000 67580 66060
rect 67500 65990 67580 66000
rect 64970 65450 66742 65478
rect 64970 65192 66742 65220
rect 63950 64350 64030 64360
rect 62510 64290 62520 64350
rect 62580 64290 62590 64350
rect 62510 64280 62590 64290
rect 59980 63740 61752 63768
rect 59980 63482 61752 63510
rect 59080 63160 59160 63170
rect 59080 63100 59090 63160
rect 59150 63100 59160 63160
rect 59080 63090 59160 63100
rect 59080 62650 59140 63090
rect 59080 62640 59160 62650
rect 59080 62580 59090 62640
rect 59150 62580 59160 62640
rect 59080 62570 59160 62580
rect 59080 60930 59140 62570
rect 59980 62058 61668 63482
rect 61732 62058 61752 63482
rect 62530 62650 62590 64280
rect 63950 64290 63960 64350
rect 64020 64290 64030 64350
rect 63950 64280 64030 64290
rect 62510 62640 62590 62650
rect 63120 62860 63260 62890
rect 63120 62790 63150 62860
rect 63230 62790 63260 62860
rect 63120 62750 63260 62790
rect 63120 62680 63150 62750
rect 63230 62680 63260 62750
rect 63120 62640 63260 62680
rect 63950 62650 64010 64280
rect 64970 63768 66658 65192
rect 66722 63768 66742 65192
rect 67520 64360 67580 65990
rect 68940 66000 68950 66060
rect 69010 66000 69020 66060
rect 68940 65990 69020 66000
rect 67500 64350 67580 64360
rect 68110 64570 68250 64600
rect 68110 64500 68140 64570
rect 68220 64500 68250 64570
rect 68110 64460 68250 64500
rect 68110 64390 68140 64460
rect 68220 64390 68250 64460
rect 68110 64350 68250 64390
rect 68940 64360 69000 65990
rect 69960 65478 71648 66902
rect 71712 65478 71732 66902
rect 74950 66902 76722 66930
rect 72490 66580 72570 66590
rect 72490 66520 72500 66580
rect 72560 66520 72570 66580
rect 72490 66510 72570 66520
rect 72510 66070 72570 66510
rect 73930 66580 74010 66590
rect 73930 66520 73940 66580
rect 74000 66520 74010 66580
rect 73930 66510 74010 66520
rect 72490 66060 72570 66070
rect 73100 66280 73240 66310
rect 73100 66210 73130 66280
rect 73210 66210 73240 66280
rect 73100 66170 73240 66210
rect 73100 66100 73130 66170
rect 73210 66100 73240 66170
rect 73100 66060 73240 66100
rect 73930 66070 73990 66510
rect 73930 66060 74010 66070
rect 72490 66000 72500 66060
rect 72560 66000 72570 66060
rect 72490 65990 72570 66000
rect 69960 65450 71732 65478
rect 69960 65192 71732 65220
rect 68940 64350 69020 64360
rect 67500 64290 67510 64350
rect 67570 64290 67580 64350
rect 67500 64280 67580 64290
rect 64970 63740 66742 63768
rect 64970 63482 66742 63510
rect 63950 62640 64030 62650
rect 62510 62580 62520 62640
rect 62580 62580 62590 62640
rect 62510 62570 62590 62580
rect 59980 62030 61752 62058
rect 59980 61772 61752 61800
rect 59080 60920 59160 60930
rect 59080 60860 59090 60920
rect 59150 60860 59160 60920
rect 59080 60850 59160 60860
rect 59080 45550 59140 60850
rect 59980 60348 61668 61772
rect 61732 60348 61752 61772
rect 62530 60940 62590 62570
rect 63950 62580 63960 62640
rect 64020 62580 64030 62640
rect 63950 62570 64030 62580
rect 62510 60930 62590 60940
rect 63120 61150 63260 61180
rect 63120 61080 63150 61150
rect 63230 61080 63260 61150
rect 63120 61040 63260 61080
rect 63120 60970 63150 61040
rect 63230 60970 63260 61040
rect 63120 60930 63260 60970
rect 63950 60940 64010 62570
rect 64970 62058 66658 63482
rect 66722 62058 66742 63482
rect 67520 62650 67580 64280
rect 68940 64290 68950 64350
rect 69010 64290 69020 64350
rect 68940 64280 69020 64290
rect 67500 62640 67580 62650
rect 68110 62860 68250 62890
rect 68110 62790 68140 62860
rect 68220 62790 68250 62860
rect 68110 62750 68250 62790
rect 68110 62680 68140 62750
rect 68220 62680 68250 62750
rect 68110 62640 68250 62680
rect 68940 62650 69000 64280
rect 69960 63768 71648 65192
rect 71712 63768 71732 65192
rect 72510 64360 72570 65990
rect 73930 66000 73940 66060
rect 74000 66000 74010 66060
rect 73930 65990 74010 66000
rect 72490 64350 72570 64360
rect 73100 64570 73240 64600
rect 73100 64500 73130 64570
rect 73210 64500 73240 64570
rect 73100 64460 73240 64500
rect 73100 64390 73130 64460
rect 73210 64390 73240 64460
rect 73100 64350 73240 64390
rect 73930 64360 73990 65990
rect 74950 65478 76638 66902
rect 76702 65478 76722 66902
rect 77480 66580 77560 66590
rect 77480 66520 77490 66580
rect 77550 66520 77560 66580
rect 77480 66510 77560 66520
rect 77500 66070 77560 66510
rect 78920 66580 79000 66590
rect 78920 66520 78930 66580
rect 78990 66520 79000 66580
rect 78920 66510 79000 66520
rect 77480 66060 77560 66070
rect 78090 66280 78230 66310
rect 78090 66210 78120 66280
rect 78200 66210 78230 66280
rect 78090 66170 78230 66210
rect 78090 66100 78120 66170
rect 78200 66100 78230 66170
rect 78090 66060 78230 66100
rect 78920 66070 78980 66510
rect 78920 66060 79000 66070
rect 77480 66000 77490 66060
rect 77550 66000 77560 66060
rect 77480 65990 77560 66000
rect 74950 65450 76722 65478
rect 74950 65192 76722 65220
rect 73930 64350 74010 64360
rect 72490 64290 72500 64350
rect 72560 64290 72570 64350
rect 72490 64280 72570 64290
rect 69960 63740 71732 63768
rect 69960 63482 71732 63510
rect 68940 62640 69020 62650
rect 67500 62580 67510 62640
rect 67570 62580 67580 62640
rect 67500 62570 67580 62580
rect 64970 62030 66742 62058
rect 64970 61772 66742 61800
rect 63950 60930 64030 60940
rect 62510 60870 62520 60930
rect 62580 60870 62590 60930
rect 62510 60860 62590 60870
rect 59980 60320 61752 60348
rect 59980 60062 61752 60090
rect 59200 59740 59280 59750
rect 59200 59680 59210 59740
rect 59270 59680 59280 59740
rect 59200 59670 59280 59680
rect 59200 59230 59260 59670
rect 59200 59220 59280 59230
rect 59200 59160 59210 59220
rect 59270 59160 59280 59220
rect 59200 59150 59280 59160
rect 59200 47260 59260 59150
rect 59980 58638 61668 60062
rect 61732 58638 61752 60062
rect 62390 59740 62470 59750
rect 62390 59680 62400 59740
rect 62460 59680 62470 59740
rect 62390 59670 62470 59680
rect 62410 59230 62470 59670
rect 62390 59220 62470 59230
rect 62390 59160 62400 59220
rect 62460 59160 62470 59220
rect 62390 59150 62470 59160
rect 59980 58610 61752 58638
rect 59980 58352 61752 58380
rect 59320 58030 59400 58040
rect 59320 57970 59330 58030
rect 59390 57970 59400 58030
rect 59320 57960 59400 57970
rect 59320 57520 59380 57960
rect 59320 57510 59400 57520
rect 59320 57450 59330 57510
rect 59390 57450 59400 57510
rect 59320 57440 59400 57450
rect 59320 55810 59380 57440
rect 59980 56928 61668 58352
rect 61732 56928 61752 58352
rect 62410 57520 62470 59150
rect 62390 57510 62470 57520
rect 62390 57450 62400 57510
rect 62460 57450 62470 57510
rect 62390 57440 62470 57450
rect 59980 56900 61752 56928
rect 59980 56642 61752 56670
rect 59320 55800 59400 55810
rect 59320 55740 59330 55800
rect 59390 55740 59400 55800
rect 59320 55730 59400 55740
rect 59320 54100 59380 55730
rect 59980 55218 61668 56642
rect 61732 55218 61752 56642
rect 62410 55810 62470 57440
rect 62390 55800 62470 55810
rect 62390 55740 62400 55800
rect 62460 55740 62470 55800
rect 62390 55730 62470 55740
rect 59980 55190 61752 55218
rect 59980 54932 61752 54960
rect 59320 54090 59400 54100
rect 59320 54030 59330 54090
rect 59390 54030 59400 54090
rect 59320 54020 59400 54030
rect 59320 52390 59380 54020
rect 59980 53508 61668 54932
rect 61732 53508 61752 54932
rect 62410 54100 62470 55730
rect 62390 54090 62470 54100
rect 62390 54030 62400 54090
rect 62460 54030 62470 54090
rect 62390 54020 62470 54030
rect 59980 53480 61752 53508
rect 59980 53222 61752 53250
rect 59320 52380 59400 52390
rect 59320 52320 59330 52380
rect 59390 52320 59400 52380
rect 59320 52310 59400 52320
rect 59320 50680 59380 52310
rect 59980 51798 61668 53222
rect 61732 51798 61752 53222
rect 62410 52390 62470 54020
rect 62390 52380 62470 52390
rect 62390 52320 62400 52380
rect 62460 52320 62470 52380
rect 62390 52310 62470 52320
rect 59980 51770 61752 51798
rect 59980 51512 61752 51540
rect 59320 50670 59400 50680
rect 59320 50610 59330 50670
rect 59390 50610 59400 50670
rect 59320 50600 59400 50610
rect 59320 48970 59380 50600
rect 59980 50088 61668 51512
rect 61732 50088 61752 51512
rect 62410 50680 62470 52310
rect 62390 50670 62470 50680
rect 62390 50610 62400 50670
rect 62460 50610 62470 50670
rect 62390 50600 62470 50610
rect 59980 50060 61752 50088
rect 59980 49802 61752 49830
rect 59320 48960 59400 48970
rect 59320 48900 59330 48960
rect 59390 48900 59400 48960
rect 59320 48890 59400 48900
rect 59980 48378 61668 49802
rect 61732 48378 61752 49802
rect 62410 48970 62470 50600
rect 62390 48960 62470 48970
rect 62390 48900 62400 48960
rect 62460 48900 62470 48960
rect 62390 48890 62470 48900
rect 59980 48350 61752 48378
rect 59980 48092 61752 48120
rect 59200 47250 59280 47260
rect 59200 47190 59210 47250
rect 59270 47190 59280 47250
rect 59200 47180 59280 47190
rect 59980 46668 61668 48092
rect 61732 46668 61752 48092
rect 62410 47260 62470 48890
rect 62390 47250 62470 47260
rect 62390 47190 62400 47250
rect 62460 47190 62470 47250
rect 62390 47180 62470 47190
rect 59980 46640 61752 46668
rect 59980 46382 61752 46410
rect 59080 45540 59160 45550
rect 59080 45480 59090 45540
rect 59150 45480 59160 45540
rect 59080 45470 59160 45480
rect 59080 43840 59140 45470
rect 59980 44958 61668 46382
rect 61732 44958 61752 46382
rect 62530 45550 62590 60860
rect 63950 60870 63960 60930
rect 64020 60870 64030 60930
rect 63950 60860 64030 60870
rect 63120 59440 63260 59470
rect 63120 59370 63150 59440
rect 63230 59370 63260 59440
rect 63120 59330 63260 59370
rect 63120 59260 63150 59330
rect 63230 59260 63260 59330
rect 63120 59220 63260 59260
rect 63120 57730 63260 57760
rect 63120 57660 63150 57730
rect 63230 57660 63260 57730
rect 63120 57620 63260 57660
rect 63120 57550 63150 57620
rect 63230 57550 63260 57620
rect 63120 57510 63260 57550
rect 63120 56020 63260 56050
rect 63120 55950 63150 56020
rect 63230 55950 63260 56020
rect 63120 55910 63260 55950
rect 63120 55840 63150 55910
rect 63230 55840 63260 55910
rect 63120 55800 63260 55840
rect 63120 54310 63260 54340
rect 63120 54240 63150 54310
rect 63230 54240 63260 54310
rect 63120 54200 63260 54240
rect 63120 54130 63150 54200
rect 63230 54130 63260 54200
rect 63120 54090 63260 54130
rect 63120 52600 63260 52630
rect 63120 52530 63150 52600
rect 63230 52530 63260 52600
rect 63120 52490 63260 52530
rect 63120 52420 63150 52490
rect 63230 52420 63260 52490
rect 63120 52380 63260 52420
rect 63120 50890 63260 50920
rect 63120 50820 63150 50890
rect 63230 50820 63260 50890
rect 63120 50780 63260 50820
rect 63120 50710 63150 50780
rect 63230 50710 63260 50780
rect 63120 50670 63260 50710
rect 63120 49180 63260 49210
rect 63120 49110 63150 49180
rect 63230 49110 63260 49180
rect 63120 49070 63260 49110
rect 63120 49000 63150 49070
rect 63230 49000 63260 49070
rect 63120 48960 63260 49000
rect 63120 47470 63260 47500
rect 63120 47400 63150 47470
rect 63230 47400 63260 47470
rect 63120 47360 63260 47400
rect 63120 47290 63150 47360
rect 63230 47290 63260 47360
rect 63120 47250 63260 47290
rect 62510 45540 62590 45550
rect 63120 45760 63260 45790
rect 63120 45690 63150 45760
rect 63230 45690 63260 45760
rect 63120 45650 63260 45690
rect 63120 45580 63150 45650
rect 63230 45580 63260 45650
rect 63120 45540 63260 45580
rect 63950 45550 64010 60860
rect 64970 60348 66658 61772
rect 66722 60348 66742 61772
rect 67520 60940 67580 62570
rect 68940 62580 68950 62640
rect 69010 62580 69020 62640
rect 68940 62570 69020 62580
rect 67500 60930 67580 60940
rect 68110 61150 68250 61180
rect 68110 61080 68140 61150
rect 68220 61080 68250 61150
rect 68110 61040 68250 61080
rect 68110 60970 68140 61040
rect 68220 60970 68250 61040
rect 68110 60930 68250 60970
rect 68940 60940 69000 62570
rect 69960 62058 71648 63482
rect 71712 62058 71732 63482
rect 72510 62650 72570 64280
rect 73930 64290 73940 64350
rect 74000 64290 74010 64350
rect 73930 64280 74010 64290
rect 72490 62640 72570 62650
rect 73100 62860 73240 62890
rect 73100 62790 73130 62860
rect 73210 62790 73240 62860
rect 73100 62750 73240 62790
rect 73100 62680 73130 62750
rect 73210 62680 73240 62750
rect 73100 62640 73240 62680
rect 73930 62650 73990 64280
rect 74950 63768 76638 65192
rect 76702 63768 76722 65192
rect 77500 64360 77560 65990
rect 78920 66000 78930 66060
rect 78990 66000 79000 66060
rect 78920 65990 79000 66000
rect 77480 64350 77560 64360
rect 78090 64570 78230 64600
rect 78090 64500 78120 64570
rect 78200 64500 78230 64570
rect 78090 64460 78230 64500
rect 78090 64390 78120 64460
rect 78200 64390 78230 64460
rect 78090 64350 78230 64390
rect 78920 64360 78980 65990
rect 78920 64350 79000 64360
rect 77480 64290 77490 64350
rect 77550 64290 77560 64350
rect 77480 64280 77560 64290
rect 74950 63740 76722 63768
rect 74950 63482 76722 63510
rect 73930 62640 74010 62650
rect 72490 62580 72500 62640
rect 72560 62580 72570 62640
rect 72490 62570 72570 62580
rect 69960 62030 71732 62058
rect 69960 61772 71732 61800
rect 68940 60930 69020 60940
rect 67500 60870 67510 60930
rect 67570 60870 67580 60930
rect 67500 60860 67580 60870
rect 64970 60320 66742 60348
rect 64970 60062 66742 60090
rect 64070 59740 64150 59750
rect 64070 59680 64080 59740
rect 64140 59680 64150 59740
rect 64070 59670 64150 59680
rect 64070 59230 64130 59670
rect 64070 59220 64150 59230
rect 64070 59160 64080 59220
rect 64140 59160 64150 59220
rect 64070 59150 64150 59160
rect 64070 57520 64130 59150
rect 64970 58638 66658 60062
rect 66722 58638 66742 60062
rect 67380 59740 67460 59750
rect 67380 59680 67390 59740
rect 67450 59680 67460 59740
rect 67380 59670 67460 59680
rect 67400 59230 67460 59670
rect 67380 59220 67460 59230
rect 67380 59160 67390 59220
rect 67450 59160 67460 59220
rect 67380 59150 67460 59160
rect 64970 58610 66742 58638
rect 64970 58352 66742 58380
rect 64070 57510 64150 57520
rect 64070 57450 64080 57510
rect 64140 57450 64150 57510
rect 64070 57440 64150 57450
rect 64070 55810 64130 57440
rect 64970 56928 66658 58352
rect 66722 56928 66742 58352
rect 67400 57520 67460 59150
rect 67380 57510 67460 57520
rect 67380 57450 67390 57510
rect 67450 57450 67460 57510
rect 67380 57440 67460 57450
rect 64970 56900 66742 56928
rect 64970 56642 66742 56670
rect 64070 55800 64150 55810
rect 64070 55740 64080 55800
rect 64140 55740 64150 55800
rect 64070 55730 64150 55740
rect 64070 54100 64130 55730
rect 64970 55218 66658 56642
rect 66722 55218 66742 56642
rect 67400 55810 67460 57440
rect 67380 55800 67460 55810
rect 67380 55740 67390 55800
rect 67450 55740 67460 55800
rect 67380 55730 67460 55740
rect 64970 55190 66742 55218
rect 64970 54932 66742 54960
rect 64070 54090 64150 54100
rect 64070 54030 64080 54090
rect 64140 54030 64150 54090
rect 64070 54020 64150 54030
rect 64070 52390 64130 54020
rect 64970 53508 66658 54932
rect 66722 53508 66742 54932
rect 67400 54100 67460 55730
rect 67380 54090 67460 54100
rect 67380 54030 67390 54090
rect 67450 54030 67460 54090
rect 67380 54020 67460 54030
rect 64970 53480 66742 53508
rect 64970 53222 66742 53250
rect 64070 52380 64150 52390
rect 64070 52320 64080 52380
rect 64140 52320 64150 52380
rect 64070 52310 64150 52320
rect 64070 50680 64130 52310
rect 64970 51798 66658 53222
rect 66722 51798 66742 53222
rect 67400 52390 67460 54020
rect 67380 52380 67460 52390
rect 67380 52320 67390 52380
rect 67450 52320 67460 52380
rect 67380 52310 67460 52320
rect 64970 51770 66742 51798
rect 64970 51512 66742 51540
rect 64070 50670 64150 50680
rect 64070 50610 64080 50670
rect 64140 50610 64150 50670
rect 64070 50600 64150 50610
rect 64070 48970 64130 50600
rect 64970 50088 66658 51512
rect 66722 50088 66742 51512
rect 67400 50680 67460 52310
rect 67380 50670 67460 50680
rect 67380 50610 67390 50670
rect 67450 50610 67460 50670
rect 67380 50600 67460 50610
rect 64970 50060 66742 50088
rect 64970 49802 66742 49830
rect 64070 48960 64150 48970
rect 64070 48900 64080 48960
rect 64140 48900 64150 48960
rect 64070 48890 64150 48900
rect 64070 47260 64130 48890
rect 64970 48378 66658 49802
rect 66722 48378 66742 49802
rect 67400 48970 67460 50600
rect 67380 48960 67460 48970
rect 67380 48900 67390 48960
rect 67450 48900 67460 48960
rect 67380 48890 67460 48900
rect 64970 48350 66742 48378
rect 64970 48092 66742 48120
rect 64070 47250 64150 47260
rect 64070 47190 64080 47250
rect 64140 47190 64150 47250
rect 64070 47180 64150 47190
rect 64970 46668 66658 48092
rect 66722 46668 66742 48092
rect 67400 47260 67460 48890
rect 67380 47250 67460 47260
rect 67380 47190 67390 47250
rect 67450 47190 67460 47250
rect 67380 47180 67460 47190
rect 64970 46640 66742 46668
rect 64970 46382 66742 46410
rect 63950 45540 64030 45550
rect 62510 45480 62520 45540
rect 62580 45480 62590 45540
rect 62510 45470 62590 45480
rect 59980 44930 61752 44958
rect 59980 44672 61752 44700
rect 59080 43830 59160 43840
rect 59080 43770 59090 43830
rect 59150 43770 59160 43830
rect 59080 43760 59160 43770
rect 59980 43248 61668 44672
rect 61732 43248 61752 44672
rect 62530 43840 62590 45470
rect 63950 45480 63960 45540
rect 64020 45480 64030 45540
rect 63950 45470 64030 45480
rect 62510 43830 62590 43840
rect 63120 44050 63260 44080
rect 63120 43980 63150 44050
rect 63230 43980 63260 44050
rect 63120 43940 63260 43980
rect 63120 43870 63150 43940
rect 63230 43870 63260 43940
rect 63120 43830 63260 43870
rect 63950 43840 64010 45470
rect 64970 44958 66658 46382
rect 66722 44958 66742 46382
rect 67520 45550 67580 60860
rect 68940 60870 68950 60930
rect 69010 60870 69020 60930
rect 68940 60860 69020 60870
rect 68110 59440 68250 59470
rect 68110 59370 68140 59440
rect 68220 59370 68250 59440
rect 68110 59330 68250 59370
rect 68110 59260 68140 59330
rect 68220 59260 68250 59330
rect 68110 59220 68250 59260
rect 68110 57730 68250 57760
rect 68110 57660 68140 57730
rect 68220 57660 68250 57730
rect 68110 57620 68250 57660
rect 68110 57550 68140 57620
rect 68220 57550 68250 57620
rect 68110 57510 68250 57550
rect 68110 56020 68250 56050
rect 68110 55950 68140 56020
rect 68220 55950 68250 56020
rect 68110 55910 68250 55950
rect 68110 55840 68140 55910
rect 68220 55840 68250 55910
rect 68110 55800 68250 55840
rect 68110 54310 68250 54340
rect 68110 54240 68140 54310
rect 68220 54240 68250 54310
rect 68110 54200 68250 54240
rect 68110 54130 68140 54200
rect 68220 54130 68250 54200
rect 68110 54090 68250 54130
rect 68110 52600 68250 52630
rect 68110 52530 68140 52600
rect 68220 52530 68250 52600
rect 68110 52490 68250 52530
rect 68110 52420 68140 52490
rect 68220 52420 68250 52490
rect 68110 52380 68250 52420
rect 68110 50890 68250 50920
rect 68110 50820 68140 50890
rect 68220 50820 68250 50890
rect 68110 50780 68250 50820
rect 68110 50710 68140 50780
rect 68220 50710 68250 50780
rect 68110 50670 68250 50710
rect 68110 49180 68250 49210
rect 68110 49110 68140 49180
rect 68220 49110 68250 49180
rect 68110 49070 68250 49110
rect 68110 49000 68140 49070
rect 68220 49000 68250 49070
rect 68110 48960 68250 49000
rect 68110 47470 68250 47500
rect 68110 47400 68140 47470
rect 68220 47400 68250 47470
rect 68110 47360 68250 47400
rect 68110 47290 68140 47360
rect 68220 47290 68250 47360
rect 68110 47250 68250 47290
rect 67500 45540 67580 45550
rect 68110 45760 68250 45790
rect 68110 45690 68140 45760
rect 68220 45690 68250 45760
rect 68110 45650 68250 45690
rect 68110 45580 68140 45650
rect 68220 45580 68250 45650
rect 68110 45540 68250 45580
rect 68940 45550 69000 60860
rect 69960 60348 71648 61772
rect 71712 60348 71732 61772
rect 72510 60940 72570 62570
rect 73930 62580 73940 62640
rect 74000 62580 74010 62640
rect 73930 62570 74010 62580
rect 72490 60930 72570 60940
rect 73100 61150 73240 61180
rect 73100 61080 73130 61150
rect 73210 61080 73240 61150
rect 73100 61040 73240 61080
rect 73100 60970 73130 61040
rect 73210 60970 73240 61040
rect 73100 60930 73240 60970
rect 73930 60940 73990 62570
rect 74950 62058 76638 63482
rect 76702 62058 76722 63482
rect 77500 62650 77560 64280
rect 78920 64290 78930 64350
rect 78990 64290 79000 64350
rect 78920 64280 79000 64290
rect 77480 62640 77560 62650
rect 78090 62860 78230 62890
rect 78090 62790 78120 62860
rect 78200 62790 78230 62860
rect 78090 62750 78230 62790
rect 78090 62680 78120 62750
rect 78200 62680 78230 62750
rect 78090 62640 78230 62680
rect 78920 62650 78980 64280
rect 78920 62640 79000 62650
rect 77480 62580 77490 62640
rect 77550 62580 77560 62640
rect 77480 62570 77560 62580
rect 74950 62030 76722 62058
rect 74950 61772 76722 61800
rect 73930 60930 74010 60940
rect 72490 60870 72500 60930
rect 72560 60870 72570 60930
rect 72490 60860 72570 60870
rect 69960 60320 71732 60348
rect 69960 60062 71732 60090
rect 69060 59740 69140 59750
rect 69060 59680 69070 59740
rect 69130 59680 69140 59740
rect 69060 59670 69140 59680
rect 69060 59230 69120 59670
rect 69060 59220 69140 59230
rect 69060 59160 69070 59220
rect 69130 59160 69140 59220
rect 69060 59150 69140 59160
rect 69060 57520 69120 59150
rect 69960 58638 71648 60062
rect 71712 58638 71732 60062
rect 72510 59230 72570 60860
rect 73930 60870 73940 60930
rect 74000 60870 74010 60930
rect 73930 60860 74010 60870
rect 72490 59220 72570 59230
rect 73100 59440 73240 59470
rect 73100 59370 73130 59440
rect 73210 59370 73240 59440
rect 73100 59330 73240 59370
rect 73100 59260 73130 59330
rect 73210 59260 73240 59330
rect 73100 59220 73240 59260
rect 73930 59230 73990 60860
rect 74950 60348 76638 61772
rect 76702 60348 76722 61772
rect 77500 60940 77560 62570
rect 78920 62580 78930 62640
rect 78990 62580 79000 62640
rect 78920 62570 79000 62580
rect 77480 60930 77560 60940
rect 78090 61150 78230 61180
rect 78090 61080 78120 61150
rect 78200 61080 78230 61150
rect 78090 61040 78230 61080
rect 78090 60970 78120 61040
rect 78200 60970 78230 61040
rect 78090 60930 78230 60970
rect 78920 60940 78980 62570
rect 78920 60930 79000 60940
rect 77480 60870 77490 60930
rect 77550 60870 77560 60930
rect 77480 60860 77560 60870
rect 74950 60320 76722 60348
rect 74950 60062 76722 60090
rect 73930 59220 74010 59230
rect 72490 59160 72500 59220
rect 72560 59160 72570 59220
rect 72490 59150 72570 59160
rect 69960 58610 71732 58638
rect 69960 58352 71732 58380
rect 69060 57510 69140 57520
rect 69060 57450 69070 57510
rect 69130 57450 69140 57510
rect 69060 57440 69140 57450
rect 69060 55810 69120 57440
rect 69960 56928 71648 58352
rect 71712 56928 71732 58352
rect 72510 57520 72570 59150
rect 73930 59160 73940 59220
rect 74000 59160 74010 59220
rect 73930 59150 74010 59160
rect 72490 57510 72570 57520
rect 73100 57730 73240 57760
rect 73100 57660 73130 57730
rect 73210 57660 73240 57730
rect 73100 57620 73240 57660
rect 73100 57550 73130 57620
rect 73210 57550 73240 57620
rect 73100 57510 73240 57550
rect 73930 57520 73990 59150
rect 74950 58638 76638 60062
rect 76702 58638 76722 60062
rect 77500 59230 77560 60860
rect 78920 60870 78930 60930
rect 78990 60870 79000 60930
rect 78920 60860 79000 60870
rect 77480 59220 77560 59230
rect 78090 59440 78230 59470
rect 78090 59370 78120 59440
rect 78200 59370 78230 59440
rect 78090 59330 78230 59370
rect 78090 59260 78120 59330
rect 78200 59260 78230 59330
rect 78090 59220 78230 59260
rect 78920 59230 78980 60860
rect 78920 59220 79000 59230
rect 77480 59160 77490 59220
rect 77550 59160 77560 59220
rect 77480 59150 77560 59160
rect 74950 58610 76722 58638
rect 74950 58352 76722 58380
rect 73930 57510 74010 57520
rect 72490 57450 72500 57510
rect 72560 57450 72570 57510
rect 72490 57440 72570 57450
rect 69960 56900 71732 56928
rect 69960 56642 71732 56670
rect 69060 55800 69140 55810
rect 69060 55740 69070 55800
rect 69130 55740 69140 55800
rect 69060 55730 69140 55740
rect 69060 54100 69120 55730
rect 69960 55218 71648 56642
rect 71712 55218 71732 56642
rect 72510 55810 72570 57440
rect 73930 57450 73940 57510
rect 74000 57450 74010 57510
rect 73930 57440 74010 57450
rect 72490 55800 72570 55810
rect 73100 56020 73240 56050
rect 73100 55950 73130 56020
rect 73210 55950 73240 56020
rect 73100 55910 73240 55950
rect 73100 55840 73130 55910
rect 73210 55840 73240 55910
rect 73100 55800 73240 55840
rect 73930 55810 73990 57440
rect 74950 56928 76638 58352
rect 76702 56928 76722 58352
rect 77500 57520 77560 59150
rect 78920 59160 78930 59220
rect 78990 59160 79000 59220
rect 78920 59150 79000 59160
rect 77480 57510 77560 57520
rect 78090 57730 78230 57760
rect 78090 57660 78120 57730
rect 78200 57660 78230 57730
rect 78090 57620 78230 57660
rect 78090 57550 78120 57620
rect 78200 57550 78230 57620
rect 78090 57510 78230 57550
rect 78920 57520 78980 59150
rect 78920 57510 79000 57520
rect 77480 57450 77490 57510
rect 77550 57450 77560 57510
rect 77480 57440 77560 57450
rect 74950 56900 76722 56928
rect 74950 56642 76722 56670
rect 73930 55800 74010 55810
rect 72490 55740 72500 55800
rect 72560 55740 72570 55800
rect 72490 55730 72570 55740
rect 69960 55190 71732 55218
rect 69960 54932 71732 54960
rect 69060 54090 69140 54100
rect 69060 54030 69070 54090
rect 69130 54030 69140 54090
rect 69060 54020 69140 54030
rect 69060 52390 69120 54020
rect 69960 53508 71648 54932
rect 71712 53508 71732 54932
rect 72510 54100 72570 55730
rect 73930 55740 73940 55800
rect 74000 55740 74010 55800
rect 73930 55730 74010 55740
rect 72490 54090 72570 54100
rect 73100 54310 73240 54340
rect 73100 54240 73130 54310
rect 73210 54240 73240 54310
rect 73100 54200 73240 54240
rect 73100 54130 73130 54200
rect 73210 54130 73240 54200
rect 73100 54090 73240 54130
rect 73930 54100 73990 55730
rect 74950 55218 76638 56642
rect 76702 55218 76722 56642
rect 77500 55810 77560 57440
rect 78920 57450 78930 57510
rect 78990 57450 79000 57510
rect 78920 57440 79000 57450
rect 77480 55800 77560 55810
rect 78090 56020 78230 56050
rect 78090 55950 78120 56020
rect 78200 55950 78230 56020
rect 78090 55910 78230 55950
rect 78090 55840 78120 55910
rect 78200 55840 78230 55910
rect 78090 55800 78230 55840
rect 78920 55810 78980 57440
rect 78920 55800 79000 55810
rect 77480 55740 77490 55800
rect 77550 55740 77560 55800
rect 77480 55730 77560 55740
rect 74950 55190 76722 55218
rect 74950 54932 76722 54960
rect 73930 54090 74010 54100
rect 72490 54030 72500 54090
rect 72560 54030 72570 54090
rect 72490 54020 72570 54030
rect 69960 53480 71732 53508
rect 69960 53222 71732 53250
rect 69060 52380 69140 52390
rect 69060 52320 69070 52380
rect 69130 52320 69140 52380
rect 69060 52310 69140 52320
rect 69060 50680 69120 52310
rect 69960 51798 71648 53222
rect 71712 51798 71732 53222
rect 72510 52390 72570 54020
rect 73930 54030 73940 54090
rect 74000 54030 74010 54090
rect 73930 54020 74010 54030
rect 72490 52380 72570 52390
rect 73100 52600 73240 52630
rect 73100 52530 73130 52600
rect 73210 52530 73240 52600
rect 73100 52490 73240 52530
rect 73100 52420 73130 52490
rect 73210 52420 73240 52490
rect 73100 52380 73240 52420
rect 73930 52390 73990 54020
rect 74950 53508 76638 54932
rect 76702 53508 76722 54932
rect 77500 54100 77560 55730
rect 78920 55740 78930 55800
rect 78990 55740 79000 55800
rect 78920 55730 79000 55740
rect 77480 54090 77560 54100
rect 78090 54310 78230 54340
rect 78090 54240 78120 54310
rect 78200 54240 78230 54310
rect 78090 54200 78230 54240
rect 78090 54130 78120 54200
rect 78200 54130 78230 54200
rect 78090 54090 78230 54130
rect 78920 54100 78980 55730
rect 78920 54090 79000 54100
rect 77480 54030 77490 54090
rect 77550 54030 77560 54090
rect 77480 54020 77560 54030
rect 74950 53480 76722 53508
rect 74950 53222 76722 53250
rect 73930 52380 74010 52390
rect 72490 52320 72500 52380
rect 72560 52320 72570 52380
rect 72490 52310 72570 52320
rect 69960 51770 71732 51798
rect 69960 51512 71732 51540
rect 69060 50670 69140 50680
rect 69060 50610 69070 50670
rect 69130 50610 69140 50670
rect 69060 50600 69140 50610
rect 69060 48970 69120 50600
rect 69960 50088 71648 51512
rect 71712 50088 71732 51512
rect 72510 50680 72570 52310
rect 73930 52320 73940 52380
rect 74000 52320 74010 52380
rect 73930 52310 74010 52320
rect 72490 50670 72570 50680
rect 73100 50890 73240 50920
rect 73100 50820 73130 50890
rect 73210 50820 73240 50890
rect 73100 50780 73240 50820
rect 73100 50710 73130 50780
rect 73210 50710 73240 50780
rect 73100 50670 73240 50710
rect 73930 50680 73990 52310
rect 74950 51798 76638 53222
rect 76702 51798 76722 53222
rect 77500 52390 77560 54020
rect 78920 54030 78930 54090
rect 78990 54030 79000 54090
rect 78920 54020 79000 54030
rect 77480 52380 77560 52390
rect 78090 52600 78230 52630
rect 78090 52530 78120 52600
rect 78200 52530 78230 52600
rect 78090 52490 78230 52530
rect 78090 52420 78120 52490
rect 78200 52420 78230 52490
rect 78090 52380 78230 52420
rect 78920 52390 78980 54020
rect 78920 52380 79000 52390
rect 77480 52320 77490 52380
rect 77550 52320 77560 52380
rect 77480 52310 77560 52320
rect 74950 51770 76722 51798
rect 74950 51512 76722 51540
rect 73930 50670 74010 50680
rect 72490 50610 72500 50670
rect 72560 50610 72570 50670
rect 72490 50600 72570 50610
rect 69960 50060 71732 50088
rect 69960 49802 71732 49830
rect 69060 48960 69140 48970
rect 69060 48900 69070 48960
rect 69130 48900 69140 48960
rect 69060 48890 69140 48900
rect 69060 47260 69120 48890
rect 69960 48378 71648 49802
rect 71712 48378 71732 49802
rect 72510 48970 72570 50600
rect 73930 50610 73940 50670
rect 74000 50610 74010 50670
rect 73930 50600 74010 50610
rect 72490 48960 72570 48970
rect 73100 49180 73240 49210
rect 73100 49110 73130 49180
rect 73210 49110 73240 49180
rect 73100 49070 73240 49110
rect 73100 49000 73130 49070
rect 73210 49000 73240 49070
rect 73100 48960 73240 49000
rect 73930 48970 73990 50600
rect 74950 50088 76638 51512
rect 76702 50088 76722 51512
rect 77500 50680 77560 52310
rect 78920 52320 78930 52380
rect 78990 52320 79000 52380
rect 78920 52310 79000 52320
rect 77480 50670 77560 50680
rect 78090 50890 78230 50920
rect 78090 50820 78120 50890
rect 78200 50820 78230 50890
rect 78090 50780 78230 50820
rect 78090 50710 78120 50780
rect 78200 50710 78230 50780
rect 78090 50670 78230 50710
rect 78920 50680 78980 52310
rect 78920 50670 79000 50680
rect 77480 50610 77490 50670
rect 77550 50610 77560 50670
rect 77480 50600 77560 50610
rect 74950 50060 76722 50088
rect 74950 49802 76722 49830
rect 73930 48960 74010 48970
rect 72490 48900 72500 48960
rect 72560 48900 72570 48960
rect 72490 48890 72570 48900
rect 69960 48350 71732 48378
rect 69960 48092 71732 48120
rect 69060 47250 69140 47260
rect 69060 47190 69070 47250
rect 69130 47190 69140 47250
rect 69060 47180 69140 47190
rect 69960 46668 71648 48092
rect 71712 46668 71732 48092
rect 72510 47260 72570 48890
rect 73930 48900 73940 48960
rect 74000 48900 74010 48960
rect 73930 48890 74010 48900
rect 72490 47250 72570 47260
rect 73100 47470 73240 47500
rect 73100 47400 73130 47470
rect 73210 47400 73240 47470
rect 73100 47360 73240 47400
rect 73100 47290 73130 47360
rect 73210 47290 73240 47360
rect 73100 47250 73240 47290
rect 73930 47260 73990 48890
rect 74950 48378 76638 49802
rect 76702 48378 76722 49802
rect 77500 48970 77560 50600
rect 78920 50610 78930 50670
rect 78990 50610 79000 50670
rect 78920 50600 79000 50610
rect 77480 48960 77560 48970
rect 78090 49180 78230 49210
rect 78090 49110 78120 49180
rect 78200 49110 78230 49180
rect 78090 49070 78230 49110
rect 78090 49000 78120 49070
rect 78200 49000 78230 49070
rect 78090 48960 78230 49000
rect 78920 48970 78980 50600
rect 78920 48960 79000 48970
rect 77480 48900 77490 48960
rect 77550 48900 77560 48960
rect 77480 48890 77560 48900
rect 74950 48350 76722 48378
rect 74950 48092 76722 48120
rect 73930 47250 74010 47260
rect 72490 47190 72500 47250
rect 72560 47190 72570 47250
rect 72490 47180 72570 47190
rect 69960 46640 71732 46668
rect 69960 46382 71732 46410
rect 68940 45540 69020 45550
rect 67500 45480 67510 45540
rect 67570 45480 67580 45540
rect 67500 45470 67580 45480
rect 64970 44930 66742 44958
rect 64970 44672 66742 44700
rect 63950 43830 64030 43840
rect 62510 43770 62520 43830
rect 62580 43770 62590 43830
rect 62510 43760 62590 43770
rect 59980 43220 61752 43248
rect 59980 42962 61752 42990
rect 58960 42120 59040 42130
rect 57520 42060 57530 42120
rect 57590 42060 57600 42120
rect 57520 42050 57600 42060
rect 54990 41510 56762 41538
rect 54990 41252 56762 41280
rect 53970 40410 54050 40420
rect 52530 40350 52540 40410
rect 52600 40350 52610 40410
rect 52530 40340 52610 40350
rect 53970 40350 53980 40410
rect 54040 40350 54050 40410
rect 53970 40340 54050 40350
rect 50000 39800 51772 39828
rect 54990 39828 56678 41252
rect 56742 39828 56762 41252
rect 57540 40420 57600 42050
rect 58960 42060 58970 42120
rect 59030 42060 59040 42120
rect 58960 42050 59040 42060
rect 57520 40410 57600 40420
rect 58130 40630 58270 40660
rect 58130 40560 58160 40630
rect 58240 40560 58270 40630
rect 58130 40520 58270 40560
rect 58130 40450 58160 40520
rect 58240 40450 58270 40520
rect 58130 40410 58270 40450
rect 58960 40420 59020 42050
rect 59980 41538 61668 42962
rect 61732 41538 61752 42962
rect 62530 42130 62590 43760
rect 63950 43770 63960 43830
rect 64020 43770 64030 43830
rect 63950 43760 64030 43770
rect 62510 42120 62590 42130
rect 63120 42340 63260 42370
rect 63120 42270 63150 42340
rect 63230 42270 63260 42340
rect 63120 42230 63260 42270
rect 63120 42160 63150 42230
rect 63230 42160 63260 42230
rect 63120 42120 63260 42160
rect 63950 42130 64010 43760
rect 64970 43248 66658 44672
rect 66722 43248 66742 44672
rect 67520 43840 67580 45470
rect 68940 45480 68950 45540
rect 69010 45480 69020 45540
rect 68940 45470 69020 45480
rect 67500 43830 67580 43840
rect 68110 44050 68250 44080
rect 68110 43980 68140 44050
rect 68220 43980 68250 44050
rect 68110 43940 68250 43980
rect 68110 43870 68140 43940
rect 68220 43870 68250 43940
rect 68110 43830 68250 43870
rect 68940 43840 69000 45470
rect 69960 44958 71648 46382
rect 71712 44958 71732 46382
rect 72510 45550 72570 47180
rect 73930 47190 73940 47250
rect 74000 47190 74010 47250
rect 73930 47180 74010 47190
rect 72490 45540 72570 45550
rect 73100 45760 73240 45790
rect 73100 45690 73130 45760
rect 73210 45690 73240 45760
rect 73100 45650 73240 45690
rect 73100 45580 73130 45650
rect 73210 45580 73240 45650
rect 73100 45540 73240 45580
rect 73930 45550 73990 47180
rect 74950 46668 76638 48092
rect 76702 46668 76722 48092
rect 77500 47260 77560 48890
rect 78920 48900 78930 48960
rect 78990 48900 79000 48960
rect 78920 48890 79000 48900
rect 77480 47250 77560 47260
rect 78090 47470 78230 47500
rect 78090 47400 78120 47470
rect 78200 47400 78230 47470
rect 78090 47360 78230 47400
rect 78090 47290 78120 47360
rect 78200 47290 78230 47360
rect 78090 47250 78230 47290
rect 78920 47260 78980 48890
rect 78920 47250 79000 47260
rect 77480 47190 77490 47250
rect 77550 47190 77560 47250
rect 77480 47180 77560 47190
rect 74950 46640 76722 46668
rect 74950 46382 76722 46410
rect 73930 45540 74010 45550
rect 72490 45480 72500 45540
rect 72560 45480 72570 45540
rect 72490 45470 72570 45480
rect 69960 44930 71732 44958
rect 69960 44672 71732 44700
rect 68940 43830 69020 43840
rect 67500 43770 67510 43830
rect 67570 43770 67580 43830
rect 67500 43760 67580 43770
rect 64970 43220 66742 43248
rect 64970 42962 66742 42990
rect 63950 42120 64030 42130
rect 62510 42060 62520 42120
rect 62580 42060 62590 42120
rect 62510 42050 62590 42060
rect 59980 41510 61752 41538
rect 59980 41252 61752 41280
rect 58960 40410 59040 40420
rect 57520 40350 57530 40410
rect 57590 40350 57600 40410
rect 57520 40340 57600 40350
rect 58960 40350 58970 40410
rect 59030 40350 59040 40410
rect 58960 40340 59040 40350
rect 54990 39800 56762 39828
rect 59980 39828 61668 41252
rect 61732 39828 61752 41252
rect 62530 40420 62590 42050
rect 63950 42060 63960 42120
rect 64020 42060 64030 42120
rect 63950 42050 64030 42060
rect 62510 40410 62590 40420
rect 63120 40630 63260 40660
rect 63120 40560 63150 40630
rect 63230 40560 63260 40630
rect 63120 40520 63260 40560
rect 63120 40450 63150 40520
rect 63230 40450 63260 40520
rect 63120 40410 63260 40450
rect 63950 40420 64010 42050
rect 64970 41538 66658 42962
rect 66722 41538 66742 42962
rect 67520 42130 67580 43760
rect 68940 43770 68950 43830
rect 69010 43770 69020 43830
rect 68940 43760 69020 43770
rect 67500 42120 67580 42130
rect 68110 42340 68250 42370
rect 68110 42270 68140 42340
rect 68220 42270 68250 42340
rect 68110 42230 68250 42270
rect 68110 42160 68140 42230
rect 68220 42160 68250 42230
rect 68110 42120 68250 42160
rect 68940 42130 69000 43760
rect 69960 43248 71648 44672
rect 71712 43248 71732 44672
rect 72510 43840 72570 45470
rect 73930 45480 73940 45540
rect 74000 45480 74010 45540
rect 73930 45470 74010 45480
rect 72490 43830 72570 43840
rect 73100 44050 73240 44080
rect 73100 43980 73130 44050
rect 73210 43980 73240 44050
rect 73100 43940 73240 43980
rect 73100 43870 73130 43940
rect 73210 43870 73240 43940
rect 73100 43830 73240 43870
rect 73930 43840 73990 45470
rect 74950 44958 76638 46382
rect 76702 44958 76722 46382
rect 77500 45550 77560 47180
rect 78920 47190 78930 47250
rect 78990 47190 79000 47250
rect 78920 47180 79000 47190
rect 77480 45540 77560 45550
rect 78090 45760 78230 45790
rect 78090 45690 78120 45760
rect 78200 45690 78230 45760
rect 78090 45650 78230 45690
rect 78090 45580 78120 45650
rect 78200 45580 78230 45650
rect 78090 45540 78230 45580
rect 78920 45550 78980 47180
rect 78920 45540 79000 45550
rect 77480 45480 77490 45540
rect 77550 45480 77560 45540
rect 77480 45470 77560 45480
rect 74950 44930 76722 44958
rect 74950 44672 76722 44700
rect 73930 43830 74010 43840
rect 72490 43770 72500 43830
rect 72560 43770 72570 43830
rect 72490 43760 72570 43770
rect 69960 43220 71732 43248
rect 69960 42962 71732 42990
rect 68940 42120 69020 42130
rect 67500 42060 67510 42120
rect 67570 42060 67580 42120
rect 67500 42050 67580 42060
rect 64970 41510 66742 41538
rect 64970 41252 66742 41280
rect 63950 40410 64030 40420
rect 62510 40350 62520 40410
rect 62580 40350 62590 40410
rect 62510 40340 62590 40350
rect 63950 40350 63960 40410
rect 64020 40350 64030 40410
rect 63950 40340 64030 40350
rect 59980 39800 61752 39828
rect 64970 39828 66658 41252
rect 66722 39828 66742 41252
rect 67520 40420 67580 42050
rect 68940 42060 68950 42120
rect 69010 42060 69020 42120
rect 68940 42050 69020 42060
rect 67500 40410 67580 40420
rect 68110 40630 68250 40660
rect 68110 40560 68140 40630
rect 68220 40560 68250 40630
rect 68110 40520 68250 40560
rect 68110 40450 68140 40520
rect 68220 40450 68250 40520
rect 68110 40410 68250 40450
rect 68940 40420 69000 42050
rect 69960 41538 71648 42962
rect 71712 41538 71732 42962
rect 72510 42130 72570 43760
rect 73930 43770 73940 43830
rect 74000 43770 74010 43830
rect 73930 43760 74010 43770
rect 72490 42120 72570 42130
rect 73100 42340 73240 42370
rect 73100 42270 73130 42340
rect 73210 42270 73240 42340
rect 73100 42230 73240 42270
rect 73100 42160 73130 42230
rect 73210 42160 73240 42230
rect 73100 42120 73240 42160
rect 73930 42130 73990 43760
rect 74950 43248 76638 44672
rect 76702 43248 76722 44672
rect 77500 43840 77560 45470
rect 78920 45480 78930 45540
rect 78990 45480 79000 45540
rect 78920 45470 79000 45480
rect 77480 43830 77560 43840
rect 78090 44050 78230 44080
rect 78090 43980 78120 44050
rect 78200 43980 78230 44050
rect 78090 43940 78230 43980
rect 78090 43870 78120 43940
rect 78200 43870 78230 43940
rect 78090 43830 78230 43870
rect 78920 43840 78980 45470
rect 78920 43830 79000 43840
rect 77480 43770 77490 43830
rect 77550 43770 77560 43830
rect 77480 43760 77560 43770
rect 74950 43220 76722 43248
rect 74950 42962 76722 42990
rect 73930 42120 74010 42130
rect 72490 42060 72500 42120
rect 72560 42060 72570 42120
rect 72490 42050 72570 42060
rect 69960 41510 71732 41538
rect 69960 41252 71732 41280
rect 68940 40410 69020 40420
rect 67500 40350 67510 40410
rect 67570 40350 67580 40410
rect 67500 40340 67580 40350
rect 68940 40350 68950 40410
rect 69010 40350 69020 40410
rect 68940 40340 69020 40350
rect 64970 39800 66742 39828
rect 69960 39828 71648 41252
rect 71712 39828 71732 41252
rect 72510 40420 72570 42050
rect 73930 42060 73940 42120
rect 74000 42060 74010 42120
rect 73930 42050 74010 42060
rect 72490 40410 72570 40420
rect 73100 40630 73240 40660
rect 73100 40560 73130 40630
rect 73210 40560 73240 40630
rect 73100 40520 73240 40560
rect 73100 40450 73130 40520
rect 73210 40450 73240 40520
rect 73100 40410 73240 40450
rect 73930 40420 73990 42050
rect 74950 41538 76638 42962
rect 76702 41538 76722 42962
rect 77500 42130 77560 43760
rect 78920 43770 78930 43830
rect 78990 43770 79000 43830
rect 78920 43760 79000 43770
rect 77480 42120 77560 42130
rect 78090 42340 78230 42370
rect 78090 42270 78120 42340
rect 78200 42270 78230 42340
rect 78090 42230 78230 42270
rect 78090 42160 78120 42230
rect 78200 42160 78230 42230
rect 78090 42120 78230 42160
rect 78920 42130 78980 43760
rect 78920 42120 79000 42130
rect 77480 42060 77490 42120
rect 77550 42060 77560 42120
rect 77480 42050 77560 42060
rect 74950 41510 76722 41538
rect 74950 41252 76722 41280
rect 73930 40410 74010 40420
rect 72490 40350 72500 40410
rect 72560 40350 72570 40410
rect 72490 40340 72570 40350
rect 73930 40350 73940 40410
rect 74000 40350 74010 40410
rect 73930 40340 74010 40350
rect 69960 39800 71732 39828
rect 74950 39828 76638 41252
rect 76702 39828 76722 41252
rect 77500 40420 77560 42050
rect 78920 42060 78930 42120
rect 78990 42060 79000 42120
rect 78920 42050 79000 42060
rect 77480 40410 77560 40420
rect 78090 40630 78230 40660
rect 78090 40560 78120 40630
rect 78200 40560 78230 40630
rect 78090 40520 78230 40560
rect 78090 40450 78120 40520
rect 78200 40450 78230 40520
rect 78090 40410 78230 40450
rect 78920 40420 78980 42050
rect 78920 40410 79000 40420
rect 77480 40350 77490 40410
rect 77550 40350 77560 40410
rect 77480 40340 77560 40350
rect 78920 40350 78930 40410
rect 78990 40350 79000 40410
rect 78920 40340 79000 40350
rect 74950 39800 76722 39828
rect 40 38830 79800 38840
rect 40 38780 2750 38830
rect 2740 38770 2750 38780
rect 2810 38780 7740 38830
rect 2810 38770 2820 38780
rect 2740 38760 2820 38770
rect 7730 38770 7740 38780
rect 7800 38780 12730 38830
rect 7800 38770 7810 38780
rect 7730 38760 7810 38770
rect 12720 38770 12730 38780
rect 12790 38780 17720 38830
rect 12790 38770 12800 38780
rect 12720 38760 12800 38770
rect 17710 38770 17720 38780
rect 17780 38780 22710 38830
rect 17780 38770 17790 38780
rect 17710 38760 17790 38770
rect 22700 38770 22710 38780
rect 22770 38780 27700 38830
rect 22770 38770 22780 38780
rect 22700 38760 22780 38770
rect 27690 38770 27700 38780
rect 27760 38780 32690 38830
rect 27760 38770 27770 38780
rect 27690 38760 27770 38770
rect 32680 38770 32690 38780
rect 32750 38780 37680 38830
rect 32750 38770 32760 38780
rect 32680 38760 32760 38770
rect 37670 38770 37680 38780
rect 37740 38780 42670 38830
rect 37740 38770 37750 38780
rect 37670 38760 37750 38770
rect 42660 38770 42670 38780
rect 42730 38780 47660 38830
rect 42730 38770 42740 38780
rect 42660 38760 42740 38770
rect 47650 38770 47660 38780
rect 47720 38780 52650 38830
rect 47720 38770 47730 38780
rect 47650 38760 47730 38770
rect 52640 38770 52650 38780
rect 52710 38780 57640 38830
rect 52710 38770 52720 38780
rect 52640 38760 52720 38770
rect 57630 38770 57640 38780
rect 57700 38780 62630 38830
rect 57700 38770 57710 38780
rect 57630 38760 57710 38770
rect 62620 38770 62630 38780
rect 62690 38780 67620 38830
rect 62690 38770 62700 38780
rect 62620 38760 62700 38770
rect 67610 38770 67620 38780
rect 67680 38780 72610 38830
rect 67680 38770 67690 38780
rect 67610 38760 67690 38770
rect 72600 38770 72610 38780
rect 72670 38780 77600 38830
rect 72670 38770 72680 38780
rect 72600 38760 72680 38770
rect 77590 38770 77600 38780
rect 77660 38780 79800 38830
rect 77660 38770 77670 38780
rect 77590 38760 77670 38770
rect 40 38690 79800 38700
rect 40 38640 3820 38690
rect 3810 38630 3820 38640
rect 3880 38640 8810 38690
rect 3880 38630 3890 38640
rect 3810 38620 3890 38630
rect 8800 38630 8810 38640
rect 8870 38640 13800 38690
rect 8870 38630 8880 38640
rect 8800 38620 8880 38630
rect 13790 38630 13800 38640
rect 13860 38640 18790 38690
rect 13860 38630 13870 38640
rect 13790 38620 13870 38630
rect 18780 38630 18790 38640
rect 18850 38640 23780 38690
rect 18850 38630 18860 38640
rect 18780 38620 18860 38630
rect 23770 38630 23780 38640
rect 23840 38640 28770 38690
rect 23840 38630 23850 38640
rect 23770 38620 23850 38630
rect 28760 38630 28770 38640
rect 28830 38640 33760 38690
rect 28830 38630 28840 38640
rect 28760 38620 28840 38630
rect 33750 38630 33760 38640
rect 33820 38640 38750 38690
rect 33820 38630 33830 38640
rect 33750 38620 33830 38630
rect 38740 38630 38750 38640
rect 38810 38640 43740 38690
rect 38810 38630 38820 38640
rect 38740 38620 38820 38630
rect 43730 38630 43740 38640
rect 43800 38640 48730 38690
rect 43800 38630 43810 38640
rect 43730 38620 43810 38630
rect 48720 38630 48730 38640
rect 48790 38640 53720 38690
rect 48790 38630 48800 38640
rect 48720 38620 48800 38630
rect 53710 38630 53720 38640
rect 53780 38640 58710 38690
rect 53780 38630 53790 38640
rect 53710 38620 53790 38630
rect 58700 38630 58710 38640
rect 58770 38640 63700 38690
rect 58770 38630 58780 38640
rect 58700 38620 58780 38630
rect 63690 38630 63700 38640
rect 63760 38640 68690 38690
rect 63760 38630 63770 38640
rect 63690 38620 63770 38630
rect 68680 38630 68690 38640
rect 68750 38640 73680 38690
rect 68750 38630 68760 38640
rect 68680 38620 68760 38630
rect 73670 38630 73680 38640
rect 73740 38640 78670 38690
rect 73740 38630 73750 38640
rect 73670 38620 73750 38630
rect 78660 38630 78670 38640
rect 78730 38640 79800 38690
rect 78730 38630 78740 38640
rect 78660 38620 78740 38630
rect 40 38550 79800 38560
rect 40 38500 36370 38550
rect 36360 38490 36370 38500
rect 36430 38500 79800 38550
rect 36430 38490 36440 38500
rect 36360 38480 36440 38490
rect 40 38410 79800 38420
rect 40 38360 36310 38410
rect 36300 38350 36310 38360
rect 36370 38360 79800 38410
rect 36370 38350 36380 38360
rect 36300 38340 36380 38350
rect 40 38270 79800 38280
rect 40 38220 41540 38270
rect 41530 38210 41540 38220
rect 41600 38220 79800 38270
rect 41600 38210 41610 38220
rect 41530 38200 41610 38210
rect 40 38130 79800 38140
rect 40 38080 41450 38130
rect 41440 38070 41450 38080
rect 41510 38080 79800 38130
rect 41510 38070 41520 38080
rect 41440 38060 41520 38070
rect 40 37990 79800 38000
rect 40 37940 36550 37990
rect 36540 37930 36550 37940
rect 36610 37940 41360 37990
rect 36610 37930 36620 37940
rect 36540 37920 36620 37930
rect 41350 37930 41360 37940
rect 41420 37940 79800 37990
rect 41420 37930 41430 37940
rect 41350 37920 41430 37930
rect 40 37850 79800 37860
rect 40 37800 36490 37850
rect 36480 37790 36490 37800
rect 36550 37800 41300 37850
rect 36550 37790 36560 37800
rect 36480 37780 36560 37790
rect 41290 37790 41300 37800
rect 41360 37800 79800 37850
rect 41360 37790 41370 37800
rect 41290 37780 41370 37790
rect 40 37710 79800 37720
rect 40 37660 31740 37710
rect 31730 37650 31740 37660
rect 31800 37660 46710 37710
rect 31800 37650 31810 37660
rect 31730 37640 31810 37650
rect 46700 37650 46710 37660
rect 46770 37660 79800 37710
rect 46770 37650 46780 37660
rect 46700 37640 46780 37650
rect 40 37570 79800 37580
rect 40 37520 31680 37570
rect 31670 37510 31680 37520
rect 31740 37520 46650 37570
rect 31740 37510 31750 37520
rect 31670 37500 31750 37510
rect 46640 37510 46650 37520
rect 46710 37520 79800 37570
rect 46710 37510 46720 37520
rect 46640 37500 46720 37510
rect 40 37430 79800 37440
rect 40 37380 31560 37430
rect 31550 37370 31560 37380
rect 31620 37380 36730 37430
rect 31620 37370 31630 37380
rect 31550 37360 31630 37370
rect 36720 37370 36730 37380
rect 36790 37380 41720 37430
rect 36790 37370 36800 37380
rect 36720 37360 36800 37370
rect 41710 37370 41720 37380
rect 41780 37380 46530 37430
rect 41780 37370 41790 37380
rect 41710 37360 41790 37370
rect 46520 37370 46530 37380
rect 46590 37380 79800 37430
rect 46590 37370 46600 37380
rect 46520 37360 46600 37370
rect 40 37290 79800 37300
rect 40 37240 31500 37290
rect 31490 37230 31500 37240
rect 31560 37240 36670 37290
rect 31560 37230 31570 37240
rect 31490 37220 31570 37230
rect 36660 37230 36670 37240
rect 36730 37240 41660 37290
rect 36730 37230 36740 37240
rect 36660 37220 36740 37230
rect 41650 37230 41660 37240
rect 41720 37240 46470 37290
rect 41720 37230 41730 37240
rect 41650 37220 41730 37230
rect 46460 37230 46470 37240
rect 46530 37240 79800 37290
rect 46530 37230 46540 37240
rect 46460 37220 46540 37230
rect 40 37150 79800 37160
rect 40 37100 22120 37150
rect 22110 37090 22120 37100
rect 22180 37100 27110 37150
rect 22180 37090 22190 37100
rect 22110 37080 22190 37090
rect 27100 37090 27110 37100
rect 27170 37100 31920 37150
rect 27170 37090 27180 37100
rect 27100 37080 27180 37090
rect 31910 37090 31920 37100
rect 31980 37100 36910 37150
rect 31980 37090 31990 37100
rect 31910 37080 31990 37090
rect 36900 37090 36910 37100
rect 36970 37100 41900 37150
rect 36970 37090 36980 37100
rect 36900 37080 36980 37090
rect 41890 37090 41900 37100
rect 41960 37100 46890 37150
rect 41960 37090 41970 37100
rect 41890 37080 41970 37090
rect 46880 37090 46890 37100
rect 46950 37100 52060 37150
rect 46950 37090 46960 37100
rect 46880 37080 46960 37090
rect 52050 37090 52060 37100
rect 52120 37100 57050 37150
rect 52120 37090 52130 37100
rect 52050 37080 52130 37090
rect 57040 37090 57050 37100
rect 57110 37100 79800 37150
rect 57110 37090 57120 37100
rect 57040 37080 57120 37090
rect 40 37010 79800 37020
rect 40 36960 22060 37010
rect 22050 36950 22060 36960
rect 22120 36960 27050 37010
rect 22120 36950 22130 36960
rect 22050 36940 22130 36950
rect 27040 36950 27050 36960
rect 27110 36960 31860 37010
rect 27110 36950 27120 36960
rect 27040 36940 27120 36950
rect 31850 36950 31860 36960
rect 31920 36960 36850 37010
rect 31920 36950 31930 36960
rect 31850 36940 31930 36950
rect 36840 36950 36850 36960
rect 36910 36960 41840 37010
rect 36910 36950 36920 36960
rect 36840 36940 36920 36950
rect 41830 36950 41840 36960
rect 41900 36960 46830 37010
rect 41900 36950 41910 36960
rect 41830 36940 41910 36950
rect 46820 36950 46830 36960
rect 46890 36960 52000 37010
rect 46890 36950 46900 36960
rect 46820 36940 46900 36950
rect 51990 36950 52000 36960
rect 52060 36960 56990 37010
rect 52060 36950 52070 36960
rect 51990 36940 52070 36950
rect 56980 36950 56990 36960
rect 57050 36960 79800 37010
rect 57050 36950 57060 36960
rect 56980 36940 57060 36950
rect 40 36870 79800 36880
rect 40 36820 21940 36870
rect 21930 36810 21940 36820
rect 22000 36820 26930 36870
rect 22000 36810 22010 36820
rect 21930 36800 22010 36810
rect 26920 36810 26930 36820
rect 26990 36820 32100 36870
rect 26990 36810 27000 36820
rect 26920 36800 27000 36810
rect 32090 36810 32100 36820
rect 32160 36820 37090 36870
rect 32160 36810 32170 36820
rect 32090 36800 32170 36810
rect 37080 36810 37090 36820
rect 37150 36820 42080 36870
rect 37150 36810 37160 36820
rect 37080 36800 37160 36810
rect 42070 36810 42080 36820
rect 42140 36820 47070 36870
rect 42140 36810 42150 36820
rect 42070 36800 42150 36810
rect 47060 36810 47070 36820
rect 47130 36820 51880 36870
rect 47130 36810 47140 36820
rect 47060 36800 47140 36810
rect 51870 36810 51880 36820
rect 51940 36820 56870 36870
rect 51940 36810 51950 36820
rect 51870 36800 51950 36810
rect 56860 36810 56870 36820
rect 56930 36820 79800 36870
rect 56930 36810 56940 36820
rect 56860 36800 56940 36810
rect 40 36730 79800 36740
rect 40 36680 21880 36730
rect 21870 36670 21880 36680
rect 21940 36680 26870 36730
rect 21940 36670 21950 36680
rect 21870 36660 21950 36670
rect 26860 36670 26870 36680
rect 26930 36680 32040 36730
rect 26930 36670 26940 36680
rect 26860 36660 26940 36670
rect 32030 36670 32040 36680
rect 32100 36680 37030 36730
rect 32100 36670 32110 36680
rect 32030 36660 32110 36670
rect 37020 36670 37030 36680
rect 37090 36680 42020 36730
rect 37090 36670 37100 36680
rect 37020 36660 37100 36670
rect 42010 36670 42020 36680
rect 42080 36680 47010 36730
rect 42080 36670 42090 36680
rect 42010 36660 42090 36670
rect 47000 36670 47010 36680
rect 47070 36680 51820 36730
rect 47070 36670 47080 36680
rect 47000 36660 47080 36670
rect 51810 36670 51820 36680
rect 51880 36680 56810 36730
rect 51880 36670 51890 36680
rect 51810 36660 51890 36670
rect 56800 36670 56810 36680
rect 56870 36680 79800 36730
rect 56870 36670 56880 36680
rect 56800 36660 56880 36670
rect 40 36590 79800 36600
rect 40 36540 12320 36590
rect 12310 36530 12320 36540
rect 12380 36540 17310 36590
rect 12380 36530 12390 36540
rect 12310 36520 12390 36530
rect 17300 36530 17310 36540
rect 17370 36540 22300 36590
rect 17370 36530 17380 36540
rect 17300 36520 17380 36530
rect 22290 36530 22300 36540
rect 22360 36540 27290 36590
rect 22360 36530 22370 36540
rect 22290 36520 22370 36530
rect 27280 36530 27290 36540
rect 27350 36540 32280 36590
rect 27350 36530 27360 36540
rect 27280 36520 27360 36530
rect 32270 36530 32280 36540
rect 32340 36540 37270 36590
rect 32340 36530 32350 36540
rect 32270 36520 32350 36530
rect 37260 36530 37270 36540
rect 37330 36540 42260 36590
rect 37330 36530 37340 36540
rect 37260 36520 37340 36530
rect 42250 36530 42260 36540
rect 42320 36540 47250 36590
rect 42320 36530 42330 36540
rect 42250 36520 42330 36530
rect 47240 36530 47250 36540
rect 47310 36540 52240 36590
rect 47310 36530 47320 36540
rect 47240 36520 47320 36530
rect 52230 36530 52240 36540
rect 52300 36540 57230 36590
rect 52300 36530 52310 36540
rect 52230 36520 52310 36530
rect 57220 36530 57230 36540
rect 57290 36540 62220 36590
rect 57290 36530 57300 36540
rect 57220 36520 57300 36530
rect 62210 36530 62220 36540
rect 62280 36540 67210 36590
rect 62280 36530 62290 36540
rect 62210 36520 62290 36530
rect 67200 36530 67210 36540
rect 67270 36540 79800 36590
rect 67270 36530 67280 36540
rect 67200 36520 67280 36530
rect 40 36450 79800 36460
rect 40 36400 12260 36450
rect 12250 36390 12260 36400
rect 12320 36400 17250 36450
rect 12320 36390 12330 36400
rect 12250 36380 12330 36390
rect 17240 36390 17250 36400
rect 17310 36400 22240 36450
rect 17310 36390 17320 36400
rect 17240 36380 17320 36390
rect 22230 36390 22240 36400
rect 22300 36400 27230 36450
rect 22300 36390 22310 36400
rect 22230 36380 22310 36390
rect 27220 36390 27230 36400
rect 27290 36400 32220 36450
rect 27290 36390 27300 36400
rect 27220 36380 27300 36390
rect 32210 36390 32220 36400
rect 32280 36400 37210 36450
rect 32280 36390 32290 36400
rect 32210 36380 32290 36390
rect 37200 36390 37210 36400
rect 37270 36400 42200 36450
rect 37270 36390 37280 36400
rect 37200 36380 37280 36390
rect 42190 36390 42200 36400
rect 42260 36400 47190 36450
rect 42260 36390 42270 36400
rect 42190 36380 42270 36390
rect 47180 36390 47190 36400
rect 47250 36400 52180 36450
rect 47250 36390 47260 36400
rect 47180 36380 47260 36390
rect 52170 36390 52180 36400
rect 52240 36400 57170 36450
rect 52240 36390 52250 36400
rect 52170 36380 52250 36390
rect 57160 36390 57170 36400
rect 57230 36400 62160 36450
rect 57230 36390 57240 36400
rect 57160 36380 57240 36390
rect 62150 36390 62160 36400
rect 62220 36400 67150 36450
rect 62220 36390 62230 36400
rect 62150 36380 62230 36390
rect 67140 36390 67150 36400
rect 67210 36400 79800 36450
rect 67210 36390 67220 36400
rect 67140 36380 67220 36390
rect 40 36310 79800 36320
rect 40 36260 2520 36310
rect 2510 36250 2520 36260
rect 2580 36260 7510 36310
rect 2580 36250 2590 36260
rect 2510 36240 2590 36250
rect 7500 36250 7510 36260
rect 7570 36260 12500 36310
rect 7570 36250 7580 36260
rect 7500 36240 7580 36250
rect 12490 36250 12500 36260
rect 12560 36260 17490 36310
rect 12560 36250 12570 36260
rect 12490 36240 12570 36250
rect 17480 36250 17490 36260
rect 17550 36260 22480 36310
rect 17550 36250 17560 36260
rect 17480 36240 17560 36250
rect 22470 36250 22480 36260
rect 22540 36260 27470 36310
rect 22540 36250 22550 36260
rect 22470 36240 22550 36250
rect 27460 36250 27470 36260
rect 27530 36260 32460 36310
rect 27530 36250 27540 36260
rect 27460 36240 27540 36250
rect 32450 36250 32460 36260
rect 32520 36260 37450 36310
rect 32520 36250 32530 36260
rect 32450 36240 32530 36250
rect 37440 36250 37450 36260
rect 37510 36260 42440 36310
rect 37510 36250 37520 36260
rect 37440 36240 37520 36250
rect 42430 36250 42440 36260
rect 42500 36260 47430 36310
rect 42500 36250 42510 36260
rect 42430 36240 42510 36250
rect 47420 36250 47430 36260
rect 47490 36260 52420 36310
rect 47490 36250 47500 36260
rect 47420 36240 47500 36250
rect 52410 36250 52420 36260
rect 52480 36260 57410 36310
rect 52480 36250 52490 36260
rect 52410 36240 52490 36250
rect 57400 36250 57410 36260
rect 57470 36260 62400 36310
rect 57470 36250 57480 36260
rect 57400 36240 57480 36250
rect 62390 36250 62400 36260
rect 62460 36260 67390 36310
rect 62460 36250 62470 36260
rect 62390 36240 62470 36250
rect 67380 36250 67390 36260
rect 67450 36260 72380 36310
rect 67450 36250 67460 36260
rect 67380 36240 67460 36250
rect 72370 36250 72380 36260
rect 72440 36260 77370 36310
rect 72440 36250 72450 36260
rect 72370 36240 72450 36250
rect 77360 36250 77370 36260
rect 77430 36260 79800 36310
rect 77430 36250 77440 36260
rect 77360 36240 77440 36250
rect 40 36170 79800 36180
rect 40 36120 2460 36170
rect 2450 36110 2460 36120
rect 2520 36120 7450 36170
rect 2520 36110 2530 36120
rect 2450 36100 2530 36110
rect 7440 36110 7450 36120
rect 7510 36120 12440 36170
rect 7510 36110 7520 36120
rect 7440 36100 7520 36110
rect 12430 36110 12440 36120
rect 12500 36120 17430 36170
rect 12500 36110 12510 36120
rect 12430 36100 12510 36110
rect 17420 36110 17430 36120
rect 17490 36120 22420 36170
rect 17490 36110 17500 36120
rect 17420 36100 17500 36110
rect 22410 36110 22420 36120
rect 22480 36120 27410 36170
rect 22480 36110 22490 36120
rect 22410 36100 22490 36110
rect 27400 36110 27410 36120
rect 27470 36120 32400 36170
rect 27470 36110 27480 36120
rect 27400 36100 27480 36110
rect 32390 36110 32400 36120
rect 32460 36120 37390 36170
rect 32460 36110 32470 36120
rect 32390 36100 32470 36110
rect 37380 36110 37390 36120
rect 37450 36120 42380 36170
rect 37450 36110 37460 36120
rect 37380 36100 37460 36110
rect 42370 36110 42380 36120
rect 42440 36120 47370 36170
rect 42440 36110 42450 36120
rect 42370 36100 42450 36110
rect 47360 36110 47370 36120
rect 47430 36120 52360 36170
rect 47430 36110 47440 36120
rect 47360 36100 47440 36110
rect 52350 36110 52360 36120
rect 52420 36120 57350 36170
rect 52420 36110 52430 36120
rect 52350 36100 52430 36110
rect 57340 36110 57350 36120
rect 57410 36120 62340 36170
rect 57410 36110 57420 36120
rect 57340 36100 57420 36110
rect 62330 36110 62340 36120
rect 62400 36120 67330 36170
rect 62400 36110 62410 36120
rect 62330 36100 62410 36110
rect 67320 36110 67330 36120
rect 67390 36120 72320 36170
rect 67390 36110 67400 36120
rect 67320 36100 67400 36110
rect 72310 36110 72320 36120
rect 72380 36120 77310 36170
rect 72380 36110 72390 36120
rect 72310 36100 72390 36110
rect 77300 36110 77310 36120
rect 77370 36120 79800 36170
rect 77370 36110 77380 36120
rect 77300 36100 77380 36110
rect 2350 30940 2430 30950
rect 2350 30930 2360 30940
rect -60 30880 2360 30930
rect 2420 30930 2430 30940
rect 7340 30940 7420 30950
rect 7340 30930 7350 30940
rect 2420 30880 7350 30930
rect 7410 30930 7420 30940
rect 12330 30940 12410 30950
rect 12330 30930 12340 30940
rect 7410 30880 12340 30930
rect 12400 30930 12410 30940
rect 17320 30940 17400 30950
rect 17320 30930 17330 30940
rect 12400 30880 17330 30930
rect 17390 30930 17400 30940
rect 22310 30940 22390 30950
rect 22310 30930 22320 30940
rect 17390 30880 22320 30930
rect 22380 30930 22390 30940
rect 27300 30940 27380 30950
rect 27300 30930 27310 30940
rect 22380 30880 27310 30930
rect 27370 30930 27380 30940
rect 32290 30940 32370 30950
rect 32290 30930 32300 30940
rect 27370 30880 32300 30930
rect 32360 30930 32370 30940
rect 37280 30940 37360 30950
rect 37280 30930 37290 30940
rect 32360 30880 37290 30930
rect 37350 30930 37360 30940
rect 42270 30940 42350 30950
rect 42270 30930 42280 30940
rect 37350 30880 42280 30930
rect 42340 30930 42350 30940
rect 47260 30940 47340 30950
rect 47260 30930 47270 30940
rect 42340 30880 47270 30930
rect 47330 30930 47340 30940
rect 52250 30940 52330 30950
rect 52250 30930 52260 30940
rect 47330 30880 52260 30930
rect 52320 30930 52330 30940
rect 57240 30940 57320 30950
rect 57240 30930 57250 30940
rect 52320 30880 57250 30930
rect 57310 30930 57320 30940
rect 62230 30940 62310 30950
rect 62230 30930 62240 30940
rect 57310 30880 62240 30930
rect 62300 30930 62310 30940
rect 67220 30940 67300 30950
rect 67220 30930 67230 30940
rect 62300 30880 67230 30930
rect 67290 30930 67300 30940
rect 72210 30940 72290 30950
rect 72210 30930 72220 30940
rect 67290 30880 72220 30930
rect 72280 30930 72290 30940
rect 77200 30940 77280 30950
rect 77200 30930 77210 30940
rect 72280 30880 77210 30930
rect 77270 30930 77280 30940
rect 77270 30880 79700 30930
rect -60 30870 79700 30880
rect 2410 30800 2490 30810
rect 2410 30790 2420 30800
rect -60 30740 2420 30790
rect 2480 30790 2490 30800
rect 7400 30800 7480 30810
rect 7400 30790 7410 30800
rect 2480 30740 7410 30790
rect 7470 30790 7480 30800
rect 12390 30800 12470 30810
rect 12390 30790 12400 30800
rect 7470 30740 12400 30790
rect 12460 30790 12470 30800
rect 17380 30800 17460 30810
rect 17380 30790 17390 30800
rect 12460 30740 17390 30790
rect 17450 30790 17460 30800
rect 22370 30800 22450 30810
rect 22370 30790 22380 30800
rect 17450 30740 22380 30790
rect 22440 30790 22450 30800
rect 27360 30800 27440 30810
rect 27360 30790 27370 30800
rect 22440 30740 27370 30790
rect 27430 30790 27440 30800
rect 32350 30800 32430 30810
rect 32350 30790 32360 30800
rect 27430 30740 32360 30790
rect 32420 30790 32430 30800
rect 37340 30800 37420 30810
rect 37340 30790 37350 30800
rect 32420 30740 37350 30790
rect 37410 30790 37420 30800
rect 42330 30800 42410 30810
rect 42330 30790 42340 30800
rect 37410 30740 42340 30790
rect 42400 30790 42410 30800
rect 47320 30800 47400 30810
rect 47320 30790 47330 30800
rect 42400 30740 47330 30790
rect 47390 30790 47400 30800
rect 52310 30800 52390 30810
rect 52310 30790 52320 30800
rect 47390 30740 52320 30790
rect 52380 30790 52390 30800
rect 57300 30800 57380 30810
rect 57300 30790 57310 30800
rect 52380 30740 57310 30790
rect 57370 30790 57380 30800
rect 62290 30800 62370 30810
rect 62290 30790 62300 30800
rect 57370 30740 62300 30790
rect 62360 30790 62370 30800
rect 67280 30800 67360 30810
rect 67280 30790 67290 30800
rect 62360 30740 67290 30790
rect 67350 30790 67360 30800
rect 72270 30800 72350 30810
rect 72270 30790 72280 30800
rect 67350 30740 72280 30790
rect 72340 30790 72350 30800
rect 77260 30800 77340 30810
rect 77260 30790 77270 30800
rect 72340 30740 77270 30790
rect 77330 30790 77340 30800
rect 77330 30740 79700 30790
rect -60 30730 79700 30740
rect 12150 30660 12230 30670
rect 12150 30650 12160 30660
rect -60 30600 12160 30650
rect 12220 30650 12230 30660
rect 17140 30660 17220 30670
rect 17140 30650 17150 30660
rect 12220 30600 17150 30650
rect 17210 30650 17220 30660
rect 22130 30660 22210 30670
rect 22130 30650 22140 30660
rect 17210 30600 22140 30650
rect 22200 30650 22210 30660
rect 27120 30660 27200 30670
rect 27120 30650 27130 30660
rect 22200 30600 27130 30650
rect 27190 30650 27200 30660
rect 32110 30660 32190 30670
rect 32110 30650 32120 30660
rect 27190 30600 32120 30650
rect 32180 30650 32190 30660
rect 37100 30660 37180 30670
rect 37100 30650 37110 30660
rect 32180 30600 37110 30650
rect 37170 30650 37180 30660
rect 42090 30660 42170 30670
rect 42090 30650 42100 30660
rect 37170 30600 42100 30650
rect 42160 30650 42170 30660
rect 47080 30660 47160 30670
rect 47080 30650 47090 30660
rect 42160 30600 47090 30650
rect 47150 30650 47160 30660
rect 52070 30660 52150 30670
rect 52070 30650 52080 30660
rect 47150 30600 52080 30650
rect 52140 30650 52150 30660
rect 57060 30660 57140 30670
rect 57060 30650 57070 30660
rect 52140 30600 57070 30650
rect 57130 30650 57140 30660
rect 62050 30660 62130 30670
rect 62050 30650 62060 30660
rect 57130 30600 62060 30650
rect 62120 30650 62130 30660
rect 67040 30660 67120 30670
rect 67040 30650 67050 30660
rect 62120 30600 67050 30650
rect 67110 30650 67120 30660
rect 67110 30600 79700 30650
rect -60 30590 79700 30600
rect 12210 30520 12290 30530
rect 12210 30510 12220 30520
rect -60 30460 12220 30510
rect 12280 30510 12290 30520
rect 17200 30520 17280 30530
rect 17200 30510 17210 30520
rect 12280 30460 17210 30510
rect 17270 30510 17280 30520
rect 22190 30520 22270 30530
rect 22190 30510 22200 30520
rect 17270 30460 22200 30510
rect 22260 30510 22270 30520
rect 27180 30520 27260 30530
rect 27180 30510 27190 30520
rect 22260 30460 27190 30510
rect 27250 30510 27260 30520
rect 32170 30520 32250 30530
rect 32170 30510 32180 30520
rect 27250 30460 32180 30510
rect 32240 30510 32250 30520
rect 37160 30520 37240 30530
rect 37160 30510 37170 30520
rect 32240 30460 37170 30510
rect 37230 30510 37240 30520
rect 42150 30520 42230 30530
rect 42150 30510 42160 30520
rect 37230 30460 42160 30510
rect 42220 30510 42230 30520
rect 47140 30520 47220 30530
rect 47140 30510 47150 30520
rect 42220 30460 47150 30510
rect 47210 30510 47220 30520
rect 52130 30520 52210 30530
rect 52130 30510 52140 30520
rect 47210 30460 52140 30510
rect 52200 30510 52210 30520
rect 57120 30520 57200 30530
rect 57120 30510 57130 30520
rect 52200 30460 57130 30510
rect 57190 30510 57200 30520
rect 62110 30520 62190 30530
rect 62110 30510 62120 30520
rect 57190 30460 62120 30510
rect 62180 30510 62190 30520
rect 67100 30520 67180 30530
rect 67100 30510 67110 30520
rect 62180 30460 67110 30510
rect 67170 30510 67180 30520
rect 67170 30460 79700 30510
rect -60 30450 79700 30460
rect 21770 30380 21850 30390
rect 21770 30370 21780 30380
rect -60 30320 21780 30370
rect 21840 30370 21850 30380
rect 26760 30380 26840 30390
rect 26760 30370 26770 30380
rect 21840 30320 26770 30370
rect 26830 30370 26840 30380
rect 31930 30380 32010 30390
rect 31930 30370 31940 30380
rect 26830 30320 31940 30370
rect 32000 30370 32010 30380
rect 36920 30380 37000 30390
rect 36920 30370 36930 30380
rect 32000 30320 36930 30370
rect 36990 30370 37000 30380
rect 41910 30380 41990 30390
rect 41910 30370 41920 30380
rect 36990 30320 41920 30370
rect 41980 30370 41990 30380
rect 46900 30380 46980 30390
rect 46900 30370 46910 30380
rect 41980 30320 46910 30370
rect 46970 30370 46980 30380
rect 51710 30380 51790 30390
rect 51710 30370 51720 30380
rect 46970 30320 51720 30370
rect 51780 30370 51790 30380
rect 56700 30380 56780 30390
rect 56700 30370 56710 30380
rect 51780 30320 56710 30370
rect 56770 30370 56780 30380
rect 56770 30320 79700 30370
rect -60 30310 79700 30320
rect 21830 30240 21910 30250
rect 21830 30230 21840 30240
rect -60 30180 21840 30230
rect 21900 30230 21910 30240
rect 26820 30240 26900 30250
rect 26820 30230 26830 30240
rect 21900 30180 26830 30230
rect 26890 30230 26900 30240
rect 31990 30240 32070 30250
rect 31990 30230 32000 30240
rect 26890 30180 32000 30230
rect 32060 30230 32070 30240
rect 36980 30240 37060 30250
rect 36980 30230 36990 30240
rect 32060 30180 36990 30230
rect 37050 30230 37060 30240
rect 41970 30240 42050 30250
rect 41970 30230 41980 30240
rect 37050 30180 41980 30230
rect 42040 30230 42050 30240
rect 46960 30240 47040 30250
rect 46960 30230 46970 30240
rect 42040 30180 46970 30230
rect 47030 30230 47040 30240
rect 51770 30240 51850 30250
rect 51770 30230 51780 30240
rect 47030 30180 51780 30230
rect 51840 30230 51850 30240
rect 56760 30240 56840 30250
rect 56760 30230 56770 30240
rect 51840 30180 56770 30230
rect 56830 30230 56840 30240
rect 56830 30180 79700 30230
rect -60 30170 79700 30180
rect 21950 30100 22030 30110
rect 21950 30090 21960 30100
rect -60 30040 21960 30090
rect 22020 30090 22030 30100
rect 26940 30100 27020 30110
rect 26940 30090 26950 30100
rect 22020 30040 26950 30090
rect 27010 30090 27020 30100
rect 31750 30100 31830 30110
rect 31750 30090 31760 30100
rect 27010 30040 31760 30090
rect 31820 30090 31830 30100
rect 36740 30100 36820 30110
rect 36740 30090 36750 30100
rect 31820 30040 36750 30090
rect 36810 30090 36820 30100
rect 41730 30100 41810 30110
rect 41730 30090 41740 30100
rect 36810 30040 41740 30090
rect 41800 30090 41810 30100
rect 46720 30100 46800 30110
rect 46720 30090 46730 30100
rect 41800 30040 46730 30090
rect 46790 30090 46800 30100
rect 51890 30100 51970 30110
rect 51890 30090 51900 30100
rect 46790 30040 51900 30090
rect 51960 30090 51970 30100
rect 56880 30100 56960 30110
rect 56880 30090 56890 30100
rect 51960 30040 56890 30090
rect 56950 30090 56960 30100
rect 56950 30040 79700 30090
rect -60 30030 79700 30040
rect 22010 29960 22090 29970
rect 22010 29950 22020 29960
rect -60 29900 22020 29950
rect 22080 29950 22090 29960
rect 27000 29960 27080 29970
rect 27000 29950 27010 29960
rect 22080 29900 27010 29950
rect 27070 29950 27080 29960
rect 31810 29960 31890 29970
rect 31810 29950 31820 29960
rect 27070 29900 31820 29950
rect 31880 29950 31890 29960
rect 36800 29960 36880 29970
rect 36800 29950 36810 29960
rect 31880 29900 36810 29950
rect 36870 29950 36880 29960
rect 41790 29960 41870 29970
rect 41790 29950 41800 29960
rect 36870 29900 41800 29950
rect 41860 29950 41870 29960
rect 46780 29960 46860 29970
rect 46780 29950 46790 29960
rect 41860 29900 46790 29950
rect 46850 29950 46860 29960
rect 51950 29960 52030 29970
rect 51950 29950 51960 29960
rect 46850 29900 51960 29950
rect 52020 29950 52030 29960
rect 56940 29960 57020 29970
rect 56940 29950 56950 29960
rect 52020 29900 56950 29950
rect 57010 29950 57020 29960
rect 57010 29900 79700 29950
rect -60 29890 79700 29900
rect 31390 29820 31470 29830
rect 31390 29810 31400 29820
rect -60 29760 31400 29810
rect 31460 29810 31470 29820
rect 36560 29820 36640 29830
rect 36560 29810 36570 29820
rect 31460 29760 36570 29810
rect 36630 29810 36640 29820
rect 41550 29820 41630 29830
rect 41550 29810 41560 29820
rect 36630 29760 41560 29810
rect 41620 29810 41630 29820
rect 46360 29820 46440 29830
rect 46360 29810 46370 29820
rect 41620 29760 46370 29810
rect 46430 29810 46440 29820
rect 46430 29760 79700 29810
rect -60 29750 79700 29760
rect 31450 29680 31530 29690
rect 31450 29670 31460 29680
rect -60 29620 31460 29670
rect 31520 29670 31530 29680
rect 36620 29680 36700 29690
rect 36620 29670 36630 29680
rect 31520 29620 36630 29670
rect 36690 29670 36700 29680
rect 41610 29680 41690 29690
rect 41610 29670 41620 29680
rect 36690 29620 41620 29670
rect 41680 29670 41690 29680
rect 46420 29680 46500 29690
rect 46420 29670 46430 29680
rect 41680 29620 46430 29670
rect 46490 29670 46500 29680
rect 46490 29620 79700 29670
rect -60 29610 79700 29620
rect 31570 29540 31650 29550
rect 31570 29530 31580 29540
rect -60 29480 31580 29530
rect 31640 29530 31650 29540
rect 46540 29540 46620 29550
rect 46540 29530 46550 29540
rect 31640 29480 46550 29530
rect 46610 29530 46620 29540
rect 46610 29480 79700 29530
rect -60 29470 79700 29480
rect 31630 29400 31710 29410
rect 31630 29390 31640 29400
rect -60 29340 31640 29390
rect 31700 29390 31710 29400
rect 46600 29400 46680 29410
rect 46600 29390 46610 29400
rect 31700 29340 46610 29390
rect 46670 29390 46680 29400
rect 46670 29340 79700 29390
rect -60 29330 79700 29340
rect 36380 29260 36460 29270
rect 36380 29250 36390 29260
rect -60 29200 36390 29250
rect 36450 29250 36460 29260
rect 41190 29260 41270 29270
rect 41190 29250 41200 29260
rect 36450 29200 41200 29250
rect 41260 29250 41270 29260
rect 41260 29200 79700 29250
rect -60 29190 79700 29200
rect 36440 29120 36520 29130
rect 36440 29110 36450 29120
rect -60 29060 36450 29110
rect 36510 29110 36520 29120
rect 41250 29120 41330 29130
rect 41250 29110 41260 29120
rect 36510 29060 41260 29110
rect 41320 29110 41330 29120
rect 41320 29060 79700 29110
rect -60 29050 79700 29060
rect 41340 28980 41420 28990
rect 41340 28970 41350 28980
rect -60 28920 41350 28970
rect 41410 28970 41420 28980
rect 41410 28920 79700 28970
rect -60 28910 79700 28920
rect 41430 28840 41510 28850
rect 41430 28830 41440 28840
rect -60 28780 41440 28830
rect 41500 28830 41510 28840
rect 41500 28780 79700 28830
rect -60 28770 79700 28780
rect 36200 28700 36280 28710
rect 36200 28690 36210 28700
rect -60 28640 36210 28690
rect 36270 28690 36280 28700
rect 36270 28640 79700 28690
rect -60 28630 79700 28640
rect 36260 28560 36340 28570
rect 36260 28550 36270 28560
rect -60 28500 36270 28550
rect 36330 28550 36340 28560
rect 36330 28500 79700 28550
rect -60 28490 79700 28500
rect 3710 28420 3790 28430
rect 3710 28410 3720 28420
rect -60 28360 3720 28410
rect 3780 28410 3790 28420
rect 8700 28420 8780 28430
rect 8700 28410 8710 28420
rect 3780 28360 8710 28410
rect 8770 28410 8780 28420
rect 13690 28420 13770 28430
rect 13690 28410 13700 28420
rect 8770 28360 13700 28410
rect 13760 28410 13770 28420
rect 18680 28420 18760 28430
rect 18680 28410 18690 28420
rect 13760 28360 18690 28410
rect 18750 28410 18760 28420
rect 23670 28420 23750 28430
rect 23670 28410 23680 28420
rect 18750 28360 23680 28410
rect 23740 28410 23750 28420
rect 28660 28420 28740 28430
rect 28660 28410 28670 28420
rect 23740 28360 28670 28410
rect 28730 28410 28740 28420
rect 33650 28420 33730 28430
rect 33650 28410 33660 28420
rect 28730 28360 33660 28410
rect 33720 28410 33730 28420
rect 38640 28420 38720 28430
rect 38640 28410 38650 28420
rect 33720 28360 38650 28410
rect 38710 28410 38720 28420
rect 43630 28420 43710 28430
rect 43630 28410 43640 28420
rect 38710 28360 43640 28410
rect 43700 28410 43710 28420
rect 48620 28420 48700 28430
rect 48620 28410 48630 28420
rect 43700 28360 48630 28410
rect 48690 28410 48700 28420
rect 53610 28420 53690 28430
rect 53610 28410 53620 28420
rect 48690 28360 53620 28410
rect 53680 28410 53690 28420
rect 58600 28420 58680 28430
rect 58600 28410 58610 28420
rect 53680 28360 58610 28410
rect 58670 28410 58680 28420
rect 63590 28420 63670 28430
rect 63590 28410 63600 28420
rect 58670 28360 63600 28410
rect 63660 28410 63670 28420
rect 68580 28420 68660 28430
rect 68580 28410 68590 28420
rect 63660 28360 68590 28410
rect 68650 28410 68660 28420
rect 73570 28420 73650 28430
rect 73570 28410 73580 28420
rect 68650 28360 73580 28410
rect 73640 28410 73650 28420
rect 78560 28420 78640 28430
rect 78560 28410 78570 28420
rect 73640 28360 78570 28410
rect 78630 28410 78640 28420
rect 78630 28360 79700 28410
rect -60 28350 79700 28360
rect 2640 28280 2720 28290
rect 2640 28270 2650 28280
rect -60 28220 2650 28270
rect 2710 28270 2720 28280
rect 7630 28280 7710 28290
rect 7630 28270 7640 28280
rect 2710 28220 7640 28270
rect 7700 28270 7710 28280
rect 12620 28280 12700 28290
rect 12620 28270 12630 28280
rect 7700 28220 12630 28270
rect 12690 28270 12700 28280
rect 17610 28280 17690 28290
rect 17610 28270 17620 28280
rect 12690 28220 17620 28270
rect 17680 28270 17690 28280
rect 22600 28280 22680 28290
rect 22600 28270 22610 28280
rect 17680 28220 22610 28270
rect 22670 28270 22680 28280
rect 27590 28280 27670 28290
rect 27590 28270 27600 28280
rect 22670 28220 27600 28270
rect 27660 28270 27670 28280
rect 32580 28280 32660 28290
rect 32580 28270 32590 28280
rect 27660 28220 32590 28270
rect 32650 28270 32660 28280
rect 37570 28280 37650 28290
rect 37570 28270 37580 28280
rect 32650 28220 37580 28270
rect 37640 28270 37650 28280
rect 42560 28280 42640 28290
rect 42560 28270 42570 28280
rect 37640 28220 42570 28270
rect 42630 28270 42640 28280
rect 47550 28280 47630 28290
rect 47550 28270 47560 28280
rect 42630 28220 47560 28270
rect 47620 28270 47630 28280
rect 52540 28280 52620 28290
rect 52540 28270 52550 28280
rect 47620 28220 52550 28270
rect 52610 28270 52620 28280
rect 57530 28280 57610 28290
rect 57530 28270 57540 28280
rect 52610 28220 57540 28270
rect 57600 28270 57610 28280
rect 62520 28280 62600 28290
rect 62520 28270 62530 28280
rect 57600 28220 62530 28270
rect 62590 28270 62600 28280
rect 67510 28280 67590 28290
rect 67510 28270 67520 28280
rect 62590 28220 67520 28270
rect 67580 28270 67590 28280
rect 72500 28280 72580 28290
rect 72500 28270 72510 28280
rect 67580 28220 72510 28270
rect 72570 28270 72580 28280
rect 77490 28280 77570 28290
rect 77490 28270 77500 28280
rect 72570 28220 77500 28270
rect 77560 28270 77570 28280
rect 77560 28220 79700 28270
rect -60 28210 79700 28220
<< via3 >>
rect 1788 65478 1852 66902
rect 3270 66210 3280 66280
rect 3280 66210 3350 66280
rect 3270 66100 3280 66170
rect 3280 66100 3350 66170
rect 1788 63768 1852 65192
rect 3270 64500 3280 64570
rect 3280 64500 3350 64570
rect 3270 64390 3280 64460
rect 3280 64390 3350 64460
rect 6778 65478 6842 66902
rect 8260 66210 8270 66280
rect 8270 66210 8340 66280
rect 8260 66100 8270 66170
rect 8270 66100 8340 66170
rect 1788 62058 1852 63482
rect 3270 62790 3280 62860
rect 3280 62790 3350 62860
rect 3270 62680 3280 62750
rect 3280 62680 3350 62750
rect 6778 63768 6842 65192
rect 8260 64500 8270 64570
rect 8270 64500 8340 64570
rect 8260 64390 8270 64460
rect 8270 64390 8340 64460
rect 11768 65478 11832 66902
rect 13250 66210 13260 66280
rect 13260 66210 13330 66280
rect 13250 66100 13260 66170
rect 13260 66100 13330 66170
rect 1788 60348 1852 61772
rect 3270 61080 3280 61150
rect 3280 61080 3350 61150
rect 3270 60970 3280 61040
rect 3280 60970 3350 61040
rect 6778 62058 6842 63482
rect 8260 62790 8270 62860
rect 8270 62790 8340 62860
rect 8260 62680 8270 62750
rect 8270 62680 8340 62750
rect 11768 63768 11832 65192
rect 13250 64500 13260 64570
rect 13260 64500 13330 64570
rect 13250 64390 13260 64460
rect 13260 64390 13330 64460
rect 16758 65478 16822 66902
rect 18240 66210 18250 66280
rect 18250 66210 18320 66280
rect 18240 66100 18250 66170
rect 18250 66100 18320 66170
rect 1788 58638 1852 60062
rect 3270 59370 3280 59440
rect 3280 59370 3350 59440
rect 3270 59260 3280 59330
rect 3280 59260 3350 59330
rect 6778 60348 6842 61772
rect 8260 61080 8270 61150
rect 8270 61080 8340 61150
rect 8260 60970 8270 61040
rect 8270 60970 8340 61040
rect 11768 62058 11832 63482
rect 13250 62790 13260 62860
rect 13260 62790 13330 62860
rect 13250 62680 13260 62750
rect 13260 62680 13330 62750
rect 16758 63768 16822 65192
rect 18240 64500 18250 64570
rect 18250 64500 18320 64570
rect 18240 64390 18250 64460
rect 18250 64390 18320 64460
rect 21748 65478 21812 66902
rect 23230 66210 23240 66280
rect 23240 66210 23310 66280
rect 23230 66100 23240 66170
rect 23240 66100 23310 66170
rect 1788 56928 1852 58352
rect 3270 57660 3280 57730
rect 3280 57660 3350 57730
rect 3270 57550 3280 57620
rect 3280 57550 3350 57620
rect 6778 58638 6842 60062
rect 8260 59370 8270 59440
rect 8270 59370 8340 59440
rect 8260 59260 8270 59330
rect 8270 59260 8340 59330
rect 11768 60348 11832 61772
rect 13250 61080 13260 61150
rect 13260 61080 13330 61150
rect 13250 60970 13260 61040
rect 13260 60970 13330 61040
rect 16758 62058 16822 63482
rect 18240 62790 18250 62860
rect 18250 62790 18320 62860
rect 18240 62680 18250 62750
rect 18250 62680 18320 62750
rect 21748 63768 21812 65192
rect 23230 64500 23240 64570
rect 23240 64500 23310 64570
rect 23230 64390 23240 64460
rect 23240 64390 23310 64460
rect 26738 65478 26802 66902
rect 28220 66210 28230 66280
rect 28230 66210 28300 66280
rect 28220 66100 28230 66170
rect 28230 66100 28300 66170
rect 1788 55218 1852 56642
rect 3270 55950 3280 56020
rect 3280 55950 3350 56020
rect 3270 55840 3280 55910
rect 3280 55840 3350 55910
rect 6778 56928 6842 58352
rect 8260 57660 8270 57730
rect 8270 57660 8340 57730
rect 8260 57550 8270 57620
rect 8270 57550 8340 57620
rect 11768 58638 11832 60062
rect 1788 53508 1852 54932
rect 3270 54240 3280 54310
rect 3280 54240 3350 54310
rect 3270 54130 3280 54200
rect 3280 54130 3350 54200
rect 6778 55218 6842 56642
rect 8260 55950 8270 56020
rect 8270 55950 8340 56020
rect 8260 55840 8270 55910
rect 8270 55840 8340 55910
rect 11768 56928 11832 58352
rect 1788 51798 1852 53222
rect 3270 52530 3280 52600
rect 3280 52530 3350 52600
rect 3270 52420 3280 52490
rect 3280 52420 3350 52490
rect 6778 53508 6842 54932
rect 8260 54240 8270 54310
rect 8270 54240 8340 54310
rect 8260 54130 8270 54200
rect 8270 54130 8340 54200
rect 11768 55218 11832 56642
rect 1788 50088 1852 51512
rect 3270 50820 3280 50890
rect 3280 50820 3350 50890
rect 3270 50710 3280 50780
rect 3280 50710 3350 50780
rect 6778 51798 6842 53222
rect 8260 52530 8270 52600
rect 8270 52530 8340 52600
rect 8260 52420 8270 52490
rect 8270 52420 8340 52490
rect 11768 53508 11832 54932
rect 1788 48378 1852 49802
rect 3270 49110 3280 49180
rect 3280 49110 3350 49180
rect 3270 49000 3280 49070
rect 3280 49000 3350 49070
rect 6778 50088 6842 51512
rect 8260 50820 8270 50890
rect 8270 50820 8340 50890
rect 8260 50710 8270 50780
rect 8270 50710 8340 50780
rect 11768 51798 11832 53222
rect 1788 46668 1852 48092
rect 3270 47400 3280 47470
rect 3280 47400 3350 47470
rect 3270 47290 3280 47360
rect 3280 47290 3350 47360
rect 6778 48378 6842 49802
rect 8260 49110 8270 49180
rect 8270 49110 8340 49180
rect 8260 49000 8270 49070
rect 8270 49000 8340 49070
rect 11768 50088 11832 51512
rect 1788 44958 1852 46382
rect 3270 45690 3280 45760
rect 3280 45690 3350 45760
rect 3270 45580 3280 45650
rect 3280 45580 3350 45650
rect 6778 46668 6842 48092
rect 8260 47400 8270 47470
rect 8270 47400 8340 47470
rect 8260 47290 8270 47360
rect 8270 47290 8340 47360
rect 11768 48378 11832 49802
rect 1788 43248 1852 44672
rect 3270 43980 3280 44050
rect 3280 43980 3350 44050
rect 3270 43870 3280 43940
rect 3280 43870 3350 43940
rect 6778 44958 6842 46382
rect 8260 45690 8270 45760
rect 8270 45690 8340 45760
rect 8260 45580 8270 45650
rect 8270 45580 8340 45650
rect 11768 46668 11832 48092
rect 1788 41538 1852 42962
rect 3270 42270 3280 42340
rect 3280 42270 3350 42340
rect 3270 42160 3280 42230
rect 3280 42160 3350 42230
rect 6778 43248 6842 44672
rect 8260 43980 8270 44050
rect 8270 43980 8340 44050
rect 8260 43870 8270 43940
rect 8270 43870 8340 43940
rect 11768 44958 11832 46382
rect 13250 59370 13260 59440
rect 13260 59370 13330 59440
rect 13250 59260 13260 59330
rect 13260 59260 13330 59330
rect 13250 57660 13260 57730
rect 13260 57660 13330 57730
rect 13250 57550 13260 57620
rect 13260 57550 13330 57620
rect 13250 55950 13260 56020
rect 13260 55950 13330 56020
rect 13250 55840 13260 55910
rect 13260 55840 13330 55910
rect 13250 54240 13260 54310
rect 13260 54240 13330 54310
rect 13250 54130 13260 54200
rect 13260 54130 13330 54200
rect 13250 52530 13260 52600
rect 13260 52530 13330 52600
rect 13250 52420 13260 52490
rect 13260 52420 13330 52490
rect 13250 50820 13260 50890
rect 13260 50820 13330 50890
rect 13250 50710 13260 50780
rect 13260 50710 13330 50780
rect 13250 49110 13260 49180
rect 13260 49110 13330 49180
rect 13250 49000 13260 49070
rect 13260 49000 13330 49070
rect 13250 47400 13260 47470
rect 13260 47400 13330 47470
rect 13250 47290 13260 47360
rect 13260 47290 13330 47360
rect 13250 45690 13260 45760
rect 13260 45690 13330 45760
rect 13250 45580 13260 45650
rect 13260 45580 13330 45650
rect 16758 60348 16822 61772
rect 18240 61080 18250 61150
rect 18250 61080 18320 61150
rect 18240 60970 18250 61040
rect 18250 60970 18320 61040
rect 21748 62058 21812 63482
rect 16758 58638 16822 60062
rect 16758 56928 16822 58352
rect 16758 55218 16822 56642
rect 16758 53508 16822 54932
rect 16758 51798 16822 53222
rect 16758 50088 16822 51512
rect 16758 48378 16822 49802
rect 16758 46668 16822 48092
rect 1788 39828 1852 41252
rect 3270 40560 3280 40630
rect 3280 40560 3350 40630
rect 3270 40450 3280 40520
rect 3280 40450 3350 40520
rect 6778 41538 6842 42962
rect 8260 42270 8270 42340
rect 8270 42270 8340 42340
rect 8260 42160 8270 42230
rect 8270 42160 8340 42230
rect 11768 43248 11832 44672
rect 13250 43980 13260 44050
rect 13260 43980 13330 44050
rect 13250 43870 13260 43940
rect 13260 43870 13330 43940
rect 16758 44958 16822 46382
rect 18240 59370 18250 59440
rect 18250 59370 18320 59440
rect 18240 59260 18250 59330
rect 18250 59260 18320 59330
rect 18240 57660 18250 57730
rect 18250 57660 18320 57730
rect 18240 57550 18250 57620
rect 18250 57550 18320 57620
rect 18240 55950 18250 56020
rect 18250 55950 18320 56020
rect 18240 55840 18250 55910
rect 18250 55840 18320 55910
rect 18240 54240 18250 54310
rect 18250 54240 18320 54310
rect 18240 54130 18250 54200
rect 18250 54130 18320 54200
rect 18240 52530 18250 52600
rect 18250 52530 18320 52600
rect 18240 52420 18250 52490
rect 18250 52420 18320 52490
rect 18240 50820 18250 50890
rect 18250 50820 18320 50890
rect 18240 50710 18250 50780
rect 18250 50710 18320 50780
rect 18240 49110 18250 49180
rect 18250 49110 18320 49180
rect 18240 49000 18250 49070
rect 18250 49000 18320 49070
rect 18240 47400 18250 47470
rect 18250 47400 18320 47470
rect 18240 47290 18250 47360
rect 18250 47290 18320 47360
rect 18240 45690 18250 45760
rect 18250 45690 18320 45760
rect 18240 45580 18250 45650
rect 18250 45580 18320 45650
rect 21748 60348 21812 61772
rect 21748 58638 21812 60062
rect 21748 56928 21812 58352
rect 21748 55218 21812 56642
rect 21748 53508 21812 54932
rect 21748 51798 21812 53222
rect 21748 50088 21812 51512
rect 21748 48378 21812 49802
rect 21748 46668 21812 48092
rect 6778 39828 6842 41252
rect 8260 40560 8270 40630
rect 8270 40560 8340 40630
rect 8260 40450 8270 40520
rect 8270 40450 8340 40520
rect 11768 41538 11832 42962
rect 13250 42270 13260 42340
rect 13260 42270 13330 42340
rect 13250 42160 13260 42230
rect 13260 42160 13330 42230
rect 16758 43248 16822 44672
rect 18240 43980 18250 44050
rect 18250 43980 18320 44050
rect 18240 43870 18250 43940
rect 18250 43870 18320 43940
rect 21748 44958 21812 46382
rect 11768 39828 11832 41252
rect 13250 40560 13260 40630
rect 13260 40560 13330 40630
rect 13250 40450 13260 40520
rect 13260 40450 13330 40520
rect 16758 41538 16822 42962
rect 18240 42270 18250 42340
rect 18250 42270 18320 42340
rect 18240 42160 18250 42230
rect 18250 42160 18320 42230
rect 21748 43248 21812 44672
rect 16758 39828 16822 41252
rect 18240 40560 18250 40630
rect 18250 40560 18320 40630
rect 18240 40450 18250 40520
rect 18250 40450 18320 40520
rect 21748 41538 21812 42962
rect 23230 62790 23240 62860
rect 23240 62790 23310 62860
rect 23230 62680 23240 62750
rect 23240 62680 23310 62750
rect 23230 61080 23240 61150
rect 23240 61080 23310 61150
rect 23230 60970 23240 61040
rect 23240 60970 23310 61040
rect 23230 59370 23240 59440
rect 23240 59370 23310 59440
rect 23230 59260 23240 59330
rect 23240 59260 23310 59330
rect 23230 57660 23240 57730
rect 23240 57660 23310 57730
rect 23230 57550 23240 57620
rect 23240 57550 23310 57620
rect 23230 55950 23240 56020
rect 23240 55950 23310 56020
rect 23230 55840 23240 55910
rect 23240 55840 23310 55910
rect 23230 54240 23240 54310
rect 23240 54240 23310 54310
rect 23230 54130 23240 54200
rect 23240 54130 23310 54200
rect 23230 52530 23240 52600
rect 23240 52530 23310 52600
rect 23230 52420 23240 52490
rect 23240 52420 23310 52490
rect 23230 50820 23240 50890
rect 23240 50820 23310 50890
rect 23230 50710 23240 50780
rect 23240 50710 23310 50780
rect 23230 49110 23240 49180
rect 23240 49110 23310 49180
rect 23230 49000 23240 49070
rect 23240 49000 23310 49070
rect 23230 47400 23240 47470
rect 23240 47400 23310 47470
rect 23230 47290 23240 47360
rect 23240 47290 23310 47360
rect 23230 45690 23240 45760
rect 23240 45690 23310 45760
rect 23230 45580 23240 45650
rect 23240 45580 23310 45650
rect 23230 43980 23240 44050
rect 23240 43980 23310 44050
rect 23230 43870 23240 43940
rect 23240 43870 23310 43940
rect 23230 42270 23240 42340
rect 23240 42270 23310 42340
rect 23230 42160 23240 42230
rect 23240 42160 23310 42230
rect 26738 63768 26802 65192
rect 28220 64500 28230 64570
rect 28230 64500 28300 64570
rect 28220 64390 28230 64460
rect 28230 64390 28300 64460
rect 31728 65478 31792 66902
rect 33210 66210 33220 66280
rect 33220 66210 33290 66280
rect 33210 66100 33220 66170
rect 33220 66100 33290 66170
rect 26738 62058 26802 63482
rect 26738 60348 26802 61772
rect 26738 58638 26802 60062
rect 26738 56928 26802 58352
rect 26738 55218 26802 56642
rect 26738 53508 26802 54932
rect 26738 51798 26802 53222
rect 26738 50088 26802 51512
rect 26738 48378 26802 49802
rect 26738 46668 26802 48092
rect 26738 44958 26802 46382
rect 26738 43248 26802 44672
rect 21748 39828 21812 41252
rect 23230 40560 23240 40630
rect 23240 40560 23310 40630
rect 23230 40450 23240 40520
rect 23240 40450 23310 40520
rect 26738 41538 26802 42962
rect 28220 62790 28230 62860
rect 28230 62790 28300 62860
rect 28220 62680 28230 62750
rect 28230 62680 28300 62750
rect 28220 61080 28230 61150
rect 28230 61080 28300 61150
rect 28220 60970 28230 61040
rect 28230 60970 28300 61040
rect 28220 59370 28230 59440
rect 28230 59370 28300 59440
rect 28220 59260 28230 59330
rect 28230 59260 28300 59330
rect 28220 57660 28230 57730
rect 28230 57660 28300 57730
rect 28220 57550 28230 57620
rect 28230 57550 28300 57620
rect 28220 55950 28230 56020
rect 28230 55950 28300 56020
rect 28220 55840 28230 55910
rect 28230 55840 28300 55910
rect 28220 54240 28230 54310
rect 28230 54240 28300 54310
rect 28220 54130 28230 54200
rect 28230 54130 28300 54200
rect 28220 52530 28230 52600
rect 28230 52530 28300 52600
rect 28220 52420 28230 52490
rect 28230 52420 28300 52490
rect 28220 50820 28230 50890
rect 28230 50820 28300 50890
rect 28220 50710 28230 50780
rect 28230 50710 28300 50780
rect 28220 49110 28230 49180
rect 28230 49110 28300 49180
rect 28220 49000 28230 49070
rect 28230 49000 28300 49070
rect 28220 47400 28230 47470
rect 28230 47400 28300 47470
rect 28220 47290 28230 47360
rect 28230 47290 28300 47360
rect 28220 45690 28230 45760
rect 28230 45690 28300 45760
rect 28220 45580 28230 45650
rect 28230 45580 28300 45650
rect 28220 43980 28230 44050
rect 28230 43980 28300 44050
rect 28220 43870 28230 43940
rect 28230 43870 28300 43940
rect 28220 42270 28230 42340
rect 28230 42270 28300 42340
rect 28220 42160 28230 42230
rect 28230 42160 28300 42230
rect 31728 63768 31792 65192
rect 33210 64500 33220 64570
rect 33220 64500 33290 64570
rect 33210 64390 33220 64460
rect 33220 64390 33290 64460
rect 36718 65478 36782 66902
rect 38200 66210 38210 66280
rect 38210 66210 38280 66280
rect 38200 66100 38210 66170
rect 38210 66100 38280 66170
rect 31728 62058 31792 63482
rect 31728 60348 31792 61772
rect 31728 58638 31792 60062
rect 31728 56928 31792 58352
rect 31728 55218 31792 56642
rect 31728 53508 31792 54932
rect 31728 51798 31792 53222
rect 31728 50088 31792 51512
rect 31728 48378 31792 49802
rect 31728 46668 31792 48092
rect 31728 44958 31792 46382
rect 31728 43248 31792 44672
rect 26738 39828 26802 41252
rect 28220 40560 28230 40630
rect 28230 40560 28300 40630
rect 28220 40450 28230 40520
rect 28230 40450 28300 40520
rect 31728 41538 31792 42962
rect 33210 62790 33220 62860
rect 33220 62790 33290 62860
rect 33210 62680 33220 62750
rect 33220 62680 33290 62750
rect 33210 61080 33220 61150
rect 33220 61080 33290 61150
rect 33210 60970 33220 61040
rect 33220 60970 33290 61040
rect 33210 59370 33220 59440
rect 33220 59370 33290 59440
rect 33210 59260 33220 59330
rect 33220 59260 33290 59330
rect 33210 57660 33220 57730
rect 33220 57660 33290 57730
rect 33210 57550 33220 57620
rect 33220 57550 33290 57620
rect 33210 55950 33220 56020
rect 33220 55950 33290 56020
rect 33210 55840 33220 55910
rect 33220 55840 33290 55910
rect 33210 54240 33220 54310
rect 33220 54240 33290 54310
rect 33210 54130 33220 54200
rect 33220 54130 33290 54200
rect 33210 52530 33220 52600
rect 33220 52530 33290 52600
rect 33210 52420 33220 52490
rect 33220 52420 33290 52490
rect 33210 50820 33220 50890
rect 33220 50820 33290 50890
rect 33210 50710 33220 50780
rect 33220 50710 33290 50780
rect 33210 49110 33220 49180
rect 33220 49110 33290 49180
rect 33210 49000 33220 49070
rect 33220 49000 33290 49070
rect 33210 47400 33220 47470
rect 33220 47400 33290 47470
rect 33210 47290 33220 47360
rect 33220 47290 33290 47360
rect 33210 45690 33220 45760
rect 33220 45690 33290 45760
rect 33210 45580 33220 45650
rect 33220 45580 33290 45650
rect 33210 43980 33220 44050
rect 33220 43980 33290 44050
rect 33210 43870 33220 43940
rect 33220 43870 33290 43940
rect 33210 42270 33220 42340
rect 33220 42270 33290 42340
rect 33210 42160 33220 42230
rect 33220 42160 33290 42230
rect 36718 63768 36782 65192
rect 38200 64500 38210 64570
rect 38210 64500 38280 64570
rect 38200 64390 38210 64460
rect 38210 64390 38280 64460
rect 41708 65478 41772 66902
rect 43190 66210 43200 66280
rect 43200 66210 43270 66280
rect 43190 66100 43200 66170
rect 43200 66100 43270 66170
rect 36718 62058 36782 63482
rect 36718 60348 36782 61772
rect 36718 58638 36782 60062
rect 36718 56928 36782 58352
rect 36718 55218 36782 56642
rect 36718 53508 36782 54932
rect 36718 51798 36782 53222
rect 36718 50088 36782 51512
rect 36718 48378 36782 49802
rect 36718 46668 36782 48092
rect 36718 44958 36782 46382
rect 36718 43248 36782 44672
rect 31728 39828 31792 41252
rect 33210 40560 33220 40630
rect 33220 40560 33290 40630
rect 33210 40450 33220 40520
rect 33220 40450 33290 40520
rect 36718 41538 36782 42962
rect 38200 62790 38210 62860
rect 38210 62790 38280 62860
rect 38200 62680 38210 62750
rect 38210 62680 38280 62750
rect 38200 61080 38210 61150
rect 38210 61080 38280 61150
rect 38200 60970 38210 61040
rect 38210 60970 38280 61040
rect 38200 59370 38210 59440
rect 38210 59370 38280 59440
rect 38200 59260 38210 59330
rect 38210 59260 38280 59330
rect 38200 57660 38210 57730
rect 38210 57660 38280 57730
rect 38200 57550 38210 57620
rect 38210 57550 38280 57620
rect 38200 55950 38210 56020
rect 38210 55950 38280 56020
rect 38200 55840 38210 55910
rect 38210 55840 38280 55910
rect 38200 54240 38210 54310
rect 38210 54240 38280 54310
rect 38200 54130 38210 54200
rect 38210 54130 38280 54200
rect 38200 52530 38210 52600
rect 38210 52530 38280 52600
rect 38200 52420 38210 52490
rect 38210 52420 38280 52490
rect 38200 50820 38210 50890
rect 38210 50820 38280 50890
rect 38200 50710 38210 50780
rect 38210 50710 38280 50780
rect 38200 49110 38210 49180
rect 38210 49110 38280 49180
rect 38200 49000 38210 49070
rect 38210 49000 38280 49070
rect 38200 47400 38210 47470
rect 38210 47400 38280 47470
rect 38200 47290 38210 47360
rect 38210 47290 38280 47360
rect 38200 45690 38210 45760
rect 38210 45690 38280 45760
rect 38200 45580 38210 45650
rect 38210 45580 38280 45650
rect 38200 43980 38210 44050
rect 38210 43980 38280 44050
rect 38200 43870 38210 43940
rect 38210 43870 38280 43940
rect 38200 42270 38210 42340
rect 38210 42270 38280 42340
rect 38200 42160 38210 42230
rect 38210 42160 38280 42230
rect 41708 63768 41772 65192
rect 43190 64500 43200 64570
rect 43200 64500 43270 64570
rect 43190 64390 43200 64460
rect 43200 64390 43270 64460
rect 46698 65478 46762 66902
rect 48180 66210 48190 66280
rect 48190 66210 48260 66280
rect 48180 66100 48190 66170
rect 48190 66100 48260 66170
rect 41708 62058 41772 63482
rect 41708 60348 41772 61772
rect 41708 58638 41772 60062
rect 41708 56928 41772 58352
rect 41708 55218 41772 56642
rect 41708 53508 41772 54932
rect 41708 51798 41772 53222
rect 41708 50088 41772 51512
rect 41708 48378 41772 49802
rect 41708 46668 41772 48092
rect 41708 44958 41772 46382
rect 41708 43248 41772 44672
rect 36718 39828 36782 41252
rect 38200 40560 38210 40630
rect 38210 40560 38280 40630
rect 38200 40450 38210 40520
rect 38210 40450 38280 40520
rect 41708 41538 41772 42962
rect 43190 62790 43200 62860
rect 43200 62790 43270 62860
rect 43190 62680 43200 62750
rect 43200 62680 43270 62750
rect 43190 61080 43200 61150
rect 43200 61080 43270 61150
rect 43190 60970 43200 61040
rect 43200 60970 43270 61040
rect 43190 59370 43200 59440
rect 43200 59370 43270 59440
rect 43190 59260 43200 59330
rect 43200 59260 43270 59330
rect 43190 57660 43200 57730
rect 43200 57660 43270 57730
rect 43190 57550 43200 57620
rect 43200 57550 43270 57620
rect 43190 55950 43200 56020
rect 43200 55950 43270 56020
rect 43190 55840 43200 55910
rect 43200 55840 43270 55910
rect 43190 54240 43200 54310
rect 43200 54240 43270 54310
rect 43190 54130 43200 54200
rect 43200 54130 43270 54200
rect 43190 52530 43200 52600
rect 43200 52530 43270 52600
rect 43190 52420 43200 52490
rect 43200 52420 43270 52490
rect 43190 50820 43200 50890
rect 43200 50820 43270 50890
rect 43190 50710 43200 50780
rect 43200 50710 43270 50780
rect 43190 49110 43200 49180
rect 43200 49110 43270 49180
rect 43190 49000 43200 49070
rect 43200 49000 43270 49070
rect 43190 47400 43200 47470
rect 43200 47400 43270 47470
rect 43190 47290 43200 47360
rect 43200 47290 43270 47360
rect 43190 45690 43200 45760
rect 43200 45690 43270 45760
rect 43190 45580 43200 45650
rect 43200 45580 43270 45650
rect 43190 43980 43200 44050
rect 43200 43980 43270 44050
rect 43190 43870 43200 43940
rect 43200 43870 43270 43940
rect 43190 42270 43200 42340
rect 43200 42270 43270 42340
rect 43190 42160 43200 42230
rect 43200 42160 43270 42230
rect 46698 63768 46762 65192
rect 48180 64500 48190 64570
rect 48190 64500 48260 64570
rect 48180 64390 48190 64460
rect 48190 64390 48260 64460
rect 51688 65478 51752 66902
rect 53170 66210 53180 66280
rect 53180 66210 53250 66280
rect 53170 66100 53180 66170
rect 53180 66100 53250 66170
rect 46698 62058 46762 63482
rect 46698 60348 46762 61772
rect 46698 58638 46762 60062
rect 46698 56928 46762 58352
rect 46698 55218 46762 56642
rect 46698 53508 46762 54932
rect 46698 51798 46762 53222
rect 46698 50088 46762 51512
rect 46698 48378 46762 49802
rect 46698 46668 46762 48092
rect 46698 44958 46762 46382
rect 46698 43248 46762 44672
rect 41708 39828 41772 41252
rect 43190 40560 43200 40630
rect 43200 40560 43270 40630
rect 43190 40450 43200 40520
rect 43200 40450 43270 40520
rect 46698 41538 46762 42962
rect 48180 62790 48190 62860
rect 48190 62790 48260 62860
rect 48180 62680 48190 62750
rect 48190 62680 48260 62750
rect 48180 61080 48190 61150
rect 48190 61080 48260 61150
rect 48180 60970 48190 61040
rect 48190 60970 48260 61040
rect 48180 59370 48190 59440
rect 48190 59370 48260 59440
rect 48180 59260 48190 59330
rect 48190 59260 48260 59330
rect 48180 57660 48190 57730
rect 48190 57660 48260 57730
rect 48180 57550 48190 57620
rect 48190 57550 48260 57620
rect 48180 55950 48190 56020
rect 48190 55950 48260 56020
rect 48180 55840 48190 55910
rect 48190 55840 48260 55910
rect 48180 54240 48190 54310
rect 48190 54240 48260 54310
rect 48180 54130 48190 54200
rect 48190 54130 48260 54200
rect 48180 52530 48190 52600
rect 48190 52530 48260 52600
rect 48180 52420 48190 52490
rect 48190 52420 48260 52490
rect 48180 50820 48190 50890
rect 48190 50820 48260 50890
rect 48180 50710 48190 50780
rect 48190 50710 48260 50780
rect 48180 49110 48190 49180
rect 48190 49110 48260 49180
rect 48180 49000 48190 49070
rect 48190 49000 48260 49070
rect 48180 47400 48190 47470
rect 48190 47400 48260 47470
rect 48180 47290 48190 47360
rect 48190 47290 48260 47360
rect 48180 45690 48190 45760
rect 48190 45690 48260 45760
rect 48180 45580 48190 45650
rect 48190 45580 48260 45650
rect 48180 43980 48190 44050
rect 48190 43980 48260 44050
rect 48180 43870 48190 43940
rect 48190 43870 48260 43940
rect 48180 42270 48190 42340
rect 48190 42270 48260 42340
rect 48180 42160 48190 42230
rect 48190 42160 48260 42230
rect 51688 63768 51752 65192
rect 53170 64500 53180 64570
rect 53180 64500 53250 64570
rect 53170 64390 53180 64460
rect 53180 64390 53250 64460
rect 56678 65478 56742 66902
rect 58160 66210 58170 66280
rect 58170 66210 58240 66280
rect 58160 66100 58170 66170
rect 58170 66100 58240 66170
rect 51688 62058 51752 63482
rect 51688 60348 51752 61772
rect 51688 58638 51752 60062
rect 51688 56928 51752 58352
rect 51688 55218 51752 56642
rect 51688 53508 51752 54932
rect 51688 51798 51752 53222
rect 51688 50088 51752 51512
rect 51688 48378 51752 49802
rect 51688 46668 51752 48092
rect 51688 44958 51752 46382
rect 51688 43248 51752 44672
rect 46698 39828 46762 41252
rect 48180 40560 48190 40630
rect 48190 40560 48260 40630
rect 48180 40450 48190 40520
rect 48190 40450 48260 40520
rect 51688 41538 51752 42962
rect 53170 62790 53180 62860
rect 53180 62790 53250 62860
rect 53170 62680 53180 62750
rect 53180 62680 53250 62750
rect 53170 61080 53180 61150
rect 53180 61080 53250 61150
rect 53170 60970 53180 61040
rect 53180 60970 53250 61040
rect 53170 59370 53180 59440
rect 53180 59370 53250 59440
rect 53170 59260 53180 59330
rect 53180 59260 53250 59330
rect 53170 57660 53180 57730
rect 53180 57660 53250 57730
rect 53170 57550 53180 57620
rect 53180 57550 53250 57620
rect 53170 55950 53180 56020
rect 53180 55950 53250 56020
rect 53170 55840 53180 55910
rect 53180 55840 53250 55910
rect 53170 54240 53180 54310
rect 53180 54240 53250 54310
rect 53170 54130 53180 54200
rect 53180 54130 53250 54200
rect 53170 52530 53180 52600
rect 53180 52530 53250 52600
rect 53170 52420 53180 52490
rect 53180 52420 53250 52490
rect 53170 50820 53180 50890
rect 53180 50820 53250 50890
rect 53170 50710 53180 50780
rect 53180 50710 53250 50780
rect 53170 49110 53180 49180
rect 53180 49110 53250 49180
rect 53170 49000 53180 49070
rect 53180 49000 53250 49070
rect 53170 47400 53180 47470
rect 53180 47400 53250 47470
rect 53170 47290 53180 47360
rect 53180 47290 53250 47360
rect 53170 45690 53180 45760
rect 53180 45690 53250 45760
rect 53170 45580 53180 45650
rect 53180 45580 53250 45650
rect 53170 43980 53180 44050
rect 53180 43980 53250 44050
rect 53170 43870 53180 43940
rect 53180 43870 53250 43940
rect 53170 42270 53180 42340
rect 53180 42270 53250 42340
rect 53170 42160 53180 42230
rect 53180 42160 53250 42230
rect 56678 63768 56742 65192
rect 58160 64500 58170 64570
rect 58170 64500 58240 64570
rect 58160 64390 58170 64460
rect 58170 64390 58240 64460
rect 61668 65478 61732 66902
rect 63150 66210 63160 66280
rect 63160 66210 63230 66280
rect 63150 66100 63160 66170
rect 63160 66100 63230 66170
rect 56678 62058 56742 63482
rect 56678 60348 56742 61772
rect 56678 58638 56742 60062
rect 56678 56928 56742 58352
rect 56678 55218 56742 56642
rect 56678 53508 56742 54932
rect 56678 51798 56742 53222
rect 56678 50088 56742 51512
rect 56678 48378 56742 49802
rect 56678 46668 56742 48092
rect 56678 44958 56742 46382
rect 56678 43248 56742 44672
rect 51688 39828 51752 41252
rect 53170 40560 53180 40630
rect 53180 40560 53250 40630
rect 53170 40450 53180 40520
rect 53180 40450 53250 40520
rect 56678 41538 56742 42962
rect 58160 62790 58170 62860
rect 58170 62790 58240 62860
rect 58160 62680 58170 62750
rect 58170 62680 58240 62750
rect 58160 61080 58170 61150
rect 58170 61080 58240 61150
rect 58160 60970 58170 61040
rect 58170 60970 58240 61040
rect 58160 59370 58170 59440
rect 58170 59370 58240 59440
rect 58160 59260 58170 59330
rect 58170 59260 58240 59330
rect 58160 57660 58170 57730
rect 58170 57660 58240 57730
rect 58160 57550 58170 57620
rect 58170 57550 58240 57620
rect 58160 55950 58170 56020
rect 58170 55950 58240 56020
rect 58160 55840 58170 55910
rect 58170 55840 58240 55910
rect 58160 54240 58170 54310
rect 58170 54240 58240 54310
rect 58160 54130 58170 54200
rect 58170 54130 58240 54200
rect 58160 52530 58170 52600
rect 58170 52530 58240 52600
rect 58160 52420 58170 52490
rect 58170 52420 58240 52490
rect 58160 50820 58170 50890
rect 58170 50820 58240 50890
rect 58160 50710 58170 50780
rect 58170 50710 58240 50780
rect 58160 49110 58170 49180
rect 58170 49110 58240 49180
rect 58160 49000 58170 49070
rect 58170 49000 58240 49070
rect 58160 47400 58170 47470
rect 58170 47400 58240 47470
rect 58160 47290 58170 47360
rect 58170 47290 58240 47360
rect 58160 45690 58170 45760
rect 58170 45690 58240 45760
rect 58160 45580 58170 45650
rect 58170 45580 58240 45650
rect 58160 43980 58170 44050
rect 58170 43980 58240 44050
rect 58160 43870 58170 43940
rect 58170 43870 58240 43940
rect 58160 42270 58170 42340
rect 58170 42270 58240 42340
rect 58160 42160 58170 42230
rect 58170 42160 58240 42230
rect 61668 63768 61732 65192
rect 63150 64500 63160 64570
rect 63160 64500 63230 64570
rect 63150 64390 63160 64460
rect 63160 64390 63230 64460
rect 66658 65478 66722 66902
rect 68140 66210 68150 66280
rect 68150 66210 68220 66280
rect 68140 66100 68150 66170
rect 68150 66100 68220 66170
rect 61668 62058 61732 63482
rect 63150 62790 63160 62860
rect 63160 62790 63230 62860
rect 63150 62680 63160 62750
rect 63160 62680 63230 62750
rect 66658 63768 66722 65192
rect 68140 64500 68150 64570
rect 68150 64500 68220 64570
rect 68140 64390 68150 64460
rect 68150 64390 68220 64460
rect 71648 65478 71712 66902
rect 73130 66210 73140 66280
rect 73140 66210 73210 66280
rect 73130 66100 73140 66170
rect 73140 66100 73210 66170
rect 61668 60348 61732 61772
rect 63150 61080 63160 61150
rect 63160 61080 63230 61150
rect 63150 60970 63160 61040
rect 63160 60970 63230 61040
rect 66658 62058 66722 63482
rect 68140 62790 68150 62860
rect 68150 62790 68220 62860
rect 68140 62680 68150 62750
rect 68150 62680 68220 62750
rect 71648 63768 71712 65192
rect 73130 64500 73140 64570
rect 73140 64500 73210 64570
rect 73130 64390 73140 64460
rect 73140 64390 73210 64460
rect 76638 65478 76702 66902
rect 78120 66210 78130 66280
rect 78130 66210 78200 66280
rect 78120 66100 78130 66170
rect 78130 66100 78200 66170
rect 61668 58638 61732 60062
rect 61668 56928 61732 58352
rect 61668 55218 61732 56642
rect 61668 53508 61732 54932
rect 61668 51798 61732 53222
rect 61668 50088 61732 51512
rect 61668 48378 61732 49802
rect 61668 46668 61732 48092
rect 61668 44958 61732 46382
rect 63150 59370 63160 59440
rect 63160 59370 63230 59440
rect 63150 59260 63160 59330
rect 63160 59260 63230 59330
rect 63150 57660 63160 57730
rect 63160 57660 63230 57730
rect 63150 57550 63160 57620
rect 63160 57550 63230 57620
rect 63150 55950 63160 56020
rect 63160 55950 63230 56020
rect 63150 55840 63160 55910
rect 63160 55840 63230 55910
rect 63150 54240 63160 54310
rect 63160 54240 63230 54310
rect 63150 54130 63160 54200
rect 63160 54130 63230 54200
rect 63150 52530 63160 52600
rect 63160 52530 63230 52600
rect 63150 52420 63160 52490
rect 63160 52420 63230 52490
rect 63150 50820 63160 50890
rect 63160 50820 63230 50890
rect 63150 50710 63160 50780
rect 63160 50710 63230 50780
rect 63150 49110 63160 49180
rect 63160 49110 63230 49180
rect 63150 49000 63160 49070
rect 63160 49000 63230 49070
rect 63150 47400 63160 47470
rect 63160 47400 63230 47470
rect 63150 47290 63160 47360
rect 63160 47290 63230 47360
rect 63150 45690 63160 45760
rect 63160 45690 63230 45760
rect 63150 45580 63160 45650
rect 63160 45580 63230 45650
rect 66658 60348 66722 61772
rect 68140 61080 68150 61150
rect 68150 61080 68220 61150
rect 68140 60970 68150 61040
rect 68150 60970 68220 61040
rect 71648 62058 71712 63482
rect 73130 62790 73140 62860
rect 73140 62790 73210 62860
rect 73130 62680 73140 62750
rect 73140 62680 73210 62750
rect 76638 63768 76702 65192
rect 78120 64500 78130 64570
rect 78130 64500 78200 64570
rect 78120 64390 78130 64460
rect 78130 64390 78200 64460
rect 66658 58638 66722 60062
rect 66658 56928 66722 58352
rect 66658 55218 66722 56642
rect 66658 53508 66722 54932
rect 66658 51798 66722 53222
rect 66658 50088 66722 51512
rect 66658 48378 66722 49802
rect 66658 46668 66722 48092
rect 61668 43248 61732 44672
rect 63150 43980 63160 44050
rect 63160 43980 63230 44050
rect 63150 43870 63160 43940
rect 63160 43870 63230 43940
rect 66658 44958 66722 46382
rect 68140 59370 68150 59440
rect 68150 59370 68220 59440
rect 68140 59260 68150 59330
rect 68150 59260 68220 59330
rect 68140 57660 68150 57730
rect 68150 57660 68220 57730
rect 68140 57550 68150 57620
rect 68150 57550 68220 57620
rect 68140 55950 68150 56020
rect 68150 55950 68220 56020
rect 68140 55840 68150 55910
rect 68150 55840 68220 55910
rect 68140 54240 68150 54310
rect 68150 54240 68220 54310
rect 68140 54130 68150 54200
rect 68150 54130 68220 54200
rect 68140 52530 68150 52600
rect 68150 52530 68220 52600
rect 68140 52420 68150 52490
rect 68150 52420 68220 52490
rect 68140 50820 68150 50890
rect 68150 50820 68220 50890
rect 68140 50710 68150 50780
rect 68150 50710 68220 50780
rect 68140 49110 68150 49180
rect 68150 49110 68220 49180
rect 68140 49000 68150 49070
rect 68150 49000 68220 49070
rect 68140 47400 68150 47470
rect 68150 47400 68220 47470
rect 68140 47290 68150 47360
rect 68150 47290 68220 47360
rect 68140 45690 68150 45760
rect 68150 45690 68220 45760
rect 68140 45580 68150 45650
rect 68150 45580 68220 45650
rect 71648 60348 71712 61772
rect 73130 61080 73140 61150
rect 73140 61080 73210 61150
rect 73130 60970 73140 61040
rect 73140 60970 73210 61040
rect 76638 62058 76702 63482
rect 78120 62790 78130 62860
rect 78130 62790 78200 62860
rect 78120 62680 78130 62750
rect 78130 62680 78200 62750
rect 71648 58638 71712 60062
rect 73130 59370 73140 59440
rect 73140 59370 73210 59440
rect 73130 59260 73140 59330
rect 73140 59260 73210 59330
rect 76638 60348 76702 61772
rect 78120 61080 78130 61150
rect 78130 61080 78200 61150
rect 78120 60970 78130 61040
rect 78130 60970 78200 61040
rect 71648 56928 71712 58352
rect 73130 57660 73140 57730
rect 73140 57660 73210 57730
rect 73130 57550 73140 57620
rect 73140 57550 73210 57620
rect 76638 58638 76702 60062
rect 78120 59370 78130 59440
rect 78130 59370 78200 59440
rect 78120 59260 78130 59330
rect 78130 59260 78200 59330
rect 71648 55218 71712 56642
rect 73130 55950 73140 56020
rect 73140 55950 73210 56020
rect 73130 55840 73140 55910
rect 73140 55840 73210 55910
rect 76638 56928 76702 58352
rect 78120 57660 78130 57730
rect 78130 57660 78200 57730
rect 78120 57550 78130 57620
rect 78130 57550 78200 57620
rect 71648 53508 71712 54932
rect 73130 54240 73140 54310
rect 73140 54240 73210 54310
rect 73130 54130 73140 54200
rect 73140 54130 73210 54200
rect 76638 55218 76702 56642
rect 78120 55950 78130 56020
rect 78130 55950 78200 56020
rect 78120 55840 78130 55910
rect 78130 55840 78200 55910
rect 71648 51798 71712 53222
rect 73130 52530 73140 52600
rect 73140 52530 73210 52600
rect 73130 52420 73140 52490
rect 73140 52420 73210 52490
rect 76638 53508 76702 54932
rect 78120 54240 78130 54310
rect 78130 54240 78200 54310
rect 78120 54130 78130 54200
rect 78130 54130 78200 54200
rect 71648 50088 71712 51512
rect 73130 50820 73140 50890
rect 73140 50820 73210 50890
rect 73130 50710 73140 50780
rect 73140 50710 73210 50780
rect 76638 51798 76702 53222
rect 78120 52530 78130 52600
rect 78130 52530 78200 52600
rect 78120 52420 78130 52490
rect 78130 52420 78200 52490
rect 71648 48378 71712 49802
rect 73130 49110 73140 49180
rect 73140 49110 73210 49180
rect 73130 49000 73140 49070
rect 73140 49000 73210 49070
rect 76638 50088 76702 51512
rect 78120 50820 78130 50890
rect 78130 50820 78200 50890
rect 78120 50710 78130 50780
rect 78130 50710 78200 50780
rect 71648 46668 71712 48092
rect 73130 47400 73140 47470
rect 73140 47400 73210 47470
rect 73130 47290 73140 47360
rect 73140 47290 73210 47360
rect 76638 48378 76702 49802
rect 78120 49110 78130 49180
rect 78130 49110 78200 49180
rect 78120 49000 78130 49070
rect 78130 49000 78200 49070
rect 56678 39828 56742 41252
rect 58160 40560 58170 40630
rect 58170 40560 58240 40630
rect 58160 40450 58170 40520
rect 58170 40450 58240 40520
rect 61668 41538 61732 42962
rect 63150 42270 63160 42340
rect 63160 42270 63230 42340
rect 63150 42160 63160 42230
rect 63160 42160 63230 42230
rect 66658 43248 66722 44672
rect 68140 43980 68150 44050
rect 68150 43980 68220 44050
rect 68140 43870 68150 43940
rect 68150 43870 68220 43940
rect 71648 44958 71712 46382
rect 73130 45690 73140 45760
rect 73140 45690 73210 45760
rect 73130 45580 73140 45650
rect 73140 45580 73210 45650
rect 76638 46668 76702 48092
rect 78120 47400 78130 47470
rect 78130 47400 78200 47470
rect 78120 47290 78130 47360
rect 78130 47290 78200 47360
rect 61668 39828 61732 41252
rect 63150 40560 63160 40630
rect 63160 40560 63230 40630
rect 63150 40450 63160 40520
rect 63160 40450 63230 40520
rect 66658 41538 66722 42962
rect 68140 42270 68150 42340
rect 68150 42270 68220 42340
rect 68140 42160 68150 42230
rect 68150 42160 68220 42230
rect 71648 43248 71712 44672
rect 73130 43980 73140 44050
rect 73140 43980 73210 44050
rect 73130 43870 73140 43940
rect 73140 43870 73210 43940
rect 76638 44958 76702 46382
rect 78120 45690 78130 45760
rect 78130 45690 78200 45760
rect 78120 45580 78130 45650
rect 78130 45580 78200 45650
rect 66658 39828 66722 41252
rect 68140 40560 68150 40630
rect 68150 40560 68220 40630
rect 68140 40450 68150 40520
rect 68150 40450 68220 40520
rect 71648 41538 71712 42962
rect 73130 42270 73140 42340
rect 73140 42270 73210 42340
rect 73130 42160 73140 42230
rect 73140 42160 73210 42230
rect 76638 43248 76702 44672
rect 78120 43980 78130 44050
rect 78130 43980 78200 44050
rect 78120 43870 78130 43940
rect 78130 43870 78200 43940
rect 71648 39828 71712 41252
rect 73130 40560 73140 40630
rect 73140 40560 73210 40630
rect 73130 40450 73140 40520
rect 73140 40450 73210 40520
rect 76638 41538 76702 42962
rect 78120 42270 78130 42340
rect 78130 42270 78200 42340
rect 78120 42160 78130 42230
rect 78130 42160 78200 42230
rect 76638 39828 76702 41252
rect 78120 40560 78130 40630
rect 78130 40560 78200 40630
rect 78120 40450 78130 40520
rect 78130 40450 78200 40520
<< mimcap >>
rect 140 66850 1540 66890
rect 140 65530 180 66850
rect 1500 65530 1540 66850
rect 140 65490 1540 65530
rect 5130 66850 6530 66890
rect 5130 65530 5170 66850
rect 6490 65530 6530 66850
rect 5130 65490 6530 65530
rect 10120 66850 11520 66890
rect 10120 65530 10160 66850
rect 11480 65530 11520 66850
rect 10120 65490 11520 65530
rect 15110 66850 16510 66890
rect 15110 65530 15150 66850
rect 16470 65530 16510 66850
rect 15110 65490 16510 65530
rect 20100 66850 21500 66890
rect 20100 65530 20140 66850
rect 21460 65530 21500 66850
rect 20100 65490 21500 65530
rect 25090 66850 26490 66890
rect 25090 65530 25130 66850
rect 26450 65530 26490 66850
rect 25090 65490 26490 65530
rect 30080 66850 31480 66890
rect 30080 65530 30120 66850
rect 31440 65530 31480 66850
rect 30080 65490 31480 65530
rect 35070 66850 36470 66890
rect 35070 65530 35110 66850
rect 36430 65530 36470 66850
rect 35070 65490 36470 65530
rect 40060 66850 41460 66890
rect 40060 65530 40100 66850
rect 41420 65530 41460 66850
rect 40060 65490 41460 65530
rect 45050 66850 46450 66890
rect 45050 65530 45090 66850
rect 46410 65530 46450 66850
rect 45050 65490 46450 65530
rect 50040 66850 51440 66890
rect 50040 65530 50080 66850
rect 51400 65530 51440 66850
rect 50040 65490 51440 65530
rect 55030 66850 56430 66890
rect 55030 65530 55070 66850
rect 56390 65530 56430 66850
rect 55030 65490 56430 65530
rect 60020 66850 61420 66890
rect 60020 65530 60060 66850
rect 61380 65530 61420 66850
rect 60020 65490 61420 65530
rect 65010 66850 66410 66890
rect 65010 65530 65050 66850
rect 66370 65530 66410 66850
rect 65010 65490 66410 65530
rect 70000 66850 71400 66890
rect 70000 65530 70040 66850
rect 71360 65530 71400 66850
rect 70000 65490 71400 65530
rect 74990 66850 76390 66890
rect 74990 65530 75030 66850
rect 76350 65530 76390 66850
rect 74990 65490 76390 65530
rect 140 65140 1540 65180
rect 140 63820 180 65140
rect 1500 63820 1540 65140
rect 140 63780 1540 63820
rect 5130 65140 6530 65180
rect 5130 63820 5170 65140
rect 6490 63820 6530 65140
rect 5130 63780 6530 63820
rect 10120 65140 11520 65180
rect 10120 63820 10160 65140
rect 11480 63820 11520 65140
rect 10120 63780 11520 63820
rect 15110 65140 16510 65180
rect 15110 63820 15150 65140
rect 16470 63820 16510 65140
rect 15110 63780 16510 63820
rect 20100 65140 21500 65180
rect 20100 63820 20140 65140
rect 21460 63820 21500 65140
rect 20100 63780 21500 63820
rect 25090 65140 26490 65180
rect 25090 63820 25130 65140
rect 26450 63820 26490 65140
rect 25090 63780 26490 63820
rect 30080 65140 31480 65180
rect 30080 63820 30120 65140
rect 31440 63820 31480 65140
rect 30080 63780 31480 63820
rect 35070 65140 36470 65180
rect 35070 63820 35110 65140
rect 36430 63820 36470 65140
rect 35070 63780 36470 63820
rect 40060 65140 41460 65180
rect 40060 63820 40100 65140
rect 41420 63820 41460 65140
rect 40060 63780 41460 63820
rect 45050 65140 46450 65180
rect 45050 63820 45090 65140
rect 46410 63820 46450 65140
rect 45050 63780 46450 63820
rect 50040 65140 51440 65180
rect 50040 63820 50080 65140
rect 51400 63820 51440 65140
rect 50040 63780 51440 63820
rect 55030 65140 56430 65180
rect 55030 63820 55070 65140
rect 56390 63820 56430 65140
rect 55030 63780 56430 63820
rect 60020 65140 61420 65180
rect 60020 63820 60060 65140
rect 61380 63820 61420 65140
rect 60020 63780 61420 63820
rect 65010 65140 66410 65180
rect 65010 63820 65050 65140
rect 66370 63820 66410 65140
rect 65010 63780 66410 63820
rect 70000 65140 71400 65180
rect 70000 63820 70040 65140
rect 71360 63820 71400 65140
rect 70000 63780 71400 63820
rect 74990 65140 76390 65180
rect 74990 63820 75030 65140
rect 76350 63820 76390 65140
rect 74990 63780 76390 63820
rect 140 63430 1540 63470
rect 140 62110 180 63430
rect 1500 62110 1540 63430
rect 140 62070 1540 62110
rect 5130 63430 6530 63470
rect 5130 62110 5170 63430
rect 6490 62110 6530 63430
rect 5130 62070 6530 62110
rect 10120 63430 11520 63470
rect 10120 62110 10160 63430
rect 11480 62110 11520 63430
rect 10120 62070 11520 62110
rect 15110 63430 16510 63470
rect 15110 62110 15150 63430
rect 16470 62110 16510 63430
rect 15110 62070 16510 62110
rect 20100 63430 21500 63470
rect 20100 62110 20140 63430
rect 21460 62110 21500 63430
rect 20100 62070 21500 62110
rect 25090 63430 26490 63470
rect 25090 62110 25130 63430
rect 26450 62110 26490 63430
rect 25090 62070 26490 62110
rect 30080 63430 31480 63470
rect 30080 62110 30120 63430
rect 31440 62110 31480 63430
rect 30080 62070 31480 62110
rect 35070 63430 36470 63470
rect 35070 62110 35110 63430
rect 36430 62110 36470 63430
rect 35070 62070 36470 62110
rect 40060 63430 41460 63470
rect 40060 62110 40100 63430
rect 41420 62110 41460 63430
rect 40060 62070 41460 62110
rect 45050 63430 46450 63470
rect 45050 62110 45090 63430
rect 46410 62110 46450 63430
rect 45050 62070 46450 62110
rect 50040 63430 51440 63470
rect 50040 62110 50080 63430
rect 51400 62110 51440 63430
rect 50040 62070 51440 62110
rect 55030 63430 56430 63470
rect 55030 62110 55070 63430
rect 56390 62110 56430 63430
rect 55030 62070 56430 62110
rect 60020 63430 61420 63470
rect 60020 62110 60060 63430
rect 61380 62110 61420 63430
rect 60020 62070 61420 62110
rect 65010 63430 66410 63470
rect 65010 62110 65050 63430
rect 66370 62110 66410 63430
rect 65010 62070 66410 62110
rect 70000 63430 71400 63470
rect 70000 62110 70040 63430
rect 71360 62110 71400 63430
rect 70000 62070 71400 62110
rect 74990 63430 76390 63470
rect 74990 62110 75030 63430
rect 76350 62110 76390 63430
rect 74990 62070 76390 62110
rect 140 61720 1540 61760
rect 140 60400 180 61720
rect 1500 60400 1540 61720
rect 140 60360 1540 60400
rect 5130 61720 6530 61760
rect 5130 60400 5170 61720
rect 6490 60400 6530 61720
rect 5130 60360 6530 60400
rect 10120 61720 11520 61760
rect 10120 60400 10160 61720
rect 11480 60400 11520 61720
rect 10120 60360 11520 60400
rect 15110 61720 16510 61760
rect 15110 60400 15150 61720
rect 16470 60400 16510 61720
rect 15110 60360 16510 60400
rect 20100 61720 21500 61760
rect 20100 60400 20140 61720
rect 21460 60400 21500 61720
rect 20100 60360 21500 60400
rect 25090 61720 26490 61760
rect 25090 60400 25130 61720
rect 26450 60400 26490 61720
rect 25090 60360 26490 60400
rect 30080 61720 31480 61760
rect 30080 60400 30120 61720
rect 31440 60400 31480 61720
rect 30080 60360 31480 60400
rect 35070 61720 36470 61760
rect 35070 60400 35110 61720
rect 36430 60400 36470 61720
rect 35070 60360 36470 60400
rect 40060 61720 41460 61760
rect 40060 60400 40100 61720
rect 41420 60400 41460 61720
rect 40060 60360 41460 60400
rect 45050 61720 46450 61760
rect 45050 60400 45090 61720
rect 46410 60400 46450 61720
rect 45050 60360 46450 60400
rect 50040 61720 51440 61760
rect 50040 60400 50080 61720
rect 51400 60400 51440 61720
rect 50040 60360 51440 60400
rect 55030 61720 56430 61760
rect 55030 60400 55070 61720
rect 56390 60400 56430 61720
rect 55030 60360 56430 60400
rect 60020 61720 61420 61760
rect 60020 60400 60060 61720
rect 61380 60400 61420 61720
rect 60020 60360 61420 60400
rect 65010 61720 66410 61760
rect 65010 60400 65050 61720
rect 66370 60400 66410 61720
rect 65010 60360 66410 60400
rect 70000 61720 71400 61760
rect 70000 60400 70040 61720
rect 71360 60400 71400 61720
rect 70000 60360 71400 60400
rect 74990 61720 76390 61760
rect 74990 60400 75030 61720
rect 76350 60400 76390 61720
rect 74990 60360 76390 60400
rect 140 60010 1540 60050
rect 140 58690 180 60010
rect 1500 58690 1540 60010
rect 140 58650 1540 58690
rect 5130 60010 6530 60050
rect 5130 58690 5170 60010
rect 6490 58690 6530 60010
rect 5130 58650 6530 58690
rect 10120 60010 11520 60050
rect 10120 58690 10160 60010
rect 11480 58690 11520 60010
rect 10120 58650 11520 58690
rect 15110 60010 16510 60050
rect 15110 58690 15150 60010
rect 16470 58690 16510 60010
rect 15110 58650 16510 58690
rect 20100 60010 21500 60050
rect 20100 58690 20140 60010
rect 21460 58690 21500 60010
rect 20100 58650 21500 58690
rect 25090 60010 26490 60050
rect 25090 58690 25130 60010
rect 26450 58690 26490 60010
rect 25090 58650 26490 58690
rect 30080 60010 31480 60050
rect 30080 58690 30120 60010
rect 31440 58690 31480 60010
rect 30080 58650 31480 58690
rect 35070 60010 36470 60050
rect 35070 58690 35110 60010
rect 36430 58690 36470 60010
rect 35070 58650 36470 58690
rect 40060 60010 41460 60050
rect 40060 58690 40100 60010
rect 41420 58690 41460 60010
rect 40060 58650 41460 58690
rect 45050 60010 46450 60050
rect 45050 58690 45090 60010
rect 46410 58690 46450 60010
rect 45050 58650 46450 58690
rect 50040 60010 51440 60050
rect 50040 58690 50080 60010
rect 51400 58690 51440 60010
rect 50040 58650 51440 58690
rect 55030 60010 56430 60050
rect 55030 58690 55070 60010
rect 56390 58690 56430 60010
rect 55030 58650 56430 58690
rect 60020 60010 61420 60050
rect 60020 58690 60060 60010
rect 61380 58690 61420 60010
rect 60020 58650 61420 58690
rect 65010 60010 66410 60050
rect 65010 58690 65050 60010
rect 66370 58690 66410 60010
rect 65010 58650 66410 58690
rect 70000 60010 71400 60050
rect 70000 58690 70040 60010
rect 71360 58690 71400 60010
rect 70000 58650 71400 58690
rect 74990 60010 76390 60050
rect 74990 58690 75030 60010
rect 76350 58690 76390 60010
rect 74990 58650 76390 58690
rect 140 58300 1540 58340
rect 140 56980 180 58300
rect 1500 56980 1540 58300
rect 140 56940 1540 56980
rect 5130 58300 6530 58340
rect 5130 56980 5170 58300
rect 6490 56980 6530 58300
rect 5130 56940 6530 56980
rect 10120 58300 11520 58340
rect 10120 56980 10160 58300
rect 11480 56980 11520 58300
rect 10120 56940 11520 56980
rect 15110 58300 16510 58340
rect 15110 56980 15150 58300
rect 16470 56980 16510 58300
rect 15110 56940 16510 56980
rect 20100 58300 21500 58340
rect 20100 56980 20140 58300
rect 21460 56980 21500 58300
rect 20100 56940 21500 56980
rect 25090 58300 26490 58340
rect 25090 56980 25130 58300
rect 26450 56980 26490 58300
rect 25090 56940 26490 56980
rect 30080 58300 31480 58340
rect 30080 56980 30120 58300
rect 31440 56980 31480 58300
rect 30080 56940 31480 56980
rect 35070 58300 36470 58340
rect 35070 56980 35110 58300
rect 36430 56980 36470 58300
rect 35070 56940 36470 56980
rect 40060 58300 41460 58340
rect 40060 56980 40100 58300
rect 41420 56980 41460 58300
rect 40060 56940 41460 56980
rect 45050 58300 46450 58340
rect 45050 56980 45090 58300
rect 46410 56980 46450 58300
rect 45050 56940 46450 56980
rect 50040 58300 51440 58340
rect 50040 56980 50080 58300
rect 51400 56980 51440 58300
rect 50040 56940 51440 56980
rect 55030 58300 56430 58340
rect 55030 56980 55070 58300
rect 56390 56980 56430 58300
rect 55030 56940 56430 56980
rect 60020 58300 61420 58340
rect 60020 56980 60060 58300
rect 61380 56980 61420 58300
rect 60020 56940 61420 56980
rect 65010 58300 66410 58340
rect 65010 56980 65050 58300
rect 66370 56980 66410 58300
rect 65010 56940 66410 56980
rect 70000 58300 71400 58340
rect 70000 56980 70040 58300
rect 71360 56980 71400 58300
rect 70000 56940 71400 56980
rect 74990 58300 76390 58340
rect 74990 56980 75030 58300
rect 76350 56980 76390 58300
rect 74990 56940 76390 56980
rect 140 56590 1540 56630
rect 140 55270 180 56590
rect 1500 55270 1540 56590
rect 140 55230 1540 55270
rect 5130 56590 6530 56630
rect 5130 55270 5170 56590
rect 6490 55270 6530 56590
rect 5130 55230 6530 55270
rect 10120 56590 11520 56630
rect 10120 55270 10160 56590
rect 11480 55270 11520 56590
rect 10120 55230 11520 55270
rect 15110 56590 16510 56630
rect 15110 55270 15150 56590
rect 16470 55270 16510 56590
rect 15110 55230 16510 55270
rect 20100 56590 21500 56630
rect 20100 55270 20140 56590
rect 21460 55270 21500 56590
rect 20100 55230 21500 55270
rect 25090 56590 26490 56630
rect 25090 55270 25130 56590
rect 26450 55270 26490 56590
rect 25090 55230 26490 55270
rect 30080 56590 31480 56630
rect 30080 55270 30120 56590
rect 31440 55270 31480 56590
rect 30080 55230 31480 55270
rect 35070 56590 36470 56630
rect 35070 55270 35110 56590
rect 36430 55270 36470 56590
rect 35070 55230 36470 55270
rect 40060 56590 41460 56630
rect 40060 55270 40100 56590
rect 41420 55270 41460 56590
rect 40060 55230 41460 55270
rect 45050 56590 46450 56630
rect 45050 55270 45090 56590
rect 46410 55270 46450 56590
rect 45050 55230 46450 55270
rect 50040 56590 51440 56630
rect 50040 55270 50080 56590
rect 51400 55270 51440 56590
rect 50040 55230 51440 55270
rect 55030 56590 56430 56630
rect 55030 55270 55070 56590
rect 56390 55270 56430 56590
rect 55030 55230 56430 55270
rect 60020 56590 61420 56630
rect 60020 55270 60060 56590
rect 61380 55270 61420 56590
rect 60020 55230 61420 55270
rect 65010 56590 66410 56630
rect 65010 55270 65050 56590
rect 66370 55270 66410 56590
rect 65010 55230 66410 55270
rect 70000 56590 71400 56630
rect 70000 55270 70040 56590
rect 71360 55270 71400 56590
rect 70000 55230 71400 55270
rect 74990 56590 76390 56630
rect 74990 55270 75030 56590
rect 76350 55270 76390 56590
rect 74990 55230 76390 55270
rect 140 54880 1540 54920
rect 140 53560 180 54880
rect 1500 53560 1540 54880
rect 140 53520 1540 53560
rect 5130 54880 6530 54920
rect 5130 53560 5170 54880
rect 6490 53560 6530 54880
rect 5130 53520 6530 53560
rect 10120 54880 11520 54920
rect 10120 53560 10160 54880
rect 11480 53560 11520 54880
rect 10120 53520 11520 53560
rect 15110 54880 16510 54920
rect 15110 53560 15150 54880
rect 16470 53560 16510 54880
rect 15110 53520 16510 53560
rect 20100 54880 21500 54920
rect 20100 53560 20140 54880
rect 21460 53560 21500 54880
rect 20100 53520 21500 53560
rect 25090 54880 26490 54920
rect 25090 53560 25130 54880
rect 26450 53560 26490 54880
rect 25090 53520 26490 53560
rect 30080 54880 31480 54920
rect 30080 53560 30120 54880
rect 31440 53560 31480 54880
rect 30080 53520 31480 53560
rect 35070 54880 36470 54920
rect 35070 53560 35110 54880
rect 36430 53560 36470 54880
rect 35070 53520 36470 53560
rect 40060 54880 41460 54920
rect 40060 53560 40100 54880
rect 41420 53560 41460 54880
rect 40060 53520 41460 53560
rect 45050 54880 46450 54920
rect 45050 53560 45090 54880
rect 46410 53560 46450 54880
rect 45050 53520 46450 53560
rect 50040 54880 51440 54920
rect 50040 53560 50080 54880
rect 51400 53560 51440 54880
rect 50040 53520 51440 53560
rect 55030 54880 56430 54920
rect 55030 53560 55070 54880
rect 56390 53560 56430 54880
rect 55030 53520 56430 53560
rect 60020 54880 61420 54920
rect 60020 53560 60060 54880
rect 61380 53560 61420 54880
rect 60020 53520 61420 53560
rect 65010 54880 66410 54920
rect 65010 53560 65050 54880
rect 66370 53560 66410 54880
rect 65010 53520 66410 53560
rect 70000 54880 71400 54920
rect 70000 53560 70040 54880
rect 71360 53560 71400 54880
rect 70000 53520 71400 53560
rect 74990 54880 76390 54920
rect 74990 53560 75030 54880
rect 76350 53560 76390 54880
rect 74990 53520 76390 53560
rect 140 53170 1540 53210
rect 140 51850 180 53170
rect 1500 51850 1540 53170
rect 140 51810 1540 51850
rect 5130 53170 6530 53210
rect 5130 51850 5170 53170
rect 6490 51850 6530 53170
rect 5130 51810 6530 51850
rect 10120 53170 11520 53210
rect 10120 51850 10160 53170
rect 11480 51850 11520 53170
rect 10120 51810 11520 51850
rect 15110 53170 16510 53210
rect 15110 51850 15150 53170
rect 16470 51850 16510 53170
rect 15110 51810 16510 51850
rect 20100 53170 21500 53210
rect 20100 51850 20140 53170
rect 21460 51850 21500 53170
rect 20100 51810 21500 51850
rect 25090 53170 26490 53210
rect 25090 51850 25130 53170
rect 26450 51850 26490 53170
rect 25090 51810 26490 51850
rect 30080 53170 31480 53210
rect 30080 51850 30120 53170
rect 31440 51850 31480 53170
rect 30080 51810 31480 51850
rect 35070 53170 36470 53210
rect 35070 51850 35110 53170
rect 36430 51850 36470 53170
rect 35070 51810 36470 51850
rect 40060 53170 41460 53210
rect 40060 51850 40100 53170
rect 41420 51850 41460 53170
rect 40060 51810 41460 51850
rect 45050 53170 46450 53210
rect 45050 51850 45090 53170
rect 46410 51850 46450 53170
rect 45050 51810 46450 51850
rect 50040 53170 51440 53210
rect 50040 51850 50080 53170
rect 51400 51850 51440 53170
rect 50040 51810 51440 51850
rect 55030 53170 56430 53210
rect 55030 51850 55070 53170
rect 56390 51850 56430 53170
rect 55030 51810 56430 51850
rect 60020 53170 61420 53210
rect 60020 51850 60060 53170
rect 61380 51850 61420 53170
rect 60020 51810 61420 51850
rect 65010 53170 66410 53210
rect 65010 51850 65050 53170
rect 66370 51850 66410 53170
rect 65010 51810 66410 51850
rect 70000 53170 71400 53210
rect 70000 51850 70040 53170
rect 71360 51850 71400 53170
rect 70000 51810 71400 51850
rect 74990 53170 76390 53210
rect 74990 51850 75030 53170
rect 76350 51850 76390 53170
rect 74990 51810 76390 51850
rect 140 51460 1540 51500
rect 140 50140 180 51460
rect 1500 50140 1540 51460
rect 140 50100 1540 50140
rect 5130 51460 6530 51500
rect 5130 50140 5170 51460
rect 6490 50140 6530 51460
rect 5130 50100 6530 50140
rect 10120 51460 11520 51500
rect 10120 50140 10160 51460
rect 11480 50140 11520 51460
rect 10120 50100 11520 50140
rect 15110 51460 16510 51500
rect 15110 50140 15150 51460
rect 16470 50140 16510 51460
rect 15110 50100 16510 50140
rect 20100 51460 21500 51500
rect 20100 50140 20140 51460
rect 21460 50140 21500 51460
rect 20100 50100 21500 50140
rect 25090 51460 26490 51500
rect 25090 50140 25130 51460
rect 26450 50140 26490 51460
rect 25090 50100 26490 50140
rect 30080 51460 31480 51500
rect 30080 50140 30120 51460
rect 31440 50140 31480 51460
rect 30080 50100 31480 50140
rect 35070 51460 36470 51500
rect 35070 50140 35110 51460
rect 36430 50140 36470 51460
rect 35070 50100 36470 50140
rect 40060 51460 41460 51500
rect 40060 50140 40100 51460
rect 41420 50140 41460 51460
rect 40060 50100 41460 50140
rect 45050 51460 46450 51500
rect 45050 50140 45090 51460
rect 46410 50140 46450 51460
rect 45050 50100 46450 50140
rect 50040 51460 51440 51500
rect 50040 50140 50080 51460
rect 51400 50140 51440 51460
rect 50040 50100 51440 50140
rect 55030 51460 56430 51500
rect 55030 50140 55070 51460
rect 56390 50140 56430 51460
rect 55030 50100 56430 50140
rect 60020 51460 61420 51500
rect 60020 50140 60060 51460
rect 61380 50140 61420 51460
rect 60020 50100 61420 50140
rect 65010 51460 66410 51500
rect 65010 50140 65050 51460
rect 66370 50140 66410 51460
rect 65010 50100 66410 50140
rect 70000 51460 71400 51500
rect 70000 50140 70040 51460
rect 71360 50140 71400 51460
rect 70000 50100 71400 50140
rect 74990 51460 76390 51500
rect 74990 50140 75030 51460
rect 76350 50140 76390 51460
rect 74990 50100 76390 50140
rect 140 49750 1540 49790
rect 140 48430 180 49750
rect 1500 48430 1540 49750
rect 140 48390 1540 48430
rect 5130 49750 6530 49790
rect 5130 48430 5170 49750
rect 6490 48430 6530 49750
rect 5130 48390 6530 48430
rect 10120 49750 11520 49790
rect 10120 48430 10160 49750
rect 11480 48430 11520 49750
rect 10120 48390 11520 48430
rect 15110 49750 16510 49790
rect 15110 48430 15150 49750
rect 16470 48430 16510 49750
rect 15110 48390 16510 48430
rect 20100 49750 21500 49790
rect 20100 48430 20140 49750
rect 21460 48430 21500 49750
rect 20100 48390 21500 48430
rect 25090 49750 26490 49790
rect 25090 48430 25130 49750
rect 26450 48430 26490 49750
rect 25090 48390 26490 48430
rect 30080 49750 31480 49790
rect 30080 48430 30120 49750
rect 31440 48430 31480 49750
rect 30080 48390 31480 48430
rect 35070 49750 36470 49790
rect 35070 48430 35110 49750
rect 36430 48430 36470 49750
rect 35070 48390 36470 48430
rect 40060 49750 41460 49790
rect 40060 48430 40100 49750
rect 41420 48430 41460 49750
rect 40060 48390 41460 48430
rect 45050 49750 46450 49790
rect 45050 48430 45090 49750
rect 46410 48430 46450 49750
rect 45050 48390 46450 48430
rect 50040 49750 51440 49790
rect 50040 48430 50080 49750
rect 51400 48430 51440 49750
rect 50040 48390 51440 48430
rect 55030 49750 56430 49790
rect 55030 48430 55070 49750
rect 56390 48430 56430 49750
rect 55030 48390 56430 48430
rect 60020 49750 61420 49790
rect 60020 48430 60060 49750
rect 61380 48430 61420 49750
rect 60020 48390 61420 48430
rect 65010 49750 66410 49790
rect 65010 48430 65050 49750
rect 66370 48430 66410 49750
rect 65010 48390 66410 48430
rect 70000 49750 71400 49790
rect 70000 48430 70040 49750
rect 71360 48430 71400 49750
rect 70000 48390 71400 48430
rect 74990 49750 76390 49790
rect 74990 48430 75030 49750
rect 76350 48430 76390 49750
rect 74990 48390 76390 48430
rect 140 48040 1540 48080
rect 140 46720 180 48040
rect 1500 46720 1540 48040
rect 140 46680 1540 46720
rect 5130 48040 6530 48080
rect 5130 46720 5170 48040
rect 6490 46720 6530 48040
rect 5130 46680 6530 46720
rect 10120 48040 11520 48080
rect 10120 46720 10160 48040
rect 11480 46720 11520 48040
rect 10120 46680 11520 46720
rect 15110 48040 16510 48080
rect 15110 46720 15150 48040
rect 16470 46720 16510 48040
rect 15110 46680 16510 46720
rect 20100 48040 21500 48080
rect 20100 46720 20140 48040
rect 21460 46720 21500 48040
rect 20100 46680 21500 46720
rect 25090 48040 26490 48080
rect 25090 46720 25130 48040
rect 26450 46720 26490 48040
rect 25090 46680 26490 46720
rect 30080 48040 31480 48080
rect 30080 46720 30120 48040
rect 31440 46720 31480 48040
rect 30080 46680 31480 46720
rect 35070 48040 36470 48080
rect 35070 46720 35110 48040
rect 36430 46720 36470 48040
rect 35070 46680 36470 46720
rect 40060 48040 41460 48080
rect 40060 46720 40100 48040
rect 41420 46720 41460 48040
rect 40060 46680 41460 46720
rect 45050 48040 46450 48080
rect 45050 46720 45090 48040
rect 46410 46720 46450 48040
rect 45050 46680 46450 46720
rect 50040 48040 51440 48080
rect 50040 46720 50080 48040
rect 51400 46720 51440 48040
rect 50040 46680 51440 46720
rect 55030 48040 56430 48080
rect 55030 46720 55070 48040
rect 56390 46720 56430 48040
rect 55030 46680 56430 46720
rect 60020 48040 61420 48080
rect 60020 46720 60060 48040
rect 61380 46720 61420 48040
rect 60020 46680 61420 46720
rect 65010 48040 66410 48080
rect 65010 46720 65050 48040
rect 66370 46720 66410 48040
rect 65010 46680 66410 46720
rect 70000 48040 71400 48080
rect 70000 46720 70040 48040
rect 71360 46720 71400 48040
rect 70000 46680 71400 46720
rect 74990 48040 76390 48080
rect 74990 46720 75030 48040
rect 76350 46720 76390 48040
rect 74990 46680 76390 46720
rect 140 46330 1540 46370
rect 140 45010 180 46330
rect 1500 45010 1540 46330
rect 140 44970 1540 45010
rect 5130 46330 6530 46370
rect 5130 45010 5170 46330
rect 6490 45010 6530 46330
rect 5130 44970 6530 45010
rect 10120 46330 11520 46370
rect 10120 45010 10160 46330
rect 11480 45010 11520 46330
rect 10120 44970 11520 45010
rect 15110 46330 16510 46370
rect 15110 45010 15150 46330
rect 16470 45010 16510 46330
rect 15110 44970 16510 45010
rect 20100 46330 21500 46370
rect 20100 45010 20140 46330
rect 21460 45010 21500 46330
rect 20100 44970 21500 45010
rect 25090 46330 26490 46370
rect 25090 45010 25130 46330
rect 26450 45010 26490 46330
rect 25090 44970 26490 45010
rect 30080 46330 31480 46370
rect 30080 45010 30120 46330
rect 31440 45010 31480 46330
rect 30080 44970 31480 45010
rect 35070 46330 36470 46370
rect 35070 45010 35110 46330
rect 36430 45010 36470 46330
rect 35070 44970 36470 45010
rect 40060 46330 41460 46370
rect 40060 45010 40100 46330
rect 41420 45010 41460 46330
rect 40060 44970 41460 45010
rect 45050 46330 46450 46370
rect 45050 45010 45090 46330
rect 46410 45010 46450 46330
rect 45050 44970 46450 45010
rect 50040 46330 51440 46370
rect 50040 45010 50080 46330
rect 51400 45010 51440 46330
rect 50040 44970 51440 45010
rect 55030 46330 56430 46370
rect 55030 45010 55070 46330
rect 56390 45010 56430 46330
rect 55030 44970 56430 45010
rect 60020 46330 61420 46370
rect 60020 45010 60060 46330
rect 61380 45010 61420 46330
rect 60020 44970 61420 45010
rect 65010 46330 66410 46370
rect 65010 45010 65050 46330
rect 66370 45010 66410 46330
rect 65010 44970 66410 45010
rect 70000 46330 71400 46370
rect 70000 45010 70040 46330
rect 71360 45010 71400 46330
rect 70000 44970 71400 45010
rect 74990 46330 76390 46370
rect 74990 45010 75030 46330
rect 76350 45010 76390 46330
rect 74990 44970 76390 45010
rect 140 44620 1540 44660
rect 140 43300 180 44620
rect 1500 43300 1540 44620
rect 140 43260 1540 43300
rect 5130 44620 6530 44660
rect 5130 43300 5170 44620
rect 6490 43300 6530 44620
rect 5130 43260 6530 43300
rect 10120 44620 11520 44660
rect 10120 43300 10160 44620
rect 11480 43300 11520 44620
rect 10120 43260 11520 43300
rect 15110 44620 16510 44660
rect 15110 43300 15150 44620
rect 16470 43300 16510 44620
rect 15110 43260 16510 43300
rect 20100 44620 21500 44660
rect 20100 43300 20140 44620
rect 21460 43300 21500 44620
rect 20100 43260 21500 43300
rect 25090 44620 26490 44660
rect 25090 43300 25130 44620
rect 26450 43300 26490 44620
rect 25090 43260 26490 43300
rect 30080 44620 31480 44660
rect 30080 43300 30120 44620
rect 31440 43300 31480 44620
rect 30080 43260 31480 43300
rect 35070 44620 36470 44660
rect 35070 43300 35110 44620
rect 36430 43300 36470 44620
rect 35070 43260 36470 43300
rect 40060 44620 41460 44660
rect 40060 43300 40100 44620
rect 41420 43300 41460 44620
rect 40060 43260 41460 43300
rect 45050 44620 46450 44660
rect 45050 43300 45090 44620
rect 46410 43300 46450 44620
rect 45050 43260 46450 43300
rect 50040 44620 51440 44660
rect 50040 43300 50080 44620
rect 51400 43300 51440 44620
rect 50040 43260 51440 43300
rect 55030 44620 56430 44660
rect 55030 43300 55070 44620
rect 56390 43300 56430 44620
rect 55030 43260 56430 43300
rect 60020 44620 61420 44660
rect 60020 43300 60060 44620
rect 61380 43300 61420 44620
rect 60020 43260 61420 43300
rect 65010 44620 66410 44660
rect 65010 43300 65050 44620
rect 66370 43300 66410 44620
rect 65010 43260 66410 43300
rect 70000 44620 71400 44660
rect 70000 43300 70040 44620
rect 71360 43300 71400 44620
rect 70000 43260 71400 43300
rect 74990 44620 76390 44660
rect 74990 43300 75030 44620
rect 76350 43300 76390 44620
rect 74990 43260 76390 43300
rect 140 42910 1540 42950
rect 140 41590 180 42910
rect 1500 41590 1540 42910
rect 140 41550 1540 41590
rect 5130 42910 6530 42950
rect 5130 41590 5170 42910
rect 6490 41590 6530 42910
rect 5130 41550 6530 41590
rect 10120 42910 11520 42950
rect 10120 41590 10160 42910
rect 11480 41590 11520 42910
rect 10120 41550 11520 41590
rect 15110 42910 16510 42950
rect 15110 41590 15150 42910
rect 16470 41590 16510 42910
rect 15110 41550 16510 41590
rect 20100 42910 21500 42950
rect 20100 41590 20140 42910
rect 21460 41590 21500 42910
rect 20100 41550 21500 41590
rect 25090 42910 26490 42950
rect 25090 41590 25130 42910
rect 26450 41590 26490 42910
rect 25090 41550 26490 41590
rect 30080 42910 31480 42950
rect 30080 41590 30120 42910
rect 31440 41590 31480 42910
rect 30080 41550 31480 41590
rect 35070 42910 36470 42950
rect 35070 41590 35110 42910
rect 36430 41590 36470 42910
rect 35070 41550 36470 41590
rect 40060 42910 41460 42950
rect 40060 41590 40100 42910
rect 41420 41590 41460 42910
rect 40060 41550 41460 41590
rect 45050 42910 46450 42950
rect 45050 41590 45090 42910
rect 46410 41590 46450 42910
rect 45050 41550 46450 41590
rect 50040 42910 51440 42950
rect 50040 41590 50080 42910
rect 51400 41590 51440 42910
rect 50040 41550 51440 41590
rect 55030 42910 56430 42950
rect 55030 41590 55070 42910
rect 56390 41590 56430 42910
rect 55030 41550 56430 41590
rect 60020 42910 61420 42950
rect 60020 41590 60060 42910
rect 61380 41590 61420 42910
rect 60020 41550 61420 41590
rect 65010 42910 66410 42950
rect 65010 41590 65050 42910
rect 66370 41590 66410 42910
rect 65010 41550 66410 41590
rect 70000 42910 71400 42950
rect 70000 41590 70040 42910
rect 71360 41590 71400 42910
rect 70000 41550 71400 41590
rect 74990 42910 76390 42950
rect 74990 41590 75030 42910
rect 76350 41590 76390 42910
rect 74990 41550 76390 41590
rect 140 41200 1540 41240
rect 140 39880 180 41200
rect 1500 39880 1540 41200
rect 140 39840 1540 39880
rect 5130 41200 6530 41240
rect 5130 39880 5170 41200
rect 6490 39880 6530 41200
rect 5130 39840 6530 39880
rect 10120 41200 11520 41240
rect 10120 39880 10160 41200
rect 11480 39880 11520 41200
rect 10120 39840 11520 39880
rect 15110 41200 16510 41240
rect 15110 39880 15150 41200
rect 16470 39880 16510 41200
rect 15110 39840 16510 39880
rect 20100 41200 21500 41240
rect 20100 39880 20140 41200
rect 21460 39880 21500 41200
rect 20100 39840 21500 39880
rect 25090 41200 26490 41240
rect 25090 39880 25130 41200
rect 26450 39880 26490 41200
rect 25090 39840 26490 39880
rect 30080 41200 31480 41240
rect 30080 39880 30120 41200
rect 31440 39880 31480 41200
rect 30080 39840 31480 39880
rect 35070 41200 36470 41240
rect 35070 39880 35110 41200
rect 36430 39880 36470 41200
rect 35070 39840 36470 39880
rect 40060 41200 41460 41240
rect 40060 39880 40100 41200
rect 41420 39880 41460 41200
rect 40060 39840 41460 39880
rect 45050 41200 46450 41240
rect 45050 39880 45090 41200
rect 46410 39880 46450 41200
rect 45050 39840 46450 39880
rect 50040 41200 51440 41240
rect 50040 39880 50080 41200
rect 51400 39880 51440 41200
rect 50040 39840 51440 39880
rect 55030 41200 56430 41240
rect 55030 39880 55070 41200
rect 56390 39880 56430 41200
rect 55030 39840 56430 39880
rect 60020 41200 61420 41240
rect 60020 39880 60060 41200
rect 61380 39880 61420 41200
rect 60020 39840 61420 39880
rect 65010 41200 66410 41240
rect 65010 39880 65050 41200
rect 66370 39880 66410 41200
rect 65010 39840 66410 39880
rect 70000 41200 71400 41240
rect 70000 39880 70040 41200
rect 71360 39880 71400 41200
rect 70000 39840 71400 39880
rect 74990 41200 76390 41240
rect 74990 39880 75030 41200
rect 76350 39880 76390 41200
rect 74990 39840 76390 39880
<< mimcapcontact >>
rect 180 65530 1500 66850
rect 5170 65530 6490 66850
rect 10160 65530 11480 66850
rect 15150 65530 16470 66850
rect 20140 65530 21460 66850
rect 25130 65530 26450 66850
rect 30120 65530 31440 66850
rect 35110 65530 36430 66850
rect 40100 65530 41420 66850
rect 45090 65530 46410 66850
rect 50080 65530 51400 66850
rect 55070 65530 56390 66850
rect 60060 65530 61380 66850
rect 65050 65530 66370 66850
rect 70040 65530 71360 66850
rect 75030 65530 76350 66850
rect 180 63820 1500 65140
rect 5170 63820 6490 65140
rect 10160 63820 11480 65140
rect 15150 63820 16470 65140
rect 20140 63820 21460 65140
rect 25130 63820 26450 65140
rect 30120 63820 31440 65140
rect 35110 63820 36430 65140
rect 40100 63820 41420 65140
rect 45090 63820 46410 65140
rect 50080 63820 51400 65140
rect 55070 63820 56390 65140
rect 60060 63820 61380 65140
rect 65050 63820 66370 65140
rect 70040 63820 71360 65140
rect 75030 63820 76350 65140
rect 180 62110 1500 63430
rect 5170 62110 6490 63430
rect 10160 62110 11480 63430
rect 15150 62110 16470 63430
rect 20140 62110 21460 63430
rect 25130 62110 26450 63430
rect 30120 62110 31440 63430
rect 35110 62110 36430 63430
rect 40100 62110 41420 63430
rect 45090 62110 46410 63430
rect 50080 62110 51400 63430
rect 55070 62110 56390 63430
rect 60060 62110 61380 63430
rect 65050 62110 66370 63430
rect 70040 62110 71360 63430
rect 75030 62110 76350 63430
rect 180 60400 1500 61720
rect 5170 60400 6490 61720
rect 10160 60400 11480 61720
rect 15150 60400 16470 61720
rect 20140 60400 21460 61720
rect 25130 60400 26450 61720
rect 30120 60400 31440 61720
rect 35110 60400 36430 61720
rect 40100 60400 41420 61720
rect 45090 60400 46410 61720
rect 50080 60400 51400 61720
rect 55070 60400 56390 61720
rect 60060 60400 61380 61720
rect 65050 60400 66370 61720
rect 70040 60400 71360 61720
rect 75030 60400 76350 61720
rect 180 58690 1500 60010
rect 5170 58690 6490 60010
rect 10160 58690 11480 60010
rect 15150 58690 16470 60010
rect 20140 58690 21460 60010
rect 25130 58690 26450 60010
rect 30120 58690 31440 60010
rect 35110 58690 36430 60010
rect 40100 58690 41420 60010
rect 45090 58690 46410 60010
rect 50080 58690 51400 60010
rect 55070 58690 56390 60010
rect 60060 58690 61380 60010
rect 65050 58690 66370 60010
rect 70040 58690 71360 60010
rect 75030 58690 76350 60010
rect 180 56980 1500 58300
rect 5170 56980 6490 58300
rect 10160 56980 11480 58300
rect 15150 56980 16470 58300
rect 20140 56980 21460 58300
rect 25130 56980 26450 58300
rect 30120 56980 31440 58300
rect 35110 56980 36430 58300
rect 40100 56980 41420 58300
rect 45090 56980 46410 58300
rect 50080 56980 51400 58300
rect 55070 56980 56390 58300
rect 60060 56980 61380 58300
rect 65050 56980 66370 58300
rect 70040 56980 71360 58300
rect 75030 56980 76350 58300
rect 180 55270 1500 56590
rect 5170 55270 6490 56590
rect 10160 55270 11480 56590
rect 15150 55270 16470 56590
rect 20140 55270 21460 56590
rect 25130 55270 26450 56590
rect 30120 55270 31440 56590
rect 35110 55270 36430 56590
rect 40100 55270 41420 56590
rect 45090 55270 46410 56590
rect 50080 55270 51400 56590
rect 55070 55270 56390 56590
rect 60060 55270 61380 56590
rect 65050 55270 66370 56590
rect 70040 55270 71360 56590
rect 75030 55270 76350 56590
rect 180 53560 1500 54880
rect 5170 53560 6490 54880
rect 10160 53560 11480 54880
rect 15150 53560 16470 54880
rect 20140 53560 21460 54880
rect 25130 53560 26450 54880
rect 30120 53560 31440 54880
rect 35110 53560 36430 54880
rect 40100 53560 41420 54880
rect 45090 53560 46410 54880
rect 50080 53560 51400 54880
rect 55070 53560 56390 54880
rect 60060 53560 61380 54880
rect 65050 53560 66370 54880
rect 70040 53560 71360 54880
rect 75030 53560 76350 54880
rect 180 51850 1500 53170
rect 5170 51850 6490 53170
rect 10160 51850 11480 53170
rect 15150 51850 16470 53170
rect 20140 51850 21460 53170
rect 25130 51850 26450 53170
rect 30120 51850 31440 53170
rect 35110 51850 36430 53170
rect 40100 51850 41420 53170
rect 45090 51850 46410 53170
rect 50080 51850 51400 53170
rect 55070 51850 56390 53170
rect 60060 51850 61380 53170
rect 65050 51850 66370 53170
rect 70040 51850 71360 53170
rect 75030 51850 76350 53170
rect 180 50140 1500 51460
rect 5170 50140 6490 51460
rect 10160 50140 11480 51460
rect 15150 50140 16470 51460
rect 20140 50140 21460 51460
rect 25130 50140 26450 51460
rect 30120 50140 31440 51460
rect 35110 50140 36430 51460
rect 40100 50140 41420 51460
rect 45090 50140 46410 51460
rect 50080 50140 51400 51460
rect 55070 50140 56390 51460
rect 60060 50140 61380 51460
rect 65050 50140 66370 51460
rect 70040 50140 71360 51460
rect 75030 50140 76350 51460
rect 180 48430 1500 49750
rect 5170 48430 6490 49750
rect 10160 48430 11480 49750
rect 15150 48430 16470 49750
rect 20140 48430 21460 49750
rect 25130 48430 26450 49750
rect 30120 48430 31440 49750
rect 35110 48430 36430 49750
rect 40100 48430 41420 49750
rect 45090 48430 46410 49750
rect 50080 48430 51400 49750
rect 55070 48430 56390 49750
rect 60060 48430 61380 49750
rect 65050 48430 66370 49750
rect 70040 48430 71360 49750
rect 75030 48430 76350 49750
rect 180 46720 1500 48040
rect 5170 46720 6490 48040
rect 10160 46720 11480 48040
rect 15150 46720 16470 48040
rect 20140 46720 21460 48040
rect 25130 46720 26450 48040
rect 30120 46720 31440 48040
rect 35110 46720 36430 48040
rect 40100 46720 41420 48040
rect 45090 46720 46410 48040
rect 50080 46720 51400 48040
rect 55070 46720 56390 48040
rect 60060 46720 61380 48040
rect 65050 46720 66370 48040
rect 70040 46720 71360 48040
rect 75030 46720 76350 48040
rect 180 45010 1500 46330
rect 5170 45010 6490 46330
rect 10160 45010 11480 46330
rect 15150 45010 16470 46330
rect 20140 45010 21460 46330
rect 25130 45010 26450 46330
rect 30120 45010 31440 46330
rect 35110 45010 36430 46330
rect 40100 45010 41420 46330
rect 45090 45010 46410 46330
rect 50080 45010 51400 46330
rect 55070 45010 56390 46330
rect 60060 45010 61380 46330
rect 65050 45010 66370 46330
rect 70040 45010 71360 46330
rect 75030 45010 76350 46330
rect 180 43300 1500 44620
rect 5170 43300 6490 44620
rect 10160 43300 11480 44620
rect 15150 43300 16470 44620
rect 20140 43300 21460 44620
rect 25130 43300 26450 44620
rect 30120 43300 31440 44620
rect 35110 43300 36430 44620
rect 40100 43300 41420 44620
rect 45090 43300 46410 44620
rect 50080 43300 51400 44620
rect 55070 43300 56390 44620
rect 60060 43300 61380 44620
rect 65050 43300 66370 44620
rect 70040 43300 71360 44620
rect 75030 43300 76350 44620
rect 180 41590 1500 42910
rect 5170 41590 6490 42910
rect 10160 41590 11480 42910
rect 15150 41590 16470 42910
rect 20140 41590 21460 42910
rect 25130 41590 26450 42910
rect 30120 41590 31440 42910
rect 35110 41590 36430 42910
rect 40100 41590 41420 42910
rect 45090 41590 46410 42910
rect 50080 41590 51400 42910
rect 55070 41590 56390 42910
rect 60060 41590 61380 42910
rect 65050 41590 66370 42910
rect 70040 41590 71360 42910
rect 75030 41590 76350 42910
rect 180 39880 1500 41200
rect 5170 39880 6490 41200
rect 10160 39880 11480 41200
rect 15150 39880 16470 41200
rect 20140 39880 21460 41200
rect 25130 39880 26450 41200
rect 30120 39880 31440 41200
rect 35110 39880 36430 41200
rect 40100 39880 41420 41200
rect 45090 39880 46410 41200
rect 50080 39880 51400 41200
rect 55070 39880 56390 41200
rect 60060 39880 61380 41200
rect 65050 39880 66370 41200
rect 70040 39880 71360 41200
rect 75030 39880 76350 41200
<< metal4 >>
rect 100 67110 79670 67170
rect 180 66851 240 67110
rect 1772 66902 1868 66918
rect 179 66850 1501 66851
rect 179 65530 180 66850
rect 1500 65530 1501 66850
rect 179 65529 1501 65530
rect 180 65141 240 65529
rect 1772 65478 1788 66902
rect 1852 66220 1868 66902
rect 5170 66851 5230 67110
rect 6762 66902 6858 66918
rect 5169 66850 6491 66851
rect 3240 66280 3380 66310
rect 3240 66220 3270 66280
rect 1852 66210 3270 66220
rect 3350 66210 3380 66280
rect 1852 66170 3380 66210
rect 1852 66160 3270 66170
rect 1852 65478 1868 66160
rect 3240 66100 3270 66160
rect 3350 66100 3380 66170
rect 3240 66060 3380 66100
rect 5169 65530 5170 66850
rect 6490 65530 6491 66850
rect 5169 65529 6491 65530
rect 1772 65462 1868 65478
rect 1772 65192 1868 65208
rect 179 65140 1501 65141
rect 179 63820 180 65140
rect 1500 63820 1501 65140
rect 179 63819 1501 63820
rect 180 63431 240 63819
rect 1772 63768 1788 65192
rect 1852 64510 1868 65192
rect 5170 65141 5230 65529
rect 6762 65478 6778 66902
rect 6842 66220 6858 66902
rect 10160 66851 10220 67110
rect 11752 66902 11848 66918
rect 10159 66850 11481 66851
rect 8230 66280 8370 66310
rect 8230 66220 8260 66280
rect 6842 66210 8260 66220
rect 8340 66210 8370 66280
rect 6842 66170 8370 66210
rect 6842 66160 8260 66170
rect 6842 65478 6858 66160
rect 8230 66100 8260 66160
rect 8340 66100 8370 66170
rect 8230 66060 8370 66100
rect 10159 65530 10160 66850
rect 11480 65530 11481 66850
rect 10159 65529 11481 65530
rect 6762 65462 6858 65478
rect 6762 65192 6858 65208
rect 5169 65140 6491 65141
rect 3240 64570 3380 64600
rect 3240 64510 3270 64570
rect 1852 64500 3270 64510
rect 3350 64500 3380 64570
rect 1852 64460 3380 64500
rect 1852 64450 3270 64460
rect 1852 63768 1868 64450
rect 3240 64390 3270 64450
rect 3350 64390 3380 64460
rect 3240 64350 3380 64390
rect 5169 63820 5170 65140
rect 6490 63820 6491 65140
rect 5169 63819 6491 63820
rect 1772 63752 1868 63768
rect 1772 63482 1868 63498
rect 179 63430 1501 63431
rect 179 62110 180 63430
rect 1500 62110 1501 63430
rect 179 62109 1501 62110
rect 180 61721 240 62109
rect 1772 62058 1788 63482
rect 1852 62800 1868 63482
rect 5170 63431 5230 63819
rect 6762 63768 6778 65192
rect 6842 64510 6858 65192
rect 10160 65141 10220 65529
rect 11752 65478 11768 66902
rect 11832 66220 11848 66902
rect 15150 66851 15210 67110
rect 16742 66902 16838 66918
rect 15149 66850 16471 66851
rect 13220 66280 13360 66310
rect 13220 66220 13250 66280
rect 11832 66210 13250 66220
rect 13330 66210 13360 66280
rect 11832 66170 13360 66210
rect 11832 66160 13250 66170
rect 11832 65478 11848 66160
rect 13220 66100 13250 66160
rect 13330 66100 13360 66170
rect 13220 66060 13360 66100
rect 15149 65530 15150 66850
rect 16470 65530 16471 66850
rect 15149 65529 16471 65530
rect 11752 65462 11848 65478
rect 11752 65192 11848 65208
rect 10159 65140 11481 65141
rect 8230 64570 8370 64600
rect 8230 64510 8260 64570
rect 6842 64500 8260 64510
rect 8340 64500 8370 64570
rect 6842 64460 8370 64500
rect 6842 64450 8260 64460
rect 6842 63768 6858 64450
rect 8230 64390 8260 64450
rect 8340 64390 8370 64460
rect 8230 64350 8370 64390
rect 10159 63820 10160 65140
rect 11480 63820 11481 65140
rect 10159 63819 11481 63820
rect 6762 63752 6858 63768
rect 6762 63482 6858 63498
rect 5169 63430 6491 63431
rect 3240 62860 3380 62890
rect 3240 62800 3270 62860
rect 1852 62790 3270 62800
rect 3350 62790 3380 62860
rect 1852 62750 3380 62790
rect 1852 62740 3270 62750
rect 1852 62058 1868 62740
rect 3240 62680 3270 62740
rect 3350 62680 3380 62750
rect 3240 62640 3380 62680
rect 5169 62110 5170 63430
rect 6490 62110 6491 63430
rect 5169 62109 6491 62110
rect 1772 62042 1868 62058
rect 1772 61772 1868 61788
rect 179 61720 1501 61721
rect 179 60400 180 61720
rect 1500 60400 1501 61720
rect 179 60399 1501 60400
rect 180 60011 240 60399
rect 1772 60348 1788 61772
rect 1852 61090 1868 61772
rect 5170 61721 5230 62109
rect 6762 62058 6778 63482
rect 6842 62800 6858 63482
rect 10160 63431 10220 63819
rect 11752 63768 11768 65192
rect 11832 64510 11848 65192
rect 15150 65141 15210 65529
rect 16742 65478 16758 66902
rect 16822 66220 16838 66902
rect 20140 66851 20200 67110
rect 21732 66902 21828 66918
rect 20139 66850 21461 66851
rect 18210 66280 18350 66310
rect 18210 66220 18240 66280
rect 16822 66210 18240 66220
rect 18320 66210 18350 66280
rect 16822 66170 18350 66210
rect 16822 66160 18240 66170
rect 16822 65478 16838 66160
rect 18210 66100 18240 66160
rect 18320 66100 18350 66170
rect 18210 66060 18350 66100
rect 20139 65530 20140 66850
rect 21460 65530 21461 66850
rect 20139 65529 21461 65530
rect 16742 65462 16838 65478
rect 16742 65192 16838 65208
rect 15149 65140 16471 65141
rect 13220 64570 13360 64600
rect 13220 64510 13250 64570
rect 11832 64500 13250 64510
rect 13330 64500 13360 64570
rect 11832 64460 13360 64500
rect 11832 64450 13250 64460
rect 11832 63768 11848 64450
rect 13220 64390 13250 64450
rect 13330 64390 13360 64460
rect 13220 64350 13360 64390
rect 15149 63820 15150 65140
rect 16470 63820 16471 65140
rect 15149 63819 16471 63820
rect 11752 63752 11848 63768
rect 11752 63482 11848 63498
rect 10159 63430 11481 63431
rect 8230 62860 8370 62890
rect 8230 62800 8260 62860
rect 6842 62790 8260 62800
rect 8340 62790 8370 62860
rect 6842 62750 8370 62790
rect 6842 62740 8260 62750
rect 6842 62058 6858 62740
rect 8230 62680 8260 62740
rect 8340 62680 8370 62750
rect 8230 62640 8370 62680
rect 10159 62110 10160 63430
rect 11480 62110 11481 63430
rect 10159 62109 11481 62110
rect 6762 62042 6858 62058
rect 6762 61772 6858 61788
rect 5169 61720 6491 61721
rect 3240 61150 3380 61180
rect 3240 61090 3270 61150
rect 1852 61080 3270 61090
rect 3350 61080 3380 61150
rect 1852 61040 3380 61080
rect 1852 61030 3270 61040
rect 1852 60348 1868 61030
rect 3240 60970 3270 61030
rect 3350 60970 3380 61040
rect 3240 60930 3380 60970
rect 5169 60400 5170 61720
rect 6490 60400 6491 61720
rect 5169 60399 6491 60400
rect 1772 60332 1868 60348
rect 1772 60062 1868 60078
rect 179 60010 1501 60011
rect 179 58690 180 60010
rect 1500 58690 1501 60010
rect 179 58689 1501 58690
rect 180 58301 240 58689
rect 1772 58638 1788 60062
rect 1852 59380 1868 60062
rect 5170 60011 5230 60399
rect 6762 60348 6778 61772
rect 6842 61090 6858 61772
rect 10160 61721 10220 62109
rect 11752 62058 11768 63482
rect 11832 62800 11848 63482
rect 15150 63431 15210 63819
rect 16742 63768 16758 65192
rect 16822 64510 16838 65192
rect 20140 65141 20200 65529
rect 21732 65478 21748 66902
rect 21812 66220 21828 66902
rect 25130 66851 25190 67110
rect 26722 66902 26818 66918
rect 25129 66850 26451 66851
rect 23200 66280 23340 66310
rect 23200 66220 23230 66280
rect 21812 66210 23230 66220
rect 23310 66210 23340 66280
rect 21812 66170 23340 66210
rect 21812 66160 23230 66170
rect 21812 65478 21828 66160
rect 23200 66100 23230 66160
rect 23310 66100 23340 66170
rect 23200 66060 23340 66100
rect 25129 65530 25130 66850
rect 26450 65530 26451 66850
rect 25129 65529 26451 65530
rect 21732 65462 21828 65478
rect 21732 65192 21828 65208
rect 20139 65140 21461 65141
rect 18210 64570 18350 64600
rect 18210 64510 18240 64570
rect 16822 64500 18240 64510
rect 18320 64500 18350 64570
rect 16822 64460 18350 64500
rect 16822 64450 18240 64460
rect 16822 63768 16838 64450
rect 18210 64390 18240 64450
rect 18320 64390 18350 64460
rect 18210 64350 18350 64390
rect 20139 63820 20140 65140
rect 21460 63820 21461 65140
rect 20139 63819 21461 63820
rect 16742 63752 16838 63768
rect 16742 63482 16838 63498
rect 15149 63430 16471 63431
rect 13220 62860 13360 62890
rect 13220 62800 13250 62860
rect 11832 62790 13250 62800
rect 13330 62790 13360 62860
rect 11832 62750 13360 62790
rect 11832 62740 13250 62750
rect 11832 62058 11848 62740
rect 13220 62680 13250 62740
rect 13330 62680 13360 62750
rect 13220 62640 13360 62680
rect 15149 62110 15150 63430
rect 16470 62110 16471 63430
rect 15149 62109 16471 62110
rect 11752 62042 11848 62058
rect 11752 61772 11848 61788
rect 10159 61720 11481 61721
rect 8230 61150 8370 61180
rect 8230 61090 8260 61150
rect 6842 61080 8260 61090
rect 8340 61080 8370 61150
rect 6842 61040 8370 61080
rect 6842 61030 8260 61040
rect 6842 60348 6858 61030
rect 8230 60970 8260 61030
rect 8340 60970 8370 61040
rect 8230 60930 8370 60970
rect 10159 60400 10160 61720
rect 11480 60400 11481 61720
rect 10159 60399 11481 60400
rect 6762 60332 6858 60348
rect 6762 60062 6858 60078
rect 5169 60010 6491 60011
rect 3240 59440 3380 59470
rect 3240 59380 3270 59440
rect 1852 59370 3270 59380
rect 3350 59370 3380 59440
rect 1852 59330 3380 59370
rect 1852 59320 3270 59330
rect 1852 58638 1868 59320
rect 3240 59260 3270 59320
rect 3350 59260 3380 59330
rect 3240 59220 3380 59260
rect 5169 58690 5170 60010
rect 6490 58690 6491 60010
rect 5169 58689 6491 58690
rect 1772 58622 1868 58638
rect 1772 58352 1868 58368
rect 179 58300 1501 58301
rect 179 56980 180 58300
rect 1500 56980 1501 58300
rect 179 56979 1501 56980
rect 180 56591 240 56979
rect 1772 56928 1788 58352
rect 1852 57670 1868 58352
rect 5170 58301 5230 58689
rect 6762 58638 6778 60062
rect 6842 59380 6858 60062
rect 10160 60011 10220 60399
rect 11752 60348 11768 61772
rect 11832 61090 11848 61772
rect 15150 61721 15210 62109
rect 16742 62058 16758 63482
rect 16822 62800 16838 63482
rect 20140 63431 20200 63819
rect 21732 63768 21748 65192
rect 21812 64510 21828 65192
rect 25130 65141 25190 65529
rect 26722 65478 26738 66902
rect 26802 66220 26818 66902
rect 30120 66851 30180 67110
rect 31712 66902 31808 66918
rect 30119 66850 31441 66851
rect 28190 66280 28330 66310
rect 28190 66220 28220 66280
rect 26802 66210 28220 66220
rect 28300 66210 28330 66280
rect 26802 66170 28330 66210
rect 26802 66160 28220 66170
rect 26802 65478 26818 66160
rect 28190 66100 28220 66160
rect 28300 66100 28330 66170
rect 28190 66060 28330 66100
rect 30119 65530 30120 66850
rect 31440 65530 31441 66850
rect 30119 65529 31441 65530
rect 26722 65462 26818 65478
rect 26722 65192 26818 65208
rect 25129 65140 26451 65141
rect 23200 64570 23340 64600
rect 23200 64510 23230 64570
rect 21812 64500 23230 64510
rect 23310 64500 23340 64570
rect 21812 64460 23340 64500
rect 21812 64450 23230 64460
rect 21812 63768 21828 64450
rect 23200 64390 23230 64450
rect 23310 64390 23340 64460
rect 23200 64350 23340 64390
rect 25129 63820 25130 65140
rect 26450 63820 26451 65140
rect 25129 63819 26451 63820
rect 21732 63752 21828 63768
rect 21732 63482 21828 63498
rect 20139 63430 21461 63431
rect 18210 62860 18350 62890
rect 18210 62800 18240 62860
rect 16822 62790 18240 62800
rect 18320 62790 18350 62860
rect 16822 62750 18350 62790
rect 16822 62740 18240 62750
rect 16822 62058 16838 62740
rect 18210 62680 18240 62740
rect 18320 62680 18350 62750
rect 18210 62640 18350 62680
rect 20139 62110 20140 63430
rect 21460 62110 21461 63430
rect 20139 62109 21461 62110
rect 16742 62042 16838 62058
rect 16742 61772 16838 61788
rect 15149 61720 16471 61721
rect 13220 61150 13360 61180
rect 13220 61090 13250 61150
rect 11832 61080 13250 61090
rect 13330 61080 13360 61150
rect 11832 61040 13360 61080
rect 11832 61030 13250 61040
rect 11832 60348 11848 61030
rect 13220 60970 13250 61030
rect 13330 60970 13360 61040
rect 13220 60930 13360 60970
rect 15149 60400 15150 61720
rect 16470 60400 16471 61720
rect 15149 60399 16471 60400
rect 11752 60332 11848 60348
rect 11752 60062 11848 60078
rect 10159 60010 11481 60011
rect 8230 59440 8370 59470
rect 8230 59380 8260 59440
rect 6842 59370 8260 59380
rect 8340 59370 8370 59440
rect 6842 59330 8370 59370
rect 6842 59320 8260 59330
rect 6842 58638 6858 59320
rect 8230 59260 8260 59320
rect 8340 59260 8370 59330
rect 8230 59220 8370 59260
rect 10159 58690 10160 60010
rect 11480 58690 11481 60010
rect 10159 58689 11481 58690
rect 6762 58622 6858 58638
rect 6762 58352 6858 58368
rect 5169 58300 6491 58301
rect 3240 57730 3380 57760
rect 3240 57670 3270 57730
rect 1852 57660 3270 57670
rect 3350 57660 3380 57730
rect 1852 57620 3380 57660
rect 1852 57610 3270 57620
rect 1852 56928 1868 57610
rect 3240 57550 3270 57610
rect 3350 57550 3380 57620
rect 3240 57510 3380 57550
rect 5169 56980 5170 58300
rect 6490 56980 6491 58300
rect 5169 56979 6491 56980
rect 1772 56912 1868 56928
rect 1772 56642 1868 56658
rect 179 56590 1501 56591
rect 179 55270 180 56590
rect 1500 55270 1501 56590
rect 179 55269 1501 55270
rect 180 54881 240 55269
rect 1772 55218 1788 56642
rect 1852 55960 1868 56642
rect 5170 56591 5230 56979
rect 6762 56928 6778 58352
rect 6842 57670 6858 58352
rect 10160 58301 10220 58689
rect 11752 58638 11768 60062
rect 11832 59380 11848 60062
rect 15150 60011 15210 60399
rect 16742 60348 16758 61772
rect 16822 61090 16838 61772
rect 20140 61721 20200 62109
rect 21732 62058 21748 63482
rect 21812 62800 21828 63482
rect 25130 63431 25190 63819
rect 26722 63768 26738 65192
rect 26802 64510 26818 65192
rect 30120 65141 30180 65529
rect 31712 65478 31728 66902
rect 31792 66220 31808 66902
rect 35110 66851 35170 67110
rect 36702 66902 36798 66918
rect 35109 66850 36431 66851
rect 33180 66280 33320 66310
rect 33180 66220 33210 66280
rect 31792 66210 33210 66220
rect 33290 66210 33320 66280
rect 31792 66170 33320 66210
rect 31792 66160 33210 66170
rect 31792 65478 31808 66160
rect 33180 66100 33210 66160
rect 33290 66100 33320 66170
rect 34010 66160 34700 66220
rect 33180 66060 33320 66100
rect 35109 65530 35110 66850
rect 36430 65530 36431 66850
rect 35109 65529 36431 65530
rect 31712 65462 31808 65478
rect 31712 65192 31808 65208
rect 30119 65140 31441 65141
rect 28190 64570 28330 64600
rect 28190 64510 28220 64570
rect 26802 64500 28220 64510
rect 28300 64500 28330 64570
rect 26802 64460 28330 64500
rect 26802 64450 28220 64460
rect 26802 63768 26818 64450
rect 28190 64390 28220 64450
rect 28300 64390 28330 64460
rect 28190 64350 28330 64390
rect 30119 63820 30120 65140
rect 31440 63820 31441 65140
rect 30119 63819 31441 63820
rect 26722 63752 26818 63768
rect 26722 63482 26818 63498
rect 25129 63430 26451 63431
rect 23200 62860 23340 62890
rect 23200 62800 23230 62860
rect 21812 62790 23230 62800
rect 23310 62790 23340 62860
rect 21812 62750 23340 62790
rect 21812 62740 23230 62750
rect 21812 62058 21828 62740
rect 23200 62680 23230 62740
rect 23310 62680 23340 62750
rect 23200 62640 23340 62680
rect 25129 62110 25130 63430
rect 26450 62110 26451 63430
rect 25129 62109 26451 62110
rect 21732 62042 21828 62058
rect 21732 61772 21828 61788
rect 20139 61720 21461 61721
rect 18210 61150 18350 61180
rect 18210 61090 18240 61150
rect 16822 61080 18240 61090
rect 18320 61080 18350 61150
rect 16822 61040 18350 61080
rect 16822 61030 18240 61040
rect 16822 60348 16838 61030
rect 18210 60970 18240 61030
rect 18320 60970 18350 61040
rect 18210 60930 18350 60970
rect 20139 60400 20140 61720
rect 21460 60400 21461 61720
rect 20139 60399 21461 60400
rect 16742 60332 16838 60348
rect 16742 60062 16838 60078
rect 15149 60010 16471 60011
rect 13220 59440 13360 59470
rect 13220 59380 13250 59440
rect 11832 59370 13250 59380
rect 13330 59370 13360 59440
rect 11832 59330 13360 59370
rect 11832 59320 13250 59330
rect 11832 58638 11848 59320
rect 13220 59260 13250 59320
rect 13330 59260 13360 59330
rect 13220 59220 13360 59260
rect 15149 58690 15150 60010
rect 16470 58690 16471 60010
rect 15149 58689 16471 58690
rect 11752 58622 11848 58638
rect 11752 58352 11848 58368
rect 10159 58300 11481 58301
rect 8230 57730 8370 57760
rect 8230 57670 8260 57730
rect 6842 57660 8260 57670
rect 8340 57660 8370 57730
rect 6842 57620 8370 57660
rect 6842 57610 8260 57620
rect 6842 56928 6858 57610
rect 8230 57550 8260 57610
rect 8340 57550 8370 57620
rect 8230 57510 8370 57550
rect 10159 56980 10160 58300
rect 11480 56980 11481 58300
rect 10159 56979 11481 56980
rect 6762 56912 6858 56928
rect 6762 56642 6858 56658
rect 5169 56590 6491 56591
rect 3240 56020 3380 56050
rect 3240 55960 3270 56020
rect 1852 55950 3270 55960
rect 3350 55950 3380 56020
rect 1852 55910 3380 55950
rect 1852 55900 3270 55910
rect 1852 55218 1868 55900
rect 3240 55840 3270 55900
rect 3350 55840 3380 55910
rect 3240 55800 3380 55840
rect 5169 55270 5170 56590
rect 6490 55270 6491 56590
rect 5169 55269 6491 55270
rect 1772 55202 1868 55218
rect 1772 54932 1868 54948
rect 179 54880 1501 54881
rect 179 53560 180 54880
rect 1500 53560 1501 54880
rect 179 53559 1501 53560
rect 180 53171 240 53559
rect 1772 53508 1788 54932
rect 1852 54250 1868 54932
rect 5170 54881 5230 55269
rect 6762 55218 6778 56642
rect 6842 55960 6858 56642
rect 10160 56591 10220 56979
rect 11752 56928 11768 58352
rect 11832 57670 11848 58352
rect 15150 58301 15210 58689
rect 16742 58638 16758 60062
rect 16822 59380 16838 60062
rect 20140 60011 20200 60399
rect 21732 60348 21748 61772
rect 21812 61090 21828 61772
rect 25130 61721 25190 62109
rect 26722 62058 26738 63482
rect 26802 62800 26818 63482
rect 30120 63431 30180 63819
rect 31712 63768 31728 65192
rect 31792 64510 31808 65192
rect 35110 65141 35170 65529
rect 36702 65478 36718 66902
rect 36782 66220 36798 66902
rect 40100 66851 40160 67110
rect 41692 66902 41788 66918
rect 40099 66850 41421 66851
rect 38170 66280 38310 66310
rect 38170 66220 38200 66280
rect 36782 66210 38200 66220
rect 38280 66210 38310 66280
rect 36782 66170 38310 66210
rect 36782 66160 38200 66170
rect 36782 65478 36798 66160
rect 38170 66100 38200 66160
rect 38280 66100 38310 66170
rect 38170 66060 38310 66100
rect 40099 65530 40100 66850
rect 41420 65530 41421 66850
rect 40099 65529 41421 65530
rect 36702 65462 36798 65478
rect 36702 65192 36798 65208
rect 35109 65140 36431 65141
rect 33180 64570 33320 64600
rect 33180 64510 33210 64570
rect 31792 64500 33210 64510
rect 33290 64500 33320 64570
rect 31792 64460 33320 64500
rect 31792 64450 33210 64460
rect 31792 63768 31808 64450
rect 33180 64390 33210 64450
rect 33290 64390 33320 64460
rect 34010 64450 34700 64510
rect 33180 64350 33320 64390
rect 35109 63820 35110 65140
rect 36430 63820 36431 65140
rect 35109 63819 36431 63820
rect 31712 63752 31808 63768
rect 31712 63482 31808 63498
rect 30119 63430 31441 63431
rect 28190 62860 28330 62890
rect 28190 62800 28220 62860
rect 26802 62790 28220 62800
rect 28300 62790 28330 62860
rect 26802 62750 28330 62790
rect 26802 62740 28220 62750
rect 26802 62058 26818 62740
rect 28190 62680 28220 62740
rect 28300 62680 28330 62750
rect 28190 62640 28330 62680
rect 30119 62110 30120 63430
rect 31440 62110 31441 63430
rect 30119 62109 31441 62110
rect 26722 62042 26818 62058
rect 26722 61772 26818 61788
rect 25129 61720 26451 61721
rect 23200 61150 23340 61180
rect 23200 61090 23230 61150
rect 21812 61080 23230 61090
rect 23310 61080 23340 61150
rect 21812 61040 23340 61080
rect 21812 61030 23230 61040
rect 21812 60348 21828 61030
rect 23200 60970 23230 61030
rect 23310 60970 23340 61040
rect 23200 60930 23340 60970
rect 25129 60400 25130 61720
rect 26450 60400 26451 61720
rect 25129 60399 26451 60400
rect 21732 60332 21828 60348
rect 21732 60062 21828 60078
rect 20139 60010 21461 60011
rect 18210 59440 18350 59470
rect 18210 59380 18240 59440
rect 16822 59370 18240 59380
rect 18320 59370 18350 59440
rect 16822 59330 18350 59370
rect 16822 59320 18240 59330
rect 16822 58638 16838 59320
rect 18210 59260 18240 59320
rect 18320 59260 18350 59330
rect 18210 59220 18350 59260
rect 20139 58690 20140 60010
rect 21460 58690 21461 60010
rect 20139 58689 21461 58690
rect 16742 58622 16838 58638
rect 16742 58352 16838 58368
rect 15149 58300 16471 58301
rect 13220 57730 13360 57760
rect 13220 57670 13250 57730
rect 11832 57660 13250 57670
rect 13330 57660 13360 57730
rect 11832 57620 13360 57660
rect 11832 57610 13250 57620
rect 11832 56928 11848 57610
rect 13220 57550 13250 57610
rect 13330 57550 13360 57620
rect 13220 57510 13360 57550
rect 15149 56980 15150 58300
rect 16470 56980 16471 58300
rect 15149 56979 16471 56980
rect 11752 56912 11848 56928
rect 11752 56642 11848 56658
rect 10159 56590 11481 56591
rect 8230 56020 8370 56050
rect 8230 55960 8260 56020
rect 6842 55950 8260 55960
rect 8340 55950 8370 56020
rect 6842 55910 8370 55950
rect 6842 55900 8260 55910
rect 6842 55218 6858 55900
rect 8230 55840 8260 55900
rect 8340 55840 8370 55910
rect 8230 55800 8370 55840
rect 10159 55270 10160 56590
rect 11480 55270 11481 56590
rect 10159 55269 11481 55270
rect 6762 55202 6858 55218
rect 6762 54932 6858 54948
rect 5169 54880 6491 54881
rect 3240 54310 3380 54340
rect 3240 54250 3270 54310
rect 1852 54240 3270 54250
rect 3350 54240 3380 54310
rect 1852 54200 3380 54240
rect 1852 54190 3270 54200
rect 1852 53508 1868 54190
rect 3240 54130 3270 54190
rect 3350 54130 3380 54200
rect 3240 54090 3380 54130
rect 5169 53560 5170 54880
rect 6490 53560 6491 54880
rect 5169 53559 6491 53560
rect 1772 53492 1868 53508
rect 1772 53222 1868 53238
rect 179 53170 1501 53171
rect 179 51850 180 53170
rect 1500 51850 1501 53170
rect 179 51849 1501 51850
rect 180 51461 240 51849
rect 1772 51798 1788 53222
rect 1852 52540 1868 53222
rect 5170 53171 5230 53559
rect 6762 53508 6778 54932
rect 6842 54250 6858 54932
rect 10160 54881 10220 55269
rect 11752 55218 11768 56642
rect 11832 55960 11848 56642
rect 15150 56591 15210 56979
rect 16742 56928 16758 58352
rect 16822 57670 16838 58352
rect 20140 58301 20200 58689
rect 21732 58638 21748 60062
rect 21812 59380 21828 60062
rect 25130 60011 25190 60399
rect 26722 60348 26738 61772
rect 26802 61090 26818 61772
rect 30120 61721 30180 62109
rect 31712 62058 31728 63482
rect 31792 62800 31808 63482
rect 35110 63431 35170 63819
rect 36702 63768 36718 65192
rect 36782 64510 36798 65192
rect 40100 65141 40160 65529
rect 41692 65478 41708 66902
rect 41772 66220 41788 66902
rect 45090 66851 45150 67110
rect 46682 66902 46778 66918
rect 45089 66850 46411 66851
rect 43160 66280 43300 66310
rect 43160 66220 43190 66280
rect 41772 66210 43190 66220
rect 43270 66210 43300 66280
rect 41772 66170 43300 66210
rect 41772 66160 43190 66170
rect 41772 65478 41788 66160
rect 43160 66100 43190 66160
rect 43270 66100 43300 66170
rect 43160 66060 43300 66100
rect 45089 65530 45090 66850
rect 46410 65530 46411 66850
rect 45089 65529 46411 65530
rect 41692 65462 41788 65478
rect 41692 65192 41788 65208
rect 40099 65140 41421 65141
rect 38170 64570 38310 64600
rect 38170 64510 38200 64570
rect 36782 64500 38200 64510
rect 38280 64500 38310 64570
rect 36782 64460 38310 64500
rect 36782 64450 38200 64460
rect 36782 63768 36798 64450
rect 38170 64390 38200 64450
rect 38280 64390 38310 64460
rect 38170 64350 38310 64390
rect 40099 63820 40100 65140
rect 41420 63820 41421 65140
rect 40099 63819 41421 63820
rect 36702 63752 36798 63768
rect 36702 63482 36798 63498
rect 35109 63430 36431 63431
rect 33180 62860 33320 62890
rect 33180 62800 33210 62860
rect 31792 62790 33210 62800
rect 33290 62790 33320 62860
rect 31792 62750 33320 62790
rect 31792 62740 33210 62750
rect 31792 62058 31808 62740
rect 33180 62680 33210 62740
rect 33290 62680 33320 62750
rect 34010 62740 34700 62800
rect 33180 62640 33320 62680
rect 35109 62110 35110 63430
rect 36430 62110 36431 63430
rect 35109 62109 36431 62110
rect 31712 62042 31808 62058
rect 31712 61772 31808 61788
rect 30119 61720 31441 61721
rect 28190 61150 28330 61180
rect 28190 61090 28220 61150
rect 26802 61080 28220 61090
rect 28300 61080 28330 61150
rect 26802 61040 28330 61080
rect 26802 61030 28220 61040
rect 26802 60348 26818 61030
rect 28190 60970 28220 61030
rect 28300 60970 28330 61040
rect 28190 60930 28330 60970
rect 30119 60400 30120 61720
rect 31440 60400 31441 61720
rect 30119 60399 31441 60400
rect 26722 60332 26818 60348
rect 26722 60062 26818 60078
rect 25129 60010 26451 60011
rect 23200 59440 23340 59470
rect 23200 59380 23230 59440
rect 21812 59370 23230 59380
rect 23310 59370 23340 59440
rect 21812 59330 23340 59370
rect 21812 59320 23230 59330
rect 21812 58638 21828 59320
rect 23200 59260 23230 59320
rect 23310 59260 23340 59330
rect 23200 59220 23340 59260
rect 25129 58690 25130 60010
rect 26450 58690 26451 60010
rect 25129 58689 26451 58690
rect 21732 58622 21828 58638
rect 21732 58352 21828 58368
rect 20139 58300 21461 58301
rect 18210 57730 18350 57760
rect 18210 57670 18240 57730
rect 16822 57660 18240 57670
rect 18320 57660 18350 57730
rect 16822 57620 18350 57660
rect 16822 57610 18240 57620
rect 16822 56928 16838 57610
rect 18210 57550 18240 57610
rect 18320 57550 18350 57620
rect 18210 57510 18350 57550
rect 20139 56980 20140 58300
rect 21460 56980 21461 58300
rect 20139 56979 21461 56980
rect 16742 56912 16838 56928
rect 16742 56642 16838 56658
rect 15149 56590 16471 56591
rect 13220 56020 13360 56050
rect 13220 55960 13250 56020
rect 11832 55950 13250 55960
rect 13330 55950 13360 56020
rect 11832 55910 13360 55950
rect 11832 55900 13250 55910
rect 11832 55218 11848 55900
rect 13220 55840 13250 55900
rect 13330 55840 13360 55910
rect 13220 55800 13360 55840
rect 15149 55270 15150 56590
rect 16470 55270 16471 56590
rect 15149 55269 16471 55270
rect 11752 55202 11848 55218
rect 11752 54932 11848 54948
rect 10159 54880 11481 54881
rect 8230 54310 8370 54340
rect 8230 54250 8260 54310
rect 6842 54240 8260 54250
rect 8340 54240 8370 54310
rect 6842 54200 8370 54240
rect 6842 54190 8260 54200
rect 6842 53508 6858 54190
rect 8230 54130 8260 54190
rect 8340 54130 8370 54200
rect 8230 54090 8370 54130
rect 10159 53560 10160 54880
rect 11480 53560 11481 54880
rect 10159 53559 11481 53560
rect 6762 53492 6858 53508
rect 6762 53222 6858 53238
rect 5169 53170 6491 53171
rect 3240 52600 3380 52630
rect 3240 52540 3270 52600
rect 1852 52530 3270 52540
rect 3350 52530 3380 52600
rect 1852 52490 3380 52530
rect 1852 52480 3270 52490
rect 1852 51798 1868 52480
rect 3240 52420 3270 52480
rect 3350 52420 3380 52490
rect 3240 52380 3380 52420
rect 5169 51850 5170 53170
rect 6490 51850 6491 53170
rect 5169 51849 6491 51850
rect 1772 51782 1868 51798
rect 1772 51512 1868 51528
rect 179 51460 1501 51461
rect 179 50140 180 51460
rect 1500 50140 1501 51460
rect 179 50139 1501 50140
rect 180 49751 240 50139
rect 1772 50088 1788 51512
rect 1852 50830 1868 51512
rect 5170 51461 5230 51849
rect 6762 51798 6778 53222
rect 6842 52540 6858 53222
rect 10160 53171 10220 53559
rect 11752 53508 11768 54932
rect 11832 54250 11848 54932
rect 15150 54881 15210 55269
rect 16742 55218 16758 56642
rect 16822 55960 16838 56642
rect 20140 56591 20200 56979
rect 21732 56928 21748 58352
rect 21812 57670 21828 58352
rect 25130 58301 25190 58689
rect 26722 58638 26738 60062
rect 26802 59380 26818 60062
rect 30120 60011 30180 60399
rect 31712 60348 31728 61772
rect 31792 61090 31808 61772
rect 35110 61721 35170 62109
rect 36702 62058 36718 63482
rect 36782 62800 36798 63482
rect 40100 63431 40160 63819
rect 41692 63768 41708 65192
rect 41772 64510 41788 65192
rect 45090 65141 45150 65529
rect 46682 65478 46698 66902
rect 46762 66220 46778 66902
rect 50080 66851 50140 67110
rect 51672 66902 51768 66918
rect 50079 66850 51401 66851
rect 48150 66280 48290 66310
rect 48150 66220 48180 66280
rect 46762 66210 48180 66220
rect 48260 66210 48290 66280
rect 46762 66170 48290 66210
rect 46762 66160 48180 66170
rect 46762 65478 46778 66160
rect 48150 66100 48180 66160
rect 48260 66100 48290 66170
rect 48980 66160 49670 66220
rect 48150 66060 48290 66100
rect 50079 65530 50080 66850
rect 51400 65530 51401 66850
rect 50079 65529 51401 65530
rect 46682 65462 46778 65478
rect 46682 65192 46778 65208
rect 45089 65140 46411 65141
rect 43160 64570 43300 64600
rect 43160 64510 43190 64570
rect 41772 64500 43190 64510
rect 43270 64500 43300 64570
rect 41772 64460 43300 64500
rect 41772 64450 43190 64460
rect 41772 63768 41788 64450
rect 43160 64390 43190 64450
rect 43270 64390 43300 64460
rect 43160 64350 43300 64390
rect 45089 63820 45090 65140
rect 46410 63820 46411 65140
rect 45089 63819 46411 63820
rect 41692 63752 41788 63768
rect 41692 63482 41788 63498
rect 40099 63430 41421 63431
rect 38170 62860 38310 62890
rect 38170 62800 38200 62860
rect 36782 62790 38200 62800
rect 38280 62790 38310 62860
rect 36782 62750 38310 62790
rect 36782 62740 38200 62750
rect 36782 62058 36798 62740
rect 38170 62680 38200 62740
rect 38280 62680 38310 62750
rect 38170 62640 38310 62680
rect 40099 62110 40100 63430
rect 41420 62110 41421 63430
rect 40099 62109 41421 62110
rect 36702 62042 36798 62058
rect 36702 61772 36798 61788
rect 35109 61720 36431 61721
rect 33180 61150 33320 61180
rect 33180 61090 33210 61150
rect 31792 61080 33210 61090
rect 33290 61080 33320 61150
rect 31792 61040 33320 61080
rect 31792 61030 33210 61040
rect 31792 60348 31808 61030
rect 33180 60970 33210 61030
rect 33290 60970 33320 61040
rect 34010 61030 34700 61090
rect 33180 60930 33320 60970
rect 35109 60400 35110 61720
rect 36430 60400 36431 61720
rect 35109 60399 36431 60400
rect 31712 60332 31808 60348
rect 31712 60062 31808 60078
rect 30119 60010 31441 60011
rect 28190 59440 28330 59470
rect 28190 59380 28220 59440
rect 26802 59370 28220 59380
rect 28300 59370 28330 59440
rect 26802 59330 28330 59370
rect 26802 59320 28220 59330
rect 26802 58638 26818 59320
rect 28190 59260 28220 59320
rect 28300 59260 28330 59330
rect 28190 59220 28330 59260
rect 30119 58690 30120 60010
rect 31440 58690 31441 60010
rect 30119 58689 31441 58690
rect 26722 58622 26818 58638
rect 26722 58352 26818 58368
rect 25129 58300 26451 58301
rect 23200 57730 23340 57760
rect 23200 57670 23230 57730
rect 21812 57660 23230 57670
rect 23310 57660 23340 57730
rect 21812 57620 23340 57660
rect 21812 57610 23230 57620
rect 21812 56928 21828 57610
rect 23200 57550 23230 57610
rect 23310 57550 23340 57620
rect 23200 57510 23340 57550
rect 25129 56980 25130 58300
rect 26450 56980 26451 58300
rect 25129 56979 26451 56980
rect 21732 56912 21828 56928
rect 21732 56642 21828 56658
rect 20139 56590 21461 56591
rect 18210 56020 18350 56050
rect 18210 55960 18240 56020
rect 16822 55950 18240 55960
rect 18320 55950 18350 56020
rect 16822 55910 18350 55950
rect 16822 55900 18240 55910
rect 16822 55218 16838 55900
rect 18210 55840 18240 55900
rect 18320 55840 18350 55910
rect 18210 55800 18350 55840
rect 20139 55270 20140 56590
rect 21460 55270 21461 56590
rect 20139 55269 21461 55270
rect 16742 55202 16838 55218
rect 16742 54932 16838 54948
rect 15149 54880 16471 54881
rect 13220 54310 13360 54340
rect 13220 54250 13250 54310
rect 11832 54240 13250 54250
rect 13330 54240 13360 54310
rect 11832 54200 13360 54240
rect 11832 54190 13250 54200
rect 11832 53508 11848 54190
rect 13220 54130 13250 54190
rect 13330 54130 13360 54200
rect 13220 54090 13360 54130
rect 15149 53560 15150 54880
rect 16470 53560 16471 54880
rect 15149 53559 16471 53560
rect 11752 53492 11848 53508
rect 11752 53222 11848 53238
rect 10159 53170 11481 53171
rect 8230 52600 8370 52630
rect 8230 52540 8260 52600
rect 6842 52530 8260 52540
rect 8340 52530 8370 52600
rect 6842 52490 8370 52530
rect 6842 52480 8260 52490
rect 6842 51798 6858 52480
rect 8230 52420 8260 52480
rect 8340 52420 8370 52490
rect 8230 52380 8370 52420
rect 10159 51850 10160 53170
rect 11480 51850 11481 53170
rect 10159 51849 11481 51850
rect 6762 51782 6858 51798
rect 6762 51512 6858 51528
rect 5169 51460 6491 51461
rect 3240 50890 3380 50920
rect 3240 50830 3270 50890
rect 1852 50820 3270 50830
rect 3350 50820 3380 50890
rect 1852 50780 3380 50820
rect 1852 50770 3270 50780
rect 1852 50088 1868 50770
rect 3240 50710 3270 50770
rect 3350 50710 3380 50780
rect 3240 50670 3380 50710
rect 5169 50140 5170 51460
rect 6490 50140 6491 51460
rect 5169 50139 6491 50140
rect 1772 50072 1868 50088
rect 1772 49802 1868 49818
rect 179 49750 1501 49751
rect 179 48430 180 49750
rect 1500 48430 1501 49750
rect 179 48429 1501 48430
rect 180 48041 240 48429
rect 1772 48378 1788 49802
rect 1852 49120 1868 49802
rect 5170 49751 5230 50139
rect 6762 50088 6778 51512
rect 6842 50830 6858 51512
rect 10160 51461 10220 51849
rect 11752 51798 11768 53222
rect 11832 52540 11848 53222
rect 15150 53171 15210 53559
rect 16742 53508 16758 54932
rect 16822 54250 16838 54932
rect 20140 54881 20200 55269
rect 21732 55218 21748 56642
rect 21812 55960 21828 56642
rect 25130 56591 25190 56979
rect 26722 56928 26738 58352
rect 26802 57670 26818 58352
rect 30120 58301 30180 58689
rect 31712 58638 31728 60062
rect 31792 59380 31808 60062
rect 35110 60011 35170 60399
rect 36702 60348 36718 61772
rect 36782 61090 36798 61772
rect 40100 61721 40160 62109
rect 41692 62058 41708 63482
rect 41772 62800 41788 63482
rect 45090 63431 45150 63819
rect 46682 63768 46698 65192
rect 46762 64510 46778 65192
rect 50080 65141 50140 65529
rect 51672 65478 51688 66902
rect 51752 66220 51768 66902
rect 55070 66851 55130 67110
rect 56662 66902 56758 66918
rect 55069 66850 56391 66851
rect 53140 66280 53280 66310
rect 53140 66220 53170 66280
rect 51752 66210 53170 66220
rect 53250 66210 53280 66280
rect 51752 66170 53280 66210
rect 51752 66160 53170 66170
rect 51752 65478 51768 66160
rect 53140 66100 53170 66160
rect 53250 66100 53280 66170
rect 53140 66060 53280 66100
rect 55069 65530 55070 66850
rect 56390 65530 56391 66850
rect 55069 65529 56391 65530
rect 51672 65462 51768 65478
rect 51672 65192 51768 65208
rect 50079 65140 51401 65141
rect 48150 64570 48290 64600
rect 48150 64510 48180 64570
rect 46762 64500 48180 64510
rect 48260 64500 48290 64570
rect 46762 64460 48290 64500
rect 46762 64450 48180 64460
rect 46762 63768 46778 64450
rect 48150 64390 48180 64450
rect 48260 64390 48290 64460
rect 48980 64450 49670 64510
rect 48150 64350 48290 64390
rect 50079 63820 50080 65140
rect 51400 63820 51401 65140
rect 50079 63819 51401 63820
rect 46682 63752 46778 63768
rect 46682 63482 46778 63498
rect 45089 63430 46411 63431
rect 43160 62860 43300 62890
rect 43160 62800 43190 62860
rect 41772 62790 43190 62800
rect 43270 62790 43300 62860
rect 41772 62750 43300 62790
rect 41772 62740 43190 62750
rect 41772 62058 41788 62740
rect 43160 62680 43190 62740
rect 43270 62680 43300 62750
rect 43160 62640 43300 62680
rect 45089 62110 45090 63430
rect 46410 62110 46411 63430
rect 45089 62109 46411 62110
rect 41692 62042 41788 62058
rect 41692 61772 41788 61788
rect 40099 61720 41421 61721
rect 38170 61150 38310 61180
rect 38170 61090 38200 61150
rect 36782 61080 38200 61090
rect 38280 61080 38310 61150
rect 36782 61040 38310 61080
rect 36782 61030 38200 61040
rect 36782 60348 36798 61030
rect 38170 60970 38200 61030
rect 38280 60970 38310 61040
rect 38170 60930 38310 60970
rect 40099 60400 40100 61720
rect 41420 60400 41421 61720
rect 40099 60399 41421 60400
rect 36702 60332 36798 60348
rect 36702 60062 36798 60078
rect 35109 60010 36431 60011
rect 33180 59440 33320 59470
rect 33180 59380 33210 59440
rect 31792 59370 33210 59380
rect 33290 59370 33320 59440
rect 31792 59330 33320 59370
rect 31792 59320 33210 59330
rect 31792 58638 31808 59320
rect 33180 59260 33210 59320
rect 33290 59260 33320 59330
rect 34010 59320 34700 59380
rect 33180 59220 33320 59260
rect 35109 58690 35110 60010
rect 36430 58690 36431 60010
rect 35109 58689 36431 58690
rect 31712 58622 31808 58638
rect 31712 58352 31808 58368
rect 30119 58300 31441 58301
rect 28190 57730 28330 57760
rect 28190 57670 28220 57730
rect 26802 57660 28220 57670
rect 28300 57660 28330 57730
rect 26802 57620 28330 57660
rect 26802 57610 28220 57620
rect 26802 56928 26818 57610
rect 28190 57550 28220 57610
rect 28300 57550 28330 57620
rect 28190 57510 28330 57550
rect 30119 56980 30120 58300
rect 31440 56980 31441 58300
rect 30119 56979 31441 56980
rect 26722 56912 26818 56928
rect 26722 56642 26818 56658
rect 25129 56590 26451 56591
rect 23200 56020 23340 56050
rect 23200 55960 23230 56020
rect 21812 55950 23230 55960
rect 23310 55950 23340 56020
rect 21812 55910 23340 55950
rect 21812 55900 23230 55910
rect 21812 55218 21828 55900
rect 23200 55840 23230 55900
rect 23310 55840 23340 55910
rect 23200 55800 23340 55840
rect 25129 55270 25130 56590
rect 26450 55270 26451 56590
rect 25129 55269 26451 55270
rect 21732 55202 21828 55218
rect 21732 54932 21828 54948
rect 20139 54880 21461 54881
rect 18210 54310 18350 54340
rect 18210 54250 18240 54310
rect 16822 54240 18240 54250
rect 18320 54240 18350 54310
rect 16822 54200 18350 54240
rect 16822 54190 18240 54200
rect 16822 53508 16838 54190
rect 18210 54130 18240 54190
rect 18320 54130 18350 54200
rect 18210 54090 18350 54130
rect 20139 53560 20140 54880
rect 21460 53560 21461 54880
rect 20139 53559 21461 53560
rect 16742 53492 16838 53508
rect 16742 53222 16838 53238
rect 15149 53170 16471 53171
rect 13220 52600 13360 52630
rect 13220 52540 13250 52600
rect 11832 52530 13250 52540
rect 13330 52530 13360 52600
rect 11832 52490 13360 52530
rect 11832 52480 13250 52490
rect 11832 51798 11848 52480
rect 13220 52420 13250 52480
rect 13330 52420 13360 52490
rect 13220 52380 13360 52420
rect 15149 51850 15150 53170
rect 16470 51850 16471 53170
rect 15149 51849 16471 51850
rect 11752 51782 11848 51798
rect 11752 51512 11848 51528
rect 10159 51460 11481 51461
rect 8230 50890 8370 50920
rect 8230 50830 8260 50890
rect 6842 50820 8260 50830
rect 8340 50820 8370 50890
rect 6842 50780 8370 50820
rect 6842 50770 8260 50780
rect 6842 50088 6858 50770
rect 8230 50710 8260 50770
rect 8340 50710 8370 50780
rect 8230 50670 8370 50710
rect 10159 50140 10160 51460
rect 11480 50140 11481 51460
rect 10159 50139 11481 50140
rect 6762 50072 6858 50088
rect 6762 49802 6858 49818
rect 5169 49750 6491 49751
rect 3240 49180 3380 49210
rect 3240 49120 3270 49180
rect 1852 49110 3270 49120
rect 3350 49110 3380 49180
rect 1852 49070 3380 49110
rect 1852 49060 3270 49070
rect 1852 48378 1868 49060
rect 3240 49000 3270 49060
rect 3350 49000 3380 49070
rect 3240 48960 3380 49000
rect 5169 48430 5170 49750
rect 6490 48430 6491 49750
rect 5169 48429 6491 48430
rect 1772 48362 1868 48378
rect 1772 48092 1868 48108
rect 179 48040 1501 48041
rect 179 46720 180 48040
rect 1500 46720 1501 48040
rect 179 46719 1501 46720
rect 180 46331 240 46719
rect 1772 46668 1788 48092
rect 1852 47410 1868 48092
rect 5170 48041 5230 48429
rect 6762 48378 6778 49802
rect 6842 49120 6858 49802
rect 10160 49751 10220 50139
rect 11752 50088 11768 51512
rect 11832 50830 11848 51512
rect 15150 51461 15210 51849
rect 16742 51798 16758 53222
rect 16822 52540 16838 53222
rect 20140 53171 20200 53559
rect 21732 53508 21748 54932
rect 21812 54250 21828 54932
rect 25130 54881 25190 55269
rect 26722 55218 26738 56642
rect 26802 55960 26818 56642
rect 30120 56591 30180 56979
rect 31712 56928 31728 58352
rect 31792 57670 31808 58352
rect 35110 58301 35170 58689
rect 36702 58638 36718 60062
rect 36782 59380 36798 60062
rect 40100 60011 40160 60399
rect 41692 60348 41708 61772
rect 41772 61090 41788 61772
rect 45090 61721 45150 62109
rect 46682 62058 46698 63482
rect 46762 62800 46778 63482
rect 50080 63431 50140 63819
rect 51672 63768 51688 65192
rect 51752 64510 51768 65192
rect 55070 65141 55130 65529
rect 56662 65478 56678 66902
rect 56742 66220 56758 66902
rect 60060 66851 60120 67110
rect 61652 66902 61748 66918
rect 60059 66850 61381 66851
rect 58130 66280 58270 66310
rect 58130 66220 58160 66280
rect 56742 66210 58160 66220
rect 58240 66210 58270 66280
rect 56742 66170 58270 66210
rect 56742 66160 58160 66170
rect 56742 65478 56758 66160
rect 58130 66100 58160 66160
rect 58240 66100 58270 66170
rect 58130 66060 58270 66100
rect 60059 65530 60060 66850
rect 61380 65530 61381 66850
rect 60059 65529 61381 65530
rect 56662 65462 56758 65478
rect 56662 65192 56758 65208
rect 55069 65140 56391 65141
rect 53140 64570 53280 64600
rect 53140 64510 53170 64570
rect 51752 64500 53170 64510
rect 53250 64500 53280 64570
rect 51752 64460 53280 64500
rect 51752 64450 53170 64460
rect 51752 63768 51768 64450
rect 53140 64390 53170 64450
rect 53250 64390 53280 64460
rect 53140 64350 53280 64390
rect 55069 63820 55070 65140
rect 56390 63820 56391 65140
rect 55069 63819 56391 63820
rect 51672 63752 51768 63768
rect 51672 63482 51768 63498
rect 50079 63430 51401 63431
rect 48150 62860 48290 62890
rect 48150 62800 48180 62860
rect 46762 62790 48180 62800
rect 48260 62790 48290 62860
rect 46762 62750 48290 62790
rect 46762 62740 48180 62750
rect 46762 62058 46778 62740
rect 48150 62680 48180 62740
rect 48260 62680 48290 62750
rect 48980 62740 49670 62800
rect 48150 62640 48290 62680
rect 50079 62110 50080 63430
rect 51400 62110 51401 63430
rect 50079 62109 51401 62110
rect 46682 62042 46778 62058
rect 46682 61772 46778 61788
rect 45089 61720 46411 61721
rect 43160 61150 43300 61180
rect 43160 61090 43190 61150
rect 41772 61080 43190 61090
rect 43270 61080 43300 61150
rect 41772 61040 43300 61080
rect 41772 61030 43190 61040
rect 41772 60348 41788 61030
rect 43160 60970 43190 61030
rect 43270 60970 43300 61040
rect 43160 60930 43300 60970
rect 45089 60400 45090 61720
rect 46410 60400 46411 61720
rect 45089 60399 46411 60400
rect 41692 60332 41788 60348
rect 41692 60062 41788 60078
rect 40099 60010 41421 60011
rect 38170 59440 38310 59470
rect 38170 59380 38200 59440
rect 36782 59370 38200 59380
rect 38280 59370 38310 59440
rect 36782 59330 38310 59370
rect 36782 59320 38200 59330
rect 36782 58638 36798 59320
rect 38170 59260 38200 59320
rect 38280 59260 38310 59330
rect 38170 59220 38310 59260
rect 40099 58690 40100 60010
rect 41420 58690 41421 60010
rect 40099 58689 41421 58690
rect 36702 58622 36798 58638
rect 36702 58352 36798 58368
rect 35109 58300 36431 58301
rect 33180 57730 33320 57760
rect 33180 57670 33210 57730
rect 31792 57660 33210 57670
rect 33290 57660 33320 57730
rect 31792 57620 33320 57660
rect 31792 57610 33210 57620
rect 31792 56928 31808 57610
rect 33180 57550 33210 57610
rect 33290 57550 33320 57620
rect 34010 57610 34700 57670
rect 33180 57510 33320 57550
rect 35109 56980 35110 58300
rect 36430 56980 36431 58300
rect 35109 56979 36431 56980
rect 31712 56912 31808 56928
rect 31712 56642 31808 56658
rect 30119 56590 31441 56591
rect 28190 56020 28330 56050
rect 28190 55960 28220 56020
rect 26802 55950 28220 55960
rect 28300 55950 28330 56020
rect 26802 55910 28330 55950
rect 26802 55900 28220 55910
rect 26802 55218 26818 55900
rect 28190 55840 28220 55900
rect 28300 55840 28330 55910
rect 28190 55800 28330 55840
rect 30119 55270 30120 56590
rect 31440 55270 31441 56590
rect 30119 55269 31441 55270
rect 26722 55202 26818 55218
rect 26722 54932 26818 54948
rect 25129 54880 26451 54881
rect 23200 54310 23340 54340
rect 23200 54250 23230 54310
rect 21812 54240 23230 54250
rect 23310 54240 23340 54310
rect 21812 54200 23340 54240
rect 21812 54190 23230 54200
rect 21812 53508 21828 54190
rect 23200 54130 23230 54190
rect 23310 54130 23340 54200
rect 23200 54090 23340 54130
rect 25129 53560 25130 54880
rect 26450 53560 26451 54880
rect 25129 53559 26451 53560
rect 21732 53492 21828 53508
rect 21732 53222 21828 53238
rect 20139 53170 21461 53171
rect 18210 52600 18350 52630
rect 18210 52540 18240 52600
rect 16822 52530 18240 52540
rect 18320 52530 18350 52600
rect 16822 52490 18350 52530
rect 16822 52480 18240 52490
rect 16822 51798 16838 52480
rect 18210 52420 18240 52480
rect 18320 52420 18350 52490
rect 18210 52380 18350 52420
rect 20139 51850 20140 53170
rect 21460 51850 21461 53170
rect 20139 51849 21461 51850
rect 16742 51782 16838 51798
rect 16742 51512 16838 51528
rect 15149 51460 16471 51461
rect 13220 50890 13360 50920
rect 13220 50830 13250 50890
rect 11832 50820 13250 50830
rect 13330 50820 13360 50890
rect 11832 50780 13360 50820
rect 11832 50770 13250 50780
rect 11832 50088 11848 50770
rect 13220 50710 13250 50770
rect 13330 50710 13360 50780
rect 13220 50670 13360 50710
rect 15149 50140 15150 51460
rect 16470 50140 16471 51460
rect 15149 50139 16471 50140
rect 11752 50072 11848 50088
rect 11752 49802 11848 49818
rect 10159 49750 11481 49751
rect 8230 49180 8370 49210
rect 8230 49120 8260 49180
rect 6842 49110 8260 49120
rect 8340 49110 8370 49180
rect 6842 49070 8370 49110
rect 6842 49060 8260 49070
rect 6842 48378 6858 49060
rect 8230 49000 8260 49060
rect 8340 49000 8370 49070
rect 8230 48960 8370 49000
rect 10159 48430 10160 49750
rect 11480 48430 11481 49750
rect 10159 48429 11481 48430
rect 6762 48362 6858 48378
rect 6762 48092 6858 48108
rect 5169 48040 6491 48041
rect 3240 47470 3380 47500
rect 3240 47410 3270 47470
rect 1852 47400 3270 47410
rect 3350 47400 3380 47470
rect 1852 47360 3380 47400
rect 1852 47350 3270 47360
rect 1852 46668 1868 47350
rect 3240 47290 3270 47350
rect 3350 47290 3380 47360
rect 3240 47250 3380 47290
rect 5169 46720 5170 48040
rect 6490 46720 6491 48040
rect 5169 46719 6491 46720
rect 1772 46652 1868 46668
rect 1772 46382 1868 46398
rect 179 46330 1501 46331
rect 179 45010 180 46330
rect 1500 45010 1501 46330
rect 179 45009 1501 45010
rect 180 44621 240 45009
rect 1772 44958 1788 46382
rect 1852 45700 1868 46382
rect 5170 46331 5230 46719
rect 6762 46668 6778 48092
rect 6842 47410 6858 48092
rect 10160 48041 10220 48429
rect 11752 48378 11768 49802
rect 11832 49120 11848 49802
rect 15150 49751 15210 50139
rect 16742 50088 16758 51512
rect 16822 50830 16838 51512
rect 20140 51461 20200 51849
rect 21732 51798 21748 53222
rect 21812 52540 21828 53222
rect 25130 53171 25190 53559
rect 26722 53508 26738 54932
rect 26802 54250 26818 54932
rect 30120 54881 30180 55269
rect 31712 55218 31728 56642
rect 31792 55960 31808 56642
rect 35110 56591 35170 56979
rect 36702 56928 36718 58352
rect 36782 57670 36798 58352
rect 40100 58301 40160 58689
rect 41692 58638 41708 60062
rect 41772 59380 41788 60062
rect 45090 60011 45150 60399
rect 46682 60348 46698 61772
rect 46762 61090 46778 61772
rect 50080 61721 50140 62109
rect 51672 62058 51688 63482
rect 51752 62800 51768 63482
rect 55070 63431 55130 63819
rect 56662 63768 56678 65192
rect 56742 64510 56758 65192
rect 60060 65141 60120 65529
rect 61652 65478 61668 66902
rect 61732 66220 61748 66902
rect 65050 66851 65110 67110
rect 66642 66902 66738 66918
rect 65049 66850 66371 66851
rect 63120 66280 63260 66310
rect 63120 66220 63150 66280
rect 61732 66210 63150 66220
rect 63230 66210 63260 66280
rect 61732 66170 63260 66210
rect 61732 66160 63150 66170
rect 61732 65478 61748 66160
rect 63120 66100 63150 66160
rect 63230 66100 63260 66170
rect 63120 66060 63260 66100
rect 65049 65530 65050 66850
rect 66370 65530 66371 66850
rect 65049 65529 66371 65530
rect 61652 65462 61748 65478
rect 61652 65192 61748 65208
rect 60059 65140 61381 65141
rect 58130 64570 58270 64600
rect 58130 64510 58160 64570
rect 56742 64500 58160 64510
rect 58240 64500 58270 64570
rect 56742 64460 58270 64500
rect 56742 64450 58160 64460
rect 56742 63768 56758 64450
rect 58130 64390 58160 64450
rect 58240 64390 58270 64460
rect 58130 64350 58270 64390
rect 60059 63820 60060 65140
rect 61380 63820 61381 65140
rect 60059 63819 61381 63820
rect 56662 63752 56758 63768
rect 56662 63482 56758 63498
rect 55069 63430 56391 63431
rect 53140 62860 53280 62890
rect 53140 62800 53170 62860
rect 51752 62790 53170 62800
rect 53250 62790 53280 62860
rect 51752 62750 53280 62790
rect 51752 62740 53170 62750
rect 51752 62058 51768 62740
rect 53140 62680 53170 62740
rect 53250 62680 53280 62750
rect 53140 62640 53280 62680
rect 55069 62110 55070 63430
rect 56390 62110 56391 63430
rect 55069 62109 56391 62110
rect 51672 62042 51768 62058
rect 51672 61772 51768 61788
rect 50079 61720 51401 61721
rect 48150 61150 48290 61180
rect 48150 61090 48180 61150
rect 46762 61080 48180 61090
rect 48260 61080 48290 61150
rect 46762 61040 48290 61080
rect 46762 61030 48180 61040
rect 46762 60348 46778 61030
rect 48150 60970 48180 61030
rect 48260 60970 48290 61040
rect 48980 61030 49670 61090
rect 48150 60930 48290 60970
rect 50079 60400 50080 61720
rect 51400 60400 51401 61720
rect 50079 60399 51401 60400
rect 46682 60332 46778 60348
rect 46682 60062 46778 60078
rect 45089 60010 46411 60011
rect 43160 59440 43300 59470
rect 43160 59380 43190 59440
rect 41772 59370 43190 59380
rect 43270 59370 43300 59440
rect 41772 59330 43300 59370
rect 41772 59320 43190 59330
rect 41772 58638 41788 59320
rect 43160 59260 43190 59320
rect 43270 59260 43300 59330
rect 43160 59220 43300 59260
rect 45089 58690 45090 60010
rect 46410 58690 46411 60010
rect 45089 58689 46411 58690
rect 41692 58622 41788 58638
rect 41692 58352 41788 58368
rect 40099 58300 41421 58301
rect 38170 57730 38310 57760
rect 38170 57670 38200 57730
rect 36782 57660 38200 57670
rect 38280 57660 38310 57730
rect 36782 57620 38310 57660
rect 36782 57610 38200 57620
rect 36782 56928 36798 57610
rect 38170 57550 38200 57610
rect 38280 57550 38310 57620
rect 38170 57510 38310 57550
rect 40099 56980 40100 58300
rect 41420 56980 41421 58300
rect 40099 56979 41421 56980
rect 36702 56912 36798 56928
rect 36702 56642 36798 56658
rect 35109 56590 36431 56591
rect 33180 56020 33320 56050
rect 33180 55960 33210 56020
rect 31792 55950 33210 55960
rect 33290 55950 33320 56020
rect 31792 55910 33320 55950
rect 31792 55900 33210 55910
rect 31792 55218 31808 55900
rect 33180 55840 33210 55900
rect 33290 55840 33320 55910
rect 34010 55900 34700 55960
rect 33180 55800 33320 55840
rect 35109 55270 35110 56590
rect 36430 55270 36431 56590
rect 35109 55269 36431 55270
rect 31712 55202 31808 55218
rect 31712 54932 31808 54948
rect 30119 54880 31441 54881
rect 28190 54310 28330 54340
rect 28190 54250 28220 54310
rect 26802 54240 28220 54250
rect 28300 54240 28330 54310
rect 26802 54200 28330 54240
rect 26802 54190 28220 54200
rect 26802 53508 26818 54190
rect 28190 54130 28220 54190
rect 28300 54130 28330 54200
rect 28190 54090 28330 54130
rect 30119 53560 30120 54880
rect 31440 53560 31441 54880
rect 30119 53559 31441 53560
rect 26722 53492 26818 53508
rect 26722 53222 26818 53238
rect 25129 53170 26451 53171
rect 23200 52600 23340 52630
rect 23200 52540 23230 52600
rect 21812 52530 23230 52540
rect 23310 52530 23340 52600
rect 21812 52490 23340 52530
rect 21812 52480 23230 52490
rect 21812 51798 21828 52480
rect 23200 52420 23230 52480
rect 23310 52420 23340 52490
rect 23200 52380 23340 52420
rect 25129 51850 25130 53170
rect 26450 51850 26451 53170
rect 25129 51849 26451 51850
rect 21732 51782 21828 51798
rect 21732 51512 21828 51528
rect 20139 51460 21461 51461
rect 18210 50890 18350 50920
rect 18210 50830 18240 50890
rect 16822 50820 18240 50830
rect 18320 50820 18350 50890
rect 16822 50780 18350 50820
rect 16822 50770 18240 50780
rect 16822 50088 16838 50770
rect 18210 50710 18240 50770
rect 18320 50710 18350 50780
rect 18210 50670 18350 50710
rect 20139 50140 20140 51460
rect 21460 50140 21461 51460
rect 20139 50139 21461 50140
rect 16742 50072 16838 50088
rect 16742 49802 16838 49818
rect 15149 49750 16471 49751
rect 13220 49180 13360 49210
rect 13220 49120 13250 49180
rect 11832 49110 13250 49120
rect 13330 49110 13360 49180
rect 11832 49070 13360 49110
rect 11832 49060 13250 49070
rect 11832 48378 11848 49060
rect 13220 49000 13250 49060
rect 13330 49000 13360 49070
rect 13220 48960 13360 49000
rect 15149 48430 15150 49750
rect 16470 48430 16471 49750
rect 15149 48429 16471 48430
rect 11752 48362 11848 48378
rect 11752 48092 11848 48108
rect 10159 48040 11481 48041
rect 8230 47470 8370 47500
rect 8230 47410 8260 47470
rect 6842 47400 8260 47410
rect 8340 47400 8370 47470
rect 6842 47360 8370 47400
rect 6842 47350 8260 47360
rect 6842 46668 6858 47350
rect 8230 47290 8260 47350
rect 8340 47290 8370 47360
rect 8230 47250 8370 47290
rect 10159 46720 10160 48040
rect 11480 46720 11481 48040
rect 10159 46719 11481 46720
rect 6762 46652 6858 46668
rect 6762 46382 6858 46398
rect 5169 46330 6491 46331
rect 3240 45760 3380 45790
rect 3240 45700 3270 45760
rect 1852 45690 3270 45700
rect 3350 45690 3380 45760
rect 1852 45650 3380 45690
rect 1852 45640 3270 45650
rect 1852 44958 1868 45640
rect 3240 45580 3270 45640
rect 3350 45580 3380 45650
rect 3240 45540 3380 45580
rect 5169 45010 5170 46330
rect 6490 45010 6491 46330
rect 5169 45009 6491 45010
rect 1772 44942 1868 44958
rect 1772 44672 1868 44688
rect 179 44620 1501 44621
rect 179 43300 180 44620
rect 1500 43300 1501 44620
rect 179 43299 1501 43300
rect 180 42911 240 43299
rect 1772 43248 1788 44672
rect 1852 43990 1868 44672
rect 5170 44621 5230 45009
rect 6762 44958 6778 46382
rect 6842 45700 6858 46382
rect 10160 46331 10220 46719
rect 11752 46668 11768 48092
rect 11832 47410 11848 48092
rect 15150 48041 15210 48429
rect 16742 48378 16758 49802
rect 16822 49120 16838 49802
rect 20140 49751 20200 50139
rect 21732 50088 21748 51512
rect 21812 50830 21828 51512
rect 25130 51461 25190 51849
rect 26722 51798 26738 53222
rect 26802 52540 26818 53222
rect 30120 53171 30180 53559
rect 31712 53508 31728 54932
rect 31792 54250 31808 54932
rect 35110 54881 35170 55269
rect 36702 55218 36718 56642
rect 36782 55960 36798 56642
rect 40100 56591 40160 56979
rect 41692 56928 41708 58352
rect 41772 57670 41788 58352
rect 45090 58301 45150 58689
rect 46682 58638 46698 60062
rect 46762 59380 46778 60062
rect 50080 60011 50140 60399
rect 51672 60348 51688 61772
rect 51752 61090 51768 61772
rect 55070 61721 55130 62109
rect 56662 62058 56678 63482
rect 56742 62800 56758 63482
rect 60060 63431 60120 63819
rect 61652 63768 61668 65192
rect 61732 64510 61748 65192
rect 65050 65141 65110 65529
rect 66642 65478 66658 66902
rect 66722 66220 66738 66902
rect 70040 66851 70100 67110
rect 71632 66902 71728 66918
rect 70039 66850 71361 66851
rect 68110 66280 68250 66310
rect 68110 66220 68140 66280
rect 66722 66210 68140 66220
rect 68220 66210 68250 66280
rect 66722 66170 68250 66210
rect 66722 66160 68140 66170
rect 66722 65478 66738 66160
rect 68110 66100 68140 66160
rect 68220 66100 68250 66170
rect 68110 66060 68250 66100
rect 70039 65530 70040 66850
rect 71360 65530 71361 66850
rect 70039 65529 71361 65530
rect 66642 65462 66738 65478
rect 66642 65192 66738 65208
rect 65049 65140 66371 65141
rect 63120 64570 63260 64600
rect 63120 64510 63150 64570
rect 61732 64500 63150 64510
rect 63230 64500 63260 64570
rect 61732 64460 63260 64500
rect 61732 64450 63150 64460
rect 61732 63768 61748 64450
rect 63120 64390 63150 64450
rect 63230 64390 63260 64460
rect 63120 64350 63260 64390
rect 65049 63820 65050 65140
rect 66370 63820 66371 65140
rect 65049 63819 66371 63820
rect 61652 63752 61748 63768
rect 61652 63482 61748 63498
rect 60059 63430 61381 63431
rect 58130 62860 58270 62890
rect 58130 62800 58160 62860
rect 56742 62790 58160 62800
rect 58240 62790 58270 62860
rect 56742 62750 58270 62790
rect 56742 62740 58160 62750
rect 56742 62058 56758 62740
rect 58130 62680 58160 62740
rect 58240 62680 58270 62750
rect 58130 62640 58270 62680
rect 60059 62110 60060 63430
rect 61380 62110 61381 63430
rect 60059 62109 61381 62110
rect 56662 62042 56758 62058
rect 56662 61772 56758 61788
rect 55069 61720 56391 61721
rect 53140 61150 53280 61180
rect 53140 61090 53170 61150
rect 51752 61080 53170 61090
rect 53250 61080 53280 61150
rect 51752 61040 53280 61080
rect 51752 61030 53170 61040
rect 51752 60348 51768 61030
rect 53140 60970 53170 61030
rect 53250 60970 53280 61040
rect 53140 60930 53280 60970
rect 55069 60400 55070 61720
rect 56390 60400 56391 61720
rect 55069 60399 56391 60400
rect 51672 60332 51768 60348
rect 51672 60062 51768 60078
rect 50079 60010 51401 60011
rect 48150 59440 48290 59470
rect 48150 59380 48180 59440
rect 46762 59370 48180 59380
rect 48260 59370 48290 59440
rect 46762 59330 48290 59370
rect 46762 59320 48180 59330
rect 46762 58638 46778 59320
rect 48150 59260 48180 59320
rect 48260 59260 48290 59330
rect 48980 59320 49670 59380
rect 48150 59220 48290 59260
rect 50079 58690 50080 60010
rect 51400 58690 51401 60010
rect 50079 58689 51401 58690
rect 46682 58622 46778 58638
rect 46682 58352 46778 58368
rect 45089 58300 46411 58301
rect 43160 57730 43300 57760
rect 43160 57670 43190 57730
rect 41772 57660 43190 57670
rect 43270 57660 43300 57730
rect 41772 57620 43300 57660
rect 41772 57610 43190 57620
rect 41772 56928 41788 57610
rect 43160 57550 43190 57610
rect 43270 57550 43300 57620
rect 43160 57510 43300 57550
rect 45089 56980 45090 58300
rect 46410 56980 46411 58300
rect 45089 56979 46411 56980
rect 41692 56912 41788 56928
rect 41692 56642 41788 56658
rect 40099 56590 41421 56591
rect 38170 56020 38310 56050
rect 38170 55960 38200 56020
rect 36782 55950 38200 55960
rect 38280 55950 38310 56020
rect 36782 55910 38310 55950
rect 36782 55900 38200 55910
rect 36782 55218 36798 55900
rect 38170 55840 38200 55900
rect 38280 55840 38310 55910
rect 38170 55800 38310 55840
rect 40099 55270 40100 56590
rect 41420 55270 41421 56590
rect 40099 55269 41421 55270
rect 36702 55202 36798 55218
rect 36702 54932 36798 54948
rect 35109 54880 36431 54881
rect 33180 54310 33320 54340
rect 33180 54250 33210 54310
rect 31792 54240 33210 54250
rect 33290 54240 33320 54310
rect 31792 54200 33320 54240
rect 31792 54190 33210 54200
rect 31792 53508 31808 54190
rect 33180 54130 33210 54190
rect 33290 54130 33320 54200
rect 34010 54190 34700 54250
rect 33180 54090 33320 54130
rect 35109 53560 35110 54880
rect 36430 53560 36431 54880
rect 35109 53559 36431 53560
rect 31712 53492 31808 53508
rect 31712 53222 31808 53238
rect 30119 53170 31441 53171
rect 28190 52600 28330 52630
rect 28190 52540 28220 52600
rect 26802 52530 28220 52540
rect 28300 52530 28330 52600
rect 26802 52490 28330 52530
rect 26802 52480 28220 52490
rect 26802 51798 26818 52480
rect 28190 52420 28220 52480
rect 28300 52420 28330 52490
rect 28190 52380 28330 52420
rect 30119 51850 30120 53170
rect 31440 51850 31441 53170
rect 30119 51849 31441 51850
rect 26722 51782 26818 51798
rect 26722 51512 26818 51528
rect 25129 51460 26451 51461
rect 23200 50890 23340 50920
rect 23200 50830 23230 50890
rect 21812 50820 23230 50830
rect 23310 50820 23340 50890
rect 21812 50780 23340 50820
rect 21812 50770 23230 50780
rect 21812 50088 21828 50770
rect 23200 50710 23230 50770
rect 23310 50710 23340 50780
rect 23200 50670 23340 50710
rect 25129 50140 25130 51460
rect 26450 50140 26451 51460
rect 25129 50139 26451 50140
rect 21732 50072 21828 50088
rect 21732 49802 21828 49818
rect 20139 49750 21461 49751
rect 18210 49180 18350 49210
rect 18210 49120 18240 49180
rect 16822 49110 18240 49120
rect 18320 49110 18350 49180
rect 16822 49070 18350 49110
rect 16822 49060 18240 49070
rect 16822 48378 16838 49060
rect 18210 49000 18240 49060
rect 18320 49000 18350 49070
rect 18210 48960 18350 49000
rect 20139 48430 20140 49750
rect 21460 48430 21461 49750
rect 20139 48429 21461 48430
rect 16742 48362 16838 48378
rect 16742 48092 16838 48108
rect 15149 48040 16471 48041
rect 13220 47470 13360 47500
rect 13220 47410 13250 47470
rect 11832 47400 13250 47410
rect 13330 47400 13360 47470
rect 11832 47360 13360 47400
rect 11832 47350 13250 47360
rect 11832 46668 11848 47350
rect 13220 47290 13250 47350
rect 13330 47290 13360 47360
rect 13220 47250 13360 47290
rect 15149 46720 15150 48040
rect 16470 46720 16471 48040
rect 15149 46719 16471 46720
rect 11752 46652 11848 46668
rect 11752 46382 11848 46398
rect 10159 46330 11481 46331
rect 8230 45760 8370 45790
rect 8230 45700 8260 45760
rect 6842 45690 8260 45700
rect 8340 45690 8370 45760
rect 6842 45650 8370 45690
rect 6842 45640 8260 45650
rect 6842 44958 6858 45640
rect 8230 45580 8260 45640
rect 8340 45580 8370 45650
rect 8230 45540 8370 45580
rect 10159 45010 10160 46330
rect 11480 45010 11481 46330
rect 10159 45009 11481 45010
rect 6762 44942 6858 44958
rect 6762 44672 6858 44688
rect 5169 44620 6491 44621
rect 3240 44050 3380 44080
rect 3240 43990 3270 44050
rect 1852 43980 3270 43990
rect 3350 43980 3380 44050
rect 1852 43940 3380 43980
rect 1852 43930 3270 43940
rect 1852 43248 1868 43930
rect 3240 43870 3270 43930
rect 3350 43870 3380 43940
rect 3240 43830 3380 43870
rect 5169 43300 5170 44620
rect 6490 43300 6491 44620
rect 5169 43299 6491 43300
rect 1772 43232 1868 43248
rect 1772 42962 1868 42978
rect 179 42910 1501 42911
rect 179 41590 180 42910
rect 1500 41590 1501 42910
rect 179 41589 1501 41590
rect 180 41201 240 41589
rect 1772 41538 1788 42962
rect 1852 42280 1868 42962
rect 5170 42911 5230 43299
rect 6762 43248 6778 44672
rect 6842 43990 6858 44672
rect 10160 44621 10220 45009
rect 11752 44958 11768 46382
rect 11832 45700 11848 46382
rect 15150 46331 15210 46719
rect 16742 46668 16758 48092
rect 16822 47410 16838 48092
rect 20140 48041 20200 48429
rect 21732 48378 21748 49802
rect 21812 49120 21828 49802
rect 25130 49751 25190 50139
rect 26722 50088 26738 51512
rect 26802 50830 26818 51512
rect 30120 51461 30180 51849
rect 31712 51798 31728 53222
rect 31792 52540 31808 53222
rect 35110 53171 35170 53559
rect 36702 53508 36718 54932
rect 36782 54250 36798 54932
rect 40100 54881 40160 55269
rect 41692 55218 41708 56642
rect 41772 55960 41788 56642
rect 45090 56591 45150 56979
rect 46682 56928 46698 58352
rect 46762 57670 46778 58352
rect 50080 58301 50140 58689
rect 51672 58638 51688 60062
rect 51752 59380 51768 60062
rect 55070 60011 55130 60399
rect 56662 60348 56678 61772
rect 56742 61090 56758 61772
rect 60060 61721 60120 62109
rect 61652 62058 61668 63482
rect 61732 62800 61748 63482
rect 65050 63431 65110 63819
rect 66642 63768 66658 65192
rect 66722 64510 66738 65192
rect 70040 65141 70100 65529
rect 71632 65478 71648 66902
rect 71712 66220 71728 66902
rect 75030 66851 75090 67110
rect 76622 66902 76718 66918
rect 75029 66850 76351 66851
rect 73100 66280 73240 66310
rect 73100 66220 73130 66280
rect 71712 66210 73130 66220
rect 73210 66210 73240 66280
rect 71712 66170 73240 66210
rect 71712 66160 73130 66170
rect 71712 65478 71728 66160
rect 73100 66100 73130 66160
rect 73210 66100 73240 66170
rect 73100 66060 73240 66100
rect 75029 65530 75030 66850
rect 76350 65530 76351 66850
rect 75029 65529 76351 65530
rect 71632 65462 71728 65478
rect 71632 65192 71728 65208
rect 70039 65140 71361 65141
rect 68110 64570 68250 64600
rect 68110 64510 68140 64570
rect 66722 64500 68140 64510
rect 68220 64500 68250 64570
rect 66722 64460 68250 64500
rect 66722 64450 68140 64460
rect 66722 63768 66738 64450
rect 68110 64390 68140 64450
rect 68220 64390 68250 64460
rect 68110 64350 68250 64390
rect 70039 63820 70040 65140
rect 71360 63820 71361 65140
rect 70039 63819 71361 63820
rect 66642 63752 66738 63768
rect 66642 63482 66738 63498
rect 65049 63430 66371 63431
rect 63120 62860 63260 62890
rect 63120 62800 63150 62860
rect 61732 62790 63150 62800
rect 63230 62790 63260 62860
rect 61732 62750 63260 62790
rect 61732 62740 63150 62750
rect 61732 62058 61748 62740
rect 63120 62680 63150 62740
rect 63230 62680 63260 62750
rect 63120 62640 63260 62680
rect 65049 62110 65050 63430
rect 66370 62110 66371 63430
rect 65049 62109 66371 62110
rect 61652 62042 61748 62058
rect 61652 61772 61748 61788
rect 60059 61720 61381 61721
rect 58130 61150 58270 61180
rect 58130 61090 58160 61150
rect 56742 61080 58160 61090
rect 58240 61080 58270 61150
rect 56742 61040 58270 61080
rect 56742 61030 58160 61040
rect 56742 60348 56758 61030
rect 58130 60970 58160 61030
rect 58240 60970 58270 61040
rect 58130 60930 58270 60970
rect 60059 60400 60060 61720
rect 61380 60400 61381 61720
rect 60059 60399 61381 60400
rect 56662 60332 56758 60348
rect 56662 60062 56758 60078
rect 55069 60010 56391 60011
rect 53140 59440 53280 59470
rect 53140 59380 53170 59440
rect 51752 59370 53170 59380
rect 53250 59370 53280 59440
rect 51752 59330 53280 59370
rect 51752 59320 53170 59330
rect 51752 58638 51768 59320
rect 53140 59260 53170 59320
rect 53250 59260 53280 59330
rect 53140 59220 53280 59260
rect 55069 58690 55070 60010
rect 56390 58690 56391 60010
rect 55069 58689 56391 58690
rect 51672 58622 51768 58638
rect 51672 58352 51768 58368
rect 50079 58300 51401 58301
rect 48150 57730 48290 57760
rect 48150 57670 48180 57730
rect 46762 57660 48180 57670
rect 48260 57660 48290 57730
rect 46762 57620 48290 57660
rect 46762 57610 48180 57620
rect 46762 56928 46778 57610
rect 48150 57550 48180 57610
rect 48260 57550 48290 57620
rect 48980 57610 49670 57670
rect 48150 57510 48290 57550
rect 50079 56980 50080 58300
rect 51400 56980 51401 58300
rect 50079 56979 51401 56980
rect 46682 56912 46778 56928
rect 46682 56642 46778 56658
rect 45089 56590 46411 56591
rect 43160 56020 43300 56050
rect 43160 55960 43190 56020
rect 41772 55950 43190 55960
rect 43270 55950 43300 56020
rect 41772 55910 43300 55950
rect 41772 55900 43190 55910
rect 41772 55218 41788 55900
rect 43160 55840 43190 55900
rect 43270 55840 43300 55910
rect 43160 55800 43300 55840
rect 45089 55270 45090 56590
rect 46410 55270 46411 56590
rect 45089 55269 46411 55270
rect 41692 55202 41788 55218
rect 41692 54932 41788 54948
rect 40099 54880 41421 54881
rect 38170 54310 38310 54340
rect 38170 54250 38200 54310
rect 36782 54240 38200 54250
rect 38280 54240 38310 54310
rect 36782 54200 38310 54240
rect 36782 54190 38200 54200
rect 36782 53508 36798 54190
rect 38170 54130 38200 54190
rect 38280 54130 38310 54200
rect 38170 54090 38310 54130
rect 40099 53560 40100 54880
rect 41420 53560 41421 54880
rect 40099 53559 41421 53560
rect 36702 53492 36798 53508
rect 36702 53222 36798 53238
rect 35109 53170 36431 53171
rect 33180 52600 33320 52630
rect 33180 52540 33210 52600
rect 31792 52530 33210 52540
rect 33290 52530 33320 52600
rect 31792 52490 33320 52530
rect 31792 52480 33210 52490
rect 31792 51798 31808 52480
rect 33180 52420 33210 52480
rect 33290 52420 33320 52490
rect 34010 52480 34700 52540
rect 33180 52380 33320 52420
rect 35109 51850 35110 53170
rect 36430 51850 36431 53170
rect 35109 51849 36431 51850
rect 31712 51782 31808 51798
rect 31712 51512 31808 51528
rect 30119 51460 31441 51461
rect 28190 50890 28330 50920
rect 28190 50830 28220 50890
rect 26802 50820 28220 50830
rect 28300 50820 28330 50890
rect 26802 50780 28330 50820
rect 26802 50770 28220 50780
rect 26802 50088 26818 50770
rect 28190 50710 28220 50770
rect 28300 50710 28330 50780
rect 28190 50670 28330 50710
rect 30119 50140 30120 51460
rect 31440 50140 31441 51460
rect 30119 50139 31441 50140
rect 26722 50072 26818 50088
rect 26722 49802 26818 49818
rect 25129 49750 26451 49751
rect 23200 49180 23340 49210
rect 23200 49120 23230 49180
rect 21812 49110 23230 49120
rect 23310 49110 23340 49180
rect 21812 49070 23340 49110
rect 21812 49060 23230 49070
rect 21812 48378 21828 49060
rect 23200 49000 23230 49060
rect 23310 49000 23340 49070
rect 23200 48960 23340 49000
rect 25129 48430 25130 49750
rect 26450 48430 26451 49750
rect 25129 48429 26451 48430
rect 21732 48362 21828 48378
rect 21732 48092 21828 48108
rect 20139 48040 21461 48041
rect 18210 47470 18350 47500
rect 18210 47410 18240 47470
rect 16822 47400 18240 47410
rect 18320 47400 18350 47470
rect 16822 47360 18350 47400
rect 16822 47350 18240 47360
rect 16822 46668 16838 47350
rect 18210 47290 18240 47350
rect 18320 47290 18350 47360
rect 18210 47250 18350 47290
rect 20139 46720 20140 48040
rect 21460 46720 21461 48040
rect 20139 46719 21461 46720
rect 16742 46652 16838 46668
rect 16742 46382 16838 46398
rect 15149 46330 16471 46331
rect 13220 45760 13360 45790
rect 13220 45700 13250 45760
rect 11832 45690 13250 45700
rect 13330 45690 13360 45760
rect 11832 45650 13360 45690
rect 11832 45640 13250 45650
rect 11832 44958 11848 45640
rect 13220 45580 13250 45640
rect 13330 45580 13360 45650
rect 13220 45540 13360 45580
rect 15149 45010 15150 46330
rect 16470 45010 16471 46330
rect 15149 45009 16471 45010
rect 11752 44942 11848 44958
rect 11752 44672 11848 44688
rect 10159 44620 11481 44621
rect 8230 44050 8370 44080
rect 8230 43990 8260 44050
rect 6842 43980 8260 43990
rect 8340 43980 8370 44050
rect 6842 43940 8370 43980
rect 6842 43930 8260 43940
rect 6842 43248 6858 43930
rect 8230 43870 8260 43930
rect 8340 43870 8370 43940
rect 8230 43830 8370 43870
rect 10159 43300 10160 44620
rect 11480 43300 11481 44620
rect 10159 43299 11481 43300
rect 6762 43232 6858 43248
rect 6762 42962 6858 42978
rect 5169 42910 6491 42911
rect 3240 42340 3380 42370
rect 3240 42280 3270 42340
rect 1852 42270 3270 42280
rect 3350 42270 3380 42340
rect 1852 42230 3380 42270
rect 1852 42220 3270 42230
rect 1852 41538 1868 42220
rect 3240 42160 3270 42220
rect 3350 42160 3380 42230
rect 3240 42120 3380 42160
rect 5169 41590 5170 42910
rect 6490 41590 6491 42910
rect 5169 41589 6491 41590
rect 1772 41522 1868 41538
rect 1772 41252 1868 41268
rect 179 41200 1501 41201
rect 179 39880 180 41200
rect 1500 39880 1501 41200
rect 179 39879 1501 39880
rect 180 39690 240 39879
rect 1772 39828 1788 41252
rect 1852 40570 1868 41252
rect 5170 41201 5230 41589
rect 6762 41538 6778 42962
rect 6842 42280 6858 42962
rect 10160 42911 10220 43299
rect 11752 43248 11768 44672
rect 11832 43990 11848 44672
rect 15150 44621 15210 45009
rect 16742 44958 16758 46382
rect 16822 45700 16838 46382
rect 20140 46331 20200 46719
rect 21732 46668 21748 48092
rect 21812 47410 21828 48092
rect 25130 48041 25190 48429
rect 26722 48378 26738 49802
rect 26802 49120 26818 49802
rect 30120 49751 30180 50139
rect 31712 50088 31728 51512
rect 31792 50830 31808 51512
rect 35110 51461 35170 51849
rect 36702 51798 36718 53222
rect 36782 52540 36798 53222
rect 40100 53171 40160 53559
rect 41692 53508 41708 54932
rect 41772 54250 41788 54932
rect 45090 54881 45150 55269
rect 46682 55218 46698 56642
rect 46762 55960 46778 56642
rect 50080 56591 50140 56979
rect 51672 56928 51688 58352
rect 51752 57670 51768 58352
rect 55070 58301 55130 58689
rect 56662 58638 56678 60062
rect 56742 59380 56758 60062
rect 60060 60011 60120 60399
rect 61652 60348 61668 61772
rect 61732 61090 61748 61772
rect 65050 61721 65110 62109
rect 66642 62058 66658 63482
rect 66722 62800 66738 63482
rect 70040 63431 70100 63819
rect 71632 63768 71648 65192
rect 71712 64510 71728 65192
rect 75030 65141 75090 65529
rect 76622 65478 76638 66902
rect 76702 66220 76718 66902
rect 78090 66280 78230 66310
rect 78090 66220 78120 66280
rect 76702 66210 78120 66220
rect 78200 66210 78230 66280
rect 76702 66170 78230 66210
rect 76702 66160 78120 66170
rect 76702 65478 76718 66160
rect 78090 66100 78120 66160
rect 78200 66100 78230 66170
rect 78090 66060 78230 66100
rect 76622 65462 76718 65478
rect 76622 65192 76718 65208
rect 75029 65140 76351 65141
rect 73100 64570 73240 64600
rect 73100 64510 73130 64570
rect 71712 64500 73130 64510
rect 73210 64500 73240 64570
rect 71712 64460 73240 64500
rect 71712 64450 73130 64460
rect 71712 63768 71728 64450
rect 73100 64390 73130 64450
rect 73210 64390 73240 64460
rect 73100 64350 73240 64390
rect 75029 63820 75030 65140
rect 76350 63820 76351 65140
rect 75029 63819 76351 63820
rect 71632 63752 71728 63768
rect 71632 63482 71728 63498
rect 70039 63430 71361 63431
rect 68110 62860 68250 62890
rect 68110 62800 68140 62860
rect 66722 62790 68140 62800
rect 68220 62790 68250 62860
rect 66722 62750 68250 62790
rect 66722 62740 68140 62750
rect 66722 62058 66738 62740
rect 68110 62680 68140 62740
rect 68220 62680 68250 62750
rect 68110 62640 68250 62680
rect 70039 62110 70040 63430
rect 71360 62110 71361 63430
rect 70039 62109 71361 62110
rect 66642 62042 66738 62058
rect 66642 61772 66738 61788
rect 65049 61720 66371 61721
rect 63120 61150 63260 61180
rect 63120 61090 63150 61150
rect 61732 61080 63150 61090
rect 63230 61080 63260 61150
rect 61732 61040 63260 61080
rect 61732 61030 63150 61040
rect 61732 60348 61748 61030
rect 63120 60970 63150 61030
rect 63230 60970 63260 61040
rect 63120 60930 63260 60970
rect 65049 60400 65050 61720
rect 66370 60400 66371 61720
rect 65049 60399 66371 60400
rect 61652 60332 61748 60348
rect 61652 60062 61748 60078
rect 60059 60010 61381 60011
rect 58130 59440 58270 59470
rect 58130 59380 58160 59440
rect 56742 59370 58160 59380
rect 58240 59370 58270 59440
rect 56742 59330 58270 59370
rect 56742 59320 58160 59330
rect 56742 58638 56758 59320
rect 58130 59260 58160 59320
rect 58240 59260 58270 59330
rect 58130 59220 58270 59260
rect 60059 58690 60060 60010
rect 61380 58690 61381 60010
rect 60059 58689 61381 58690
rect 56662 58622 56758 58638
rect 56662 58352 56758 58368
rect 55069 58300 56391 58301
rect 53140 57730 53280 57760
rect 53140 57670 53170 57730
rect 51752 57660 53170 57670
rect 53250 57660 53280 57730
rect 51752 57620 53280 57660
rect 51752 57610 53170 57620
rect 51752 56928 51768 57610
rect 53140 57550 53170 57610
rect 53250 57550 53280 57620
rect 53140 57510 53280 57550
rect 55069 56980 55070 58300
rect 56390 56980 56391 58300
rect 55069 56979 56391 56980
rect 51672 56912 51768 56928
rect 51672 56642 51768 56658
rect 50079 56590 51401 56591
rect 48150 56020 48290 56050
rect 48150 55960 48180 56020
rect 46762 55950 48180 55960
rect 48260 55950 48290 56020
rect 46762 55910 48290 55950
rect 46762 55900 48180 55910
rect 46762 55218 46778 55900
rect 48150 55840 48180 55900
rect 48260 55840 48290 55910
rect 48980 55900 49670 55960
rect 48150 55800 48290 55840
rect 50079 55270 50080 56590
rect 51400 55270 51401 56590
rect 50079 55269 51401 55270
rect 46682 55202 46778 55218
rect 46682 54932 46778 54948
rect 45089 54880 46411 54881
rect 43160 54310 43300 54340
rect 43160 54250 43190 54310
rect 41772 54240 43190 54250
rect 43270 54240 43300 54310
rect 41772 54200 43300 54240
rect 41772 54190 43190 54200
rect 41772 53508 41788 54190
rect 43160 54130 43190 54190
rect 43270 54130 43300 54200
rect 43160 54090 43300 54130
rect 45089 53560 45090 54880
rect 46410 53560 46411 54880
rect 45089 53559 46411 53560
rect 41692 53492 41788 53508
rect 41692 53222 41788 53238
rect 40099 53170 41421 53171
rect 38170 52600 38310 52630
rect 38170 52540 38200 52600
rect 36782 52530 38200 52540
rect 38280 52530 38310 52600
rect 36782 52490 38310 52530
rect 36782 52480 38200 52490
rect 36782 51798 36798 52480
rect 38170 52420 38200 52480
rect 38280 52420 38310 52490
rect 38170 52380 38310 52420
rect 40099 51850 40100 53170
rect 41420 51850 41421 53170
rect 40099 51849 41421 51850
rect 36702 51782 36798 51798
rect 36702 51512 36798 51528
rect 35109 51460 36431 51461
rect 33180 50890 33320 50920
rect 33180 50830 33210 50890
rect 31792 50820 33210 50830
rect 33290 50820 33320 50890
rect 31792 50780 33320 50820
rect 31792 50770 33210 50780
rect 31792 50088 31808 50770
rect 33180 50710 33210 50770
rect 33290 50710 33320 50780
rect 34010 50770 34700 50830
rect 33180 50670 33320 50710
rect 35109 50140 35110 51460
rect 36430 50140 36431 51460
rect 35109 50139 36431 50140
rect 31712 50072 31808 50088
rect 31712 49802 31808 49818
rect 30119 49750 31441 49751
rect 28190 49180 28330 49210
rect 28190 49120 28220 49180
rect 26802 49110 28220 49120
rect 28300 49110 28330 49180
rect 26802 49070 28330 49110
rect 26802 49060 28220 49070
rect 26802 48378 26818 49060
rect 28190 49000 28220 49060
rect 28300 49000 28330 49070
rect 28190 48960 28330 49000
rect 30119 48430 30120 49750
rect 31440 48430 31441 49750
rect 30119 48429 31441 48430
rect 26722 48362 26818 48378
rect 26722 48092 26818 48108
rect 25129 48040 26451 48041
rect 23200 47470 23340 47500
rect 23200 47410 23230 47470
rect 21812 47400 23230 47410
rect 23310 47400 23340 47470
rect 21812 47360 23340 47400
rect 21812 47350 23230 47360
rect 21812 46668 21828 47350
rect 23200 47290 23230 47350
rect 23310 47290 23340 47360
rect 23200 47250 23340 47290
rect 25129 46720 25130 48040
rect 26450 46720 26451 48040
rect 25129 46719 26451 46720
rect 21732 46652 21828 46668
rect 21732 46382 21828 46398
rect 20139 46330 21461 46331
rect 18210 45760 18350 45790
rect 18210 45700 18240 45760
rect 16822 45690 18240 45700
rect 18320 45690 18350 45760
rect 16822 45650 18350 45690
rect 16822 45640 18240 45650
rect 16822 44958 16838 45640
rect 18210 45580 18240 45640
rect 18320 45580 18350 45650
rect 18210 45540 18350 45580
rect 20139 45010 20140 46330
rect 21460 45010 21461 46330
rect 20139 45009 21461 45010
rect 16742 44942 16838 44958
rect 16742 44672 16838 44688
rect 15149 44620 16471 44621
rect 13220 44050 13360 44080
rect 13220 43990 13250 44050
rect 11832 43980 13250 43990
rect 13330 43980 13360 44050
rect 11832 43940 13360 43980
rect 11832 43930 13250 43940
rect 11832 43248 11848 43930
rect 13220 43870 13250 43930
rect 13330 43870 13360 43940
rect 13220 43830 13360 43870
rect 15149 43300 15150 44620
rect 16470 43300 16471 44620
rect 15149 43299 16471 43300
rect 11752 43232 11848 43248
rect 11752 42962 11848 42978
rect 10159 42910 11481 42911
rect 8230 42340 8370 42370
rect 8230 42280 8260 42340
rect 6842 42270 8260 42280
rect 8340 42270 8370 42340
rect 6842 42230 8370 42270
rect 6842 42220 8260 42230
rect 6842 41538 6858 42220
rect 8230 42160 8260 42220
rect 8340 42160 8370 42230
rect 8230 42120 8370 42160
rect 10159 41590 10160 42910
rect 11480 41590 11481 42910
rect 10159 41589 11481 41590
rect 6762 41522 6858 41538
rect 6762 41252 6858 41268
rect 5169 41200 6491 41201
rect 3240 40630 3380 40660
rect 3240 40570 3270 40630
rect 1852 40560 3270 40570
rect 3350 40560 3380 40630
rect 1852 40520 3380 40560
rect 1852 40510 3270 40520
rect 1852 39828 1868 40510
rect 3240 40450 3270 40510
rect 3350 40450 3380 40520
rect 3240 40410 3380 40450
rect 5169 39880 5170 41200
rect 6490 39880 6491 41200
rect 5169 39879 6491 39880
rect 1772 39812 1868 39828
rect 5170 39690 5230 39879
rect 6762 39828 6778 41252
rect 6842 40570 6858 41252
rect 10160 41201 10220 41589
rect 11752 41538 11768 42962
rect 11832 42280 11848 42962
rect 15150 42911 15210 43299
rect 16742 43248 16758 44672
rect 16822 43990 16838 44672
rect 20140 44621 20200 45009
rect 21732 44958 21748 46382
rect 21812 45700 21828 46382
rect 25130 46331 25190 46719
rect 26722 46668 26738 48092
rect 26802 47410 26818 48092
rect 30120 48041 30180 48429
rect 31712 48378 31728 49802
rect 31792 49120 31808 49802
rect 35110 49751 35170 50139
rect 36702 50088 36718 51512
rect 36782 50830 36798 51512
rect 40100 51461 40160 51849
rect 41692 51798 41708 53222
rect 41772 52540 41788 53222
rect 45090 53171 45150 53559
rect 46682 53508 46698 54932
rect 46762 54250 46778 54932
rect 50080 54881 50140 55269
rect 51672 55218 51688 56642
rect 51752 55960 51768 56642
rect 55070 56591 55130 56979
rect 56662 56928 56678 58352
rect 56742 57670 56758 58352
rect 60060 58301 60120 58689
rect 61652 58638 61668 60062
rect 61732 59380 61748 60062
rect 65050 60011 65110 60399
rect 66642 60348 66658 61772
rect 66722 61090 66738 61772
rect 70040 61721 70100 62109
rect 71632 62058 71648 63482
rect 71712 62800 71728 63482
rect 75030 63431 75090 63819
rect 76622 63768 76638 65192
rect 76702 64510 76718 65192
rect 78090 64570 78230 64600
rect 78090 64510 78120 64570
rect 76702 64500 78120 64510
rect 78200 64500 78230 64570
rect 76702 64460 78230 64500
rect 76702 64450 78120 64460
rect 76702 63768 76718 64450
rect 78090 64390 78120 64450
rect 78200 64390 78230 64460
rect 78090 64350 78230 64390
rect 76622 63752 76718 63768
rect 76622 63482 76718 63498
rect 75029 63430 76351 63431
rect 73100 62860 73240 62890
rect 73100 62800 73130 62860
rect 71712 62790 73130 62800
rect 73210 62790 73240 62860
rect 71712 62750 73240 62790
rect 71712 62740 73130 62750
rect 71712 62058 71728 62740
rect 73100 62680 73130 62740
rect 73210 62680 73240 62750
rect 73100 62640 73240 62680
rect 75029 62110 75030 63430
rect 76350 62110 76351 63430
rect 75029 62109 76351 62110
rect 71632 62042 71728 62058
rect 71632 61772 71728 61788
rect 70039 61720 71361 61721
rect 68110 61150 68250 61180
rect 68110 61090 68140 61150
rect 66722 61080 68140 61090
rect 68220 61080 68250 61150
rect 66722 61040 68250 61080
rect 66722 61030 68140 61040
rect 66722 60348 66738 61030
rect 68110 60970 68140 61030
rect 68220 60970 68250 61040
rect 68110 60930 68250 60970
rect 70039 60400 70040 61720
rect 71360 60400 71361 61720
rect 70039 60399 71361 60400
rect 66642 60332 66738 60348
rect 66642 60062 66738 60078
rect 65049 60010 66371 60011
rect 63120 59440 63260 59470
rect 63120 59380 63150 59440
rect 61732 59370 63150 59380
rect 63230 59370 63260 59440
rect 61732 59330 63260 59370
rect 61732 59320 63150 59330
rect 61732 58638 61748 59320
rect 63120 59260 63150 59320
rect 63230 59260 63260 59330
rect 63120 59220 63260 59260
rect 65049 58690 65050 60010
rect 66370 58690 66371 60010
rect 65049 58689 66371 58690
rect 61652 58622 61748 58638
rect 61652 58352 61748 58368
rect 60059 58300 61381 58301
rect 58130 57730 58270 57760
rect 58130 57670 58160 57730
rect 56742 57660 58160 57670
rect 58240 57660 58270 57730
rect 56742 57620 58270 57660
rect 56742 57610 58160 57620
rect 56742 56928 56758 57610
rect 58130 57550 58160 57610
rect 58240 57550 58270 57620
rect 58130 57510 58270 57550
rect 60059 56980 60060 58300
rect 61380 56980 61381 58300
rect 60059 56979 61381 56980
rect 56662 56912 56758 56928
rect 56662 56642 56758 56658
rect 55069 56590 56391 56591
rect 53140 56020 53280 56050
rect 53140 55960 53170 56020
rect 51752 55950 53170 55960
rect 53250 55950 53280 56020
rect 51752 55910 53280 55950
rect 51752 55900 53170 55910
rect 51752 55218 51768 55900
rect 53140 55840 53170 55900
rect 53250 55840 53280 55910
rect 53140 55800 53280 55840
rect 55069 55270 55070 56590
rect 56390 55270 56391 56590
rect 55069 55269 56391 55270
rect 51672 55202 51768 55218
rect 51672 54932 51768 54948
rect 50079 54880 51401 54881
rect 48150 54310 48290 54340
rect 48150 54250 48180 54310
rect 46762 54240 48180 54250
rect 48260 54240 48290 54310
rect 46762 54200 48290 54240
rect 46762 54190 48180 54200
rect 46762 53508 46778 54190
rect 48150 54130 48180 54190
rect 48260 54130 48290 54200
rect 48980 54190 49670 54250
rect 48150 54090 48290 54130
rect 50079 53560 50080 54880
rect 51400 53560 51401 54880
rect 50079 53559 51401 53560
rect 46682 53492 46778 53508
rect 46682 53222 46778 53238
rect 45089 53170 46411 53171
rect 43160 52600 43300 52630
rect 43160 52540 43190 52600
rect 41772 52530 43190 52540
rect 43270 52530 43300 52600
rect 41772 52490 43300 52530
rect 41772 52480 43190 52490
rect 41772 51798 41788 52480
rect 43160 52420 43190 52480
rect 43270 52420 43300 52490
rect 43160 52380 43300 52420
rect 45089 51850 45090 53170
rect 46410 51850 46411 53170
rect 45089 51849 46411 51850
rect 41692 51782 41788 51798
rect 41692 51512 41788 51528
rect 40099 51460 41421 51461
rect 38170 50890 38310 50920
rect 38170 50830 38200 50890
rect 36782 50820 38200 50830
rect 38280 50820 38310 50890
rect 36782 50780 38310 50820
rect 36782 50770 38200 50780
rect 36782 50088 36798 50770
rect 38170 50710 38200 50770
rect 38280 50710 38310 50780
rect 38170 50670 38310 50710
rect 40099 50140 40100 51460
rect 41420 50140 41421 51460
rect 40099 50139 41421 50140
rect 36702 50072 36798 50088
rect 36702 49802 36798 49818
rect 35109 49750 36431 49751
rect 33180 49180 33320 49210
rect 33180 49120 33210 49180
rect 31792 49110 33210 49120
rect 33290 49110 33320 49180
rect 31792 49070 33320 49110
rect 31792 49060 33210 49070
rect 31792 48378 31808 49060
rect 33180 49000 33210 49060
rect 33290 49000 33320 49070
rect 34010 49060 34700 49120
rect 33180 48960 33320 49000
rect 35109 48430 35110 49750
rect 36430 48430 36431 49750
rect 35109 48429 36431 48430
rect 31712 48362 31808 48378
rect 31712 48092 31808 48108
rect 30119 48040 31441 48041
rect 28190 47470 28330 47500
rect 28190 47410 28220 47470
rect 26802 47400 28220 47410
rect 28300 47400 28330 47470
rect 26802 47360 28330 47400
rect 26802 47350 28220 47360
rect 26802 46668 26818 47350
rect 28190 47290 28220 47350
rect 28300 47290 28330 47360
rect 28190 47250 28330 47290
rect 30119 46720 30120 48040
rect 31440 46720 31441 48040
rect 30119 46719 31441 46720
rect 26722 46652 26818 46668
rect 26722 46382 26818 46398
rect 25129 46330 26451 46331
rect 23200 45760 23340 45790
rect 23200 45700 23230 45760
rect 21812 45690 23230 45700
rect 23310 45690 23340 45760
rect 21812 45650 23340 45690
rect 21812 45640 23230 45650
rect 21812 44958 21828 45640
rect 23200 45580 23230 45640
rect 23310 45580 23340 45650
rect 23200 45540 23340 45580
rect 25129 45010 25130 46330
rect 26450 45010 26451 46330
rect 25129 45009 26451 45010
rect 21732 44942 21828 44958
rect 21732 44672 21828 44688
rect 20139 44620 21461 44621
rect 18210 44050 18350 44080
rect 18210 43990 18240 44050
rect 16822 43980 18240 43990
rect 18320 43980 18350 44050
rect 16822 43940 18350 43980
rect 16822 43930 18240 43940
rect 16822 43248 16838 43930
rect 18210 43870 18240 43930
rect 18320 43870 18350 43940
rect 18210 43830 18350 43870
rect 20139 43300 20140 44620
rect 21460 43300 21461 44620
rect 20139 43299 21461 43300
rect 16742 43232 16838 43248
rect 16742 42962 16838 42978
rect 15149 42910 16471 42911
rect 13220 42340 13360 42370
rect 13220 42280 13250 42340
rect 11832 42270 13250 42280
rect 13330 42270 13360 42340
rect 11832 42230 13360 42270
rect 11832 42220 13250 42230
rect 11832 41538 11848 42220
rect 13220 42160 13250 42220
rect 13330 42160 13360 42230
rect 13220 42120 13360 42160
rect 15149 41590 15150 42910
rect 16470 41590 16471 42910
rect 15149 41589 16471 41590
rect 11752 41522 11848 41538
rect 11752 41252 11848 41268
rect 10159 41200 11481 41201
rect 8230 40630 8370 40660
rect 8230 40570 8260 40630
rect 6842 40560 8260 40570
rect 8340 40560 8370 40630
rect 6842 40520 8370 40560
rect 6842 40510 8260 40520
rect 6842 39828 6858 40510
rect 8230 40450 8260 40510
rect 8340 40450 8370 40520
rect 8230 40410 8370 40450
rect 10159 39880 10160 41200
rect 11480 39880 11481 41200
rect 10159 39879 11481 39880
rect 6762 39812 6858 39828
rect 10160 39690 10220 39879
rect 11752 39828 11768 41252
rect 11832 40570 11848 41252
rect 15150 41201 15210 41589
rect 16742 41538 16758 42962
rect 16822 42280 16838 42962
rect 20140 42911 20200 43299
rect 21732 43248 21748 44672
rect 21812 43990 21828 44672
rect 25130 44621 25190 45009
rect 26722 44958 26738 46382
rect 26802 45700 26818 46382
rect 30120 46331 30180 46719
rect 31712 46668 31728 48092
rect 31792 47410 31808 48092
rect 35110 48041 35170 48429
rect 36702 48378 36718 49802
rect 36782 49120 36798 49802
rect 40100 49751 40160 50139
rect 41692 50088 41708 51512
rect 41772 50830 41788 51512
rect 45090 51461 45150 51849
rect 46682 51798 46698 53222
rect 46762 52540 46778 53222
rect 50080 53171 50140 53559
rect 51672 53508 51688 54932
rect 51752 54250 51768 54932
rect 55070 54881 55130 55269
rect 56662 55218 56678 56642
rect 56742 55960 56758 56642
rect 60060 56591 60120 56979
rect 61652 56928 61668 58352
rect 61732 57670 61748 58352
rect 65050 58301 65110 58689
rect 66642 58638 66658 60062
rect 66722 59380 66738 60062
rect 70040 60011 70100 60399
rect 71632 60348 71648 61772
rect 71712 61090 71728 61772
rect 75030 61721 75090 62109
rect 76622 62058 76638 63482
rect 76702 62800 76718 63482
rect 78090 62860 78230 62890
rect 78090 62800 78120 62860
rect 76702 62790 78120 62800
rect 78200 62790 78230 62860
rect 76702 62750 78230 62790
rect 76702 62740 78120 62750
rect 76702 62058 76718 62740
rect 78090 62680 78120 62740
rect 78200 62680 78230 62750
rect 78090 62640 78230 62680
rect 76622 62042 76718 62058
rect 76622 61772 76718 61788
rect 75029 61720 76351 61721
rect 73100 61150 73240 61180
rect 73100 61090 73130 61150
rect 71712 61080 73130 61090
rect 73210 61080 73240 61150
rect 71712 61040 73240 61080
rect 71712 61030 73130 61040
rect 71712 60348 71728 61030
rect 73100 60970 73130 61030
rect 73210 60970 73240 61040
rect 73100 60930 73240 60970
rect 75029 60400 75030 61720
rect 76350 60400 76351 61720
rect 75029 60399 76351 60400
rect 71632 60332 71728 60348
rect 71632 60062 71728 60078
rect 70039 60010 71361 60011
rect 68110 59440 68250 59470
rect 68110 59380 68140 59440
rect 66722 59370 68140 59380
rect 68220 59370 68250 59440
rect 66722 59330 68250 59370
rect 66722 59320 68140 59330
rect 66722 58638 66738 59320
rect 68110 59260 68140 59320
rect 68220 59260 68250 59330
rect 68110 59220 68250 59260
rect 70039 58690 70040 60010
rect 71360 58690 71361 60010
rect 70039 58689 71361 58690
rect 66642 58622 66738 58638
rect 66642 58352 66738 58368
rect 65049 58300 66371 58301
rect 63120 57730 63260 57760
rect 63120 57670 63150 57730
rect 61732 57660 63150 57670
rect 63230 57660 63260 57730
rect 61732 57620 63260 57660
rect 61732 57610 63150 57620
rect 61732 56928 61748 57610
rect 63120 57550 63150 57610
rect 63230 57550 63260 57620
rect 63120 57510 63260 57550
rect 65049 56980 65050 58300
rect 66370 56980 66371 58300
rect 65049 56979 66371 56980
rect 61652 56912 61748 56928
rect 61652 56642 61748 56658
rect 60059 56590 61381 56591
rect 58130 56020 58270 56050
rect 58130 55960 58160 56020
rect 56742 55950 58160 55960
rect 58240 55950 58270 56020
rect 56742 55910 58270 55950
rect 56742 55900 58160 55910
rect 56742 55218 56758 55900
rect 58130 55840 58160 55900
rect 58240 55840 58270 55910
rect 58130 55800 58270 55840
rect 60059 55270 60060 56590
rect 61380 55270 61381 56590
rect 60059 55269 61381 55270
rect 56662 55202 56758 55218
rect 56662 54932 56758 54948
rect 55069 54880 56391 54881
rect 53140 54310 53280 54340
rect 53140 54250 53170 54310
rect 51752 54240 53170 54250
rect 53250 54240 53280 54310
rect 51752 54200 53280 54240
rect 51752 54190 53170 54200
rect 51752 53508 51768 54190
rect 53140 54130 53170 54190
rect 53250 54130 53280 54200
rect 53140 54090 53280 54130
rect 55069 53560 55070 54880
rect 56390 53560 56391 54880
rect 55069 53559 56391 53560
rect 51672 53492 51768 53508
rect 51672 53222 51768 53238
rect 50079 53170 51401 53171
rect 48150 52600 48290 52630
rect 48150 52540 48180 52600
rect 46762 52530 48180 52540
rect 48260 52530 48290 52600
rect 46762 52490 48290 52530
rect 46762 52480 48180 52490
rect 46762 51798 46778 52480
rect 48150 52420 48180 52480
rect 48260 52420 48290 52490
rect 48980 52480 49670 52540
rect 48150 52380 48290 52420
rect 50079 51850 50080 53170
rect 51400 51850 51401 53170
rect 50079 51849 51401 51850
rect 46682 51782 46778 51798
rect 46682 51512 46778 51528
rect 45089 51460 46411 51461
rect 43160 50890 43300 50920
rect 43160 50830 43190 50890
rect 41772 50820 43190 50830
rect 43270 50820 43300 50890
rect 41772 50780 43300 50820
rect 41772 50770 43190 50780
rect 41772 50088 41788 50770
rect 43160 50710 43190 50770
rect 43270 50710 43300 50780
rect 43160 50670 43300 50710
rect 45089 50140 45090 51460
rect 46410 50140 46411 51460
rect 45089 50139 46411 50140
rect 41692 50072 41788 50088
rect 41692 49802 41788 49818
rect 40099 49750 41421 49751
rect 38170 49180 38310 49210
rect 38170 49120 38200 49180
rect 36782 49110 38200 49120
rect 38280 49110 38310 49180
rect 36782 49070 38310 49110
rect 36782 49060 38200 49070
rect 36782 48378 36798 49060
rect 38170 49000 38200 49060
rect 38280 49000 38310 49070
rect 38170 48960 38310 49000
rect 40099 48430 40100 49750
rect 41420 48430 41421 49750
rect 40099 48429 41421 48430
rect 36702 48362 36798 48378
rect 36702 48092 36798 48108
rect 35109 48040 36431 48041
rect 33180 47470 33320 47500
rect 33180 47410 33210 47470
rect 31792 47400 33210 47410
rect 33290 47400 33320 47470
rect 31792 47360 33320 47400
rect 31792 47350 33210 47360
rect 31792 46668 31808 47350
rect 33180 47290 33210 47350
rect 33290 47290 33320 47360
rect 34010 47350 34700 47410
rect 33180 47250 33320 47290
rect 35109 46720 35110 48040
rect 36430 46720 36431 48040
rect 35109 46719 36431 46720
rect 31712 46652 31808 46668
rect 31712 46382 31808 46398
rect 30119 46330 31441 46331
rect 28190 45760 28330 45790
rect 28190 45700 28220 45760
rect 26802 45690 28220 45700
rect 28300 45690 28330 45760
rect 26802 45650 28330 45690
rect 26802 45640 28220 45650
rect 26802 44958 26818 45640
rect 28190 45580 28220 45640
rect 28300 45580 28330 45650
rect 28190 45540 28330 45580
rect 30119 45010 30120 46330
rect 31440 45010 31441 46330
rect 30119 45009 31441 45010
rect 26722 44942 26818 44958
rect 26722 44672 26818 44688
rect 25129 44620 26451 44621
rect 23200 44050 23340 44080
rect 23200 43990 23230 44050
rect 21812 43980 23230 43990
rect 23310 43980 23340 44050
rect 21812 43940 23340 43980
rect 21812 43930 23230 43940
rect 21812 43248 21828 43930
rect 23200 43870 23230 43930
rect 23310 43870 23340 43940
rect 23200 43830 23340 43870
rect 25129 43300 25130 44620
rect 26450 43300 26451 44620
rect 25129 43299 26451 43300
rect 21732 43232 21828 43248
rect 21732 42962 21828 42978
rect 20139 42910 21461 42911
rect 18210 42340 18350 42370
rect 18210 42280 18240 42340
rect 16822 42270 18240 42280
rect 18320 42270 18350 42340
rect 16822 42230 18350 42270
rect 16822 42220 18240 42230
rect 16822 41538 16838 42220
rect 18210 42160 18240 42220
rect 18320 42160 18350 42230
rect 18210 42120 18350 42160
rect 20139 41590 20140 42910
rect 21460 41590 21461 42910
rect 20139 41589 21461 41590
rect 16742 41522 16838 41538
rect 16742 41252 16838 41268
rect 15149 41200 16471 41201
rect 13220 40630 13360 40660
rect 13220 40570 13250 40630
rect 11832 40560 13250 40570
rect 13330 40560 13360 40630
rect 11832 40520 13360 40560
rect 11832 40510 13250 40520
rect 11832 39828 11848 40510
rect 13220 40450 13250 40510
rect 13330 40450 13360 40520
rect 13220 40410 13360 40450
rect 15149 39880 15150 41200
rect 16470 39880 16471 41200
rect 15149 39879 16471 39880
rect 11752 39812 11848 39828
rect 15150 39690 15210 39879
rect 16742 39828 16758 41252
rect 16822 40570 16838 41252
rect 20140 41201 20200 41589
rect 21732 41538 21748 42962
rect 21812 42280 21828 42962
rect 25130 42911 25190 43299
rect 26722 43248 26738 44672
rect 26802 43990 26818 44672
rect 30120 44621 30180 45009
rect 31712 44958 31728 46382
rect 31792 45700 31808 46382
rect 35110 46331 35170 46719
rect 36702 46668 36718 48092
rect 36782 47410 36798 48092
rect 40100 48041 40160 48429
rect 41692 48378 41708 49802
rect 41772 49120 41788 49802
rect 45090 49751 45150 50139
rect 46682 50088 46698 51512
rect 46762 50830 46778 51512
rect 50080 51461 50140 51849
rect 51672 51798 51688 53222
rect 51752 52540 51768 53222
rect 55070 53171 55130 53559
rect 56662 53508 56678 54932
rect 56742 54250 56758 54932
rect 60060 54881 60120 55269
rect 61652 55218 61668 56642
rect 61732 55960 61748 56642
rect 65050 56591 65110 56979
rect 66642 56928 66658 58352
rect 66722 57670 66738 58352
rect 70040 58301 70100 58689
rect 71632 58638 71648 60062
rect 71712 59380 71728 60062
rect 75030 60011 75090 60399
rect 76622 60348 76638 61772
rect 76702 61090 76718 61772
rect 78090 61150 78230 61180
rect 78090 61090 78120 61150
rect 76702 61080 78120 61090
rect 78200 61080 78230 61150
rect 76702 61040 78230 61080
rect 76702 61030 78120 61040
rect 76702 60348 76718 61030
rect 78090 60970 78120 61030
rect 78200 60970 78230 61040
rect 78090 60930 78230 60970
rect 76622 60332 76718 60348
rect 76622 60062 76718 60078
rect 75029 60010 76351 60011
rect 73100 59440 73240 59470
rect 73100 59380 73130 59440
rect 71712 59370 73130 59380
rect 73210 59370 73240 59440
rect 71712 59330 73240 59370
rect 71712 59320 73130 59330
rect 71712 58638 71728 59320
rect 73100 59260 73130 59320
rect 73210 59260 73240 59330
rect 73100 59220 73240 59260
rect 75029 58690 75030 60010
rect 76350 58690 76351 60010
rect 75029 58689 76351 58690
rect 71632 58622 71728 58638
rect 71632 58352 71728 58368
rect 70039 58300 71361 58301
rect 68110 57730 68250 57760
rect 68110 57670 68140 57730
rect 66722 57660 68140 57670
rect 68220 57660 68250 57730
rect 66722 57620 68250 57660
rect 66722 57610 68140 57620
rect 66722 56928 66738 57610
rect 68110 57550 68140 57610
rect 68220 57550 68250 57620
rect 68110 57510 68250 57550
rect 70039 56980 70040 58300
rect 71360 56980 71361 58300
rect 70039 56979 71361 56980
rect 66642 56912 66738 56928
rect 66642 56642 66738 56658
rect 65049 56590 66371 56591
rect 63120 56020 63260 56050
rect 63120 55960 63150 56020
rect 61732 55950 63150 55960
rect 63230 55950 63260 56020
rect 61732 55910 63260 55950
rect 61732 55900 63150 55910
rect 61732 55218 61748 55900
rect 63120 55840 63150 55900
rect 63230 55840 63260 55910
rect 63120 55800 63260 55840
rect 65049 55270 65050 56590
rect 66370 55270 66371 56590
rect 65049 55269 66371 55270
rect 61652 55202 61748 55218
rect 61652 54932 61748 54948
rect 60059 54880 61381 54881
rect 58130 54310 58270 54340
rect 58130 54250 58160 54310
rect 56742 54240 58160 54250
rect 58240 54240 58270 54310
rect 56742 54200 58270 54240
rect 56742 54190 58160 54200
rect 56742 53508 56758 54190
rect 58130 54130 58160 54190
rect 58240 54130 58270 54200
rect 58130 54090 58270 54130
rect 60059 53560 60060 54880
rect 61380 53560 61381 54880
rect 60059 53559 61381 53560
rect 56662 53492 56758 53508
rect 56662 53222 56758 53238
rect 55069 53170 56391 53171
rect 53140 52600 53280 52630
rect 53140 52540 53170 52600
rect 51752 52530 53170 52540
rect 53250 52530 53280 52600
rect 51752 52490 53280 52530
rect 51752 52480 53170 52490
rect 51752 51798 51768 52480
rect 53140 52420 53170 52480
rect 53250 52420 53280 52490
rect 53140 52380 53280 52420
rect 55069 51850 55070 53170
rect 56390 51850 56391 53170
rect 55069 51849 56391 51850
rect 51672 51782 51768 51798
rect 51672 51512 51768 51528
rect 50079 51460 51401 51461
rect 48150 50890 48290 50920
rect 48150 50830 48180 50890
rect 46762 50820 48180 50830
rect 48260 50820 48290 50890
rect 46762 50780 48290 50820
rect 46762 50770 48180 50780
rect 46762 50088 46778 50770
rect 48150 50710 48180 50770
rect 48260 50710 48290 50780
rect 48980 50770 49670 50830
rect 48150 50670 48290 50710
rect 50079 50140 50080 51460
rect 51400 50140 51401 51460
rect 50079 50139 51401 50140
rect 46682 50072 46778 50088
rect 46682 49802 46778 49818
rect 45089 49750 46411 49751
rect 43160 49180 43300 49210
rect 43160 49120 43190 49180
rect 41772 49110 43190 49120
rect 43270 49110 43300 49180
rect 41772 49070 43300 49110
rect 41772 49060 43190 49070
rect 41772 48378 41788 49060
rect 43160 49000 43190 49060
rect 43270 49000 43300 49070
rect 43160 48960 43300 49000
rect 45089 48430 45090 49750
rect 46410 48430 46411 49750
rect 45089 48429 46411 48430
rect 41692 48362 41788 48378
rect 41692 48092 41788 48108
rect 40099 48040 41421 48041
rect 38170 47470 38310 47500
rect 38170 47410 38200 47470
rect 36782 47400 38200 47410
rect 38280 47400 38310 47470
rect 36782 47360 38310 47400
rect 36782 47350 38200 47360
rect 36782 46668 36798 47350
rect 38170 47290 38200 47350
rect 38280 47290 38310 47360
rect 38170 47250 38310 47290
rect 40099 46720 40100 48040
rect 41420 46720 41421 48040
rect 40099 46719 41421 46720
rect 36702 46652 36798 46668
rect 36702 46382 36798 46398
rect 35109 46330 36431 46331
rect 33180 45760 33320 45790
rect 33180 45700 33210 45760
rect 31792 45690 33210 45700
rect 33290 45690 33320 45760
rect 31792 45650 33320 45690
rect 31792 45640 33210 45650
rect 31792 44958 31808 45640
rect 33180 45580 33210 45640
rect 33290 45580 33320 45650
rect 34010 45640 34700 45700
rect 33180 45540 33320 45580
rect 35109 45010 35110 46330
rect 36430 45010 36431 46330
rect 35109 45009 36431 45010
rect 31712 44942 31808 44958
rect 31712 44672 31808 44688
rect 30119 44620 31441 44621
rect 28190 44050 28330 44080
rect 28190 43990 28220 44050
rect 26802 43980 28220 43990
rect 28300 43980 28330 44050
rect 26802 43940 28330 43980
rect 26802 43930 28220 43940
rect 26802 43248 26818 43930
rect 28190 43870 28220 43930
rect 28300 43870 28330 43940
rect 28190 43830 28330 43870
rect 30119 43300 30120 44620
rect 31440 43300 31441 44620
rect 30119 43299 31441 43300
rect 26722 43232 26818 43248
rect 26722 42962 26818 42978
rect 25129 42910 26451 42911
rect 23200 42340 23340 42370
rect 23200 42280 23230 42340
rect 21812 42270 23230 42280
rect 23310 42270 23340 42340
rect 21812 42230 23340 42270
rect 21812 42220 23230 42230
rect 21812 41538 21828 42220
rect 23200 42160 23230 42220
rect 23310 42160 23340 42230
rect 23200 42120 23340 42160
rect 25129 41590 25130 42910
rect 26450 41590 26451 42910
rect 25129 41589 26451 41590
rect 21732 41522 21828 41538
rect 21732 41252 21828 41268
rect 20139 41200 21461 41201
rect 18210 40630 18350 40660
rect 18210 40570 18240 40630
rect 16822 40560 18240 40570
rect 18320 40560 18350 40630
rect 16822 40520 18350 40560
rect 16822 40510 18240 40520
rect 16822 39828 16838 40510
rect 18210 40450 18240 40510
rect 18320 40450 18350 40520
rect 18210 40410 18350 40450
rect 20139 39880 20140 41200
rect 21460 39880 21461 41200
rect 20139 39879 21461 39880
rect 16742 39812 16838 39828
rect 20140 39690 20200 39879
rect 21732 39828 21748 41252
rect 21812 40570 21828 41252
rect 25130 41201 25190 41589
rect 26722 41538 26738 42962
rect 26802 42280 26818 42962
rect 30120 42911 30180 43299
rect 31712 43248 31728 44672
rect 31792 43990 31808 44672
rect 35110 44621 35170 45009
rect 36702 44958 36718 46382
rect 36782 45700 36798 46382
rect 40100 46331 40160 46719
rect 41692 46668 41708 48092
rect 41772 47410 41788 48092
rect 45090 48041 45150 48429
rect 46682 48378 46698 49802
rect 46762 49120 46778 49802
rect 50080 49751 50140 50139
rect 51672 50088 51688 51512
rect 51752 50830 51768 51512
rect 55070 51461 55130 51849
rect 56662 51798 56678 53222
rect 56742 52540 56758 53222
rect 60060 53171 60120 53559
rect 61652 53508 61668 54932
rect 61732 54250 61748 54932
rect 65050 54881 65110 55269
rect 66642 55218 66658 56642
rect 66722 55960 66738 56642
rect 70040 56591 70100 56979
rect 71632 56928 71648 58352
rect 71712 57670 71728 58352
rect 75030 58301 75090 58689
rect 76622 58638 76638 60062
rect 76702 59380 76718 60062
rect 78090 59440 78230 59470
rect 78090 59380 78120 59440
rect 76702 59370 78120 59380
rect 78200 59370 78230 59440
rect 76702 59330 78230 59370
rect 76702 59320 78120 59330
rect 76702 58638 76718 59320
rect 78090 59260 78120 59320
rect 78200 59260 78230 59330
rect 78090 59220 78230 59260
rect 76622 58622 76718 58638
rect 76622 58352 76718 58368
rect 75029 58300 76351 58301
rect 73100 57730 73240 57760
rect 73100 57670 73130 57730
rect 71712 57660 73130 57670
rect 73210 57660 73240 57730
rect 71712 57620 73240 57660
rect 71712 57610 73130 57620
rect 71712 56928 71728 57610
rect 73100 57550 73130 57610
rect 73210 57550 73240 57620
rect 73100 57510 73240 57550
rect 75029 56980 75030 58300
rect 76350 56980 76351 58300
rect 75029 56979 76351 56980
rect 71632 56912 71728 56928
rect 71632 56642 71728 56658
rect 70039 56590 71361 56591
rect 68110 56020 68250 56050
rect 68110 55960 68140 56020
rect 66722 55950 68140 55960
rect 68220 55950 68250 56020
rect 66722 55910 68250 55950
rect 66722 55900 68140 55910
rect 66722 55218 66738 55900
rect 68110 55840 68140 55900
rect 68220 55840 68250 55910
rect 68110 55800 68250 55840
rect 70039 55270 70040 56590
rect 71360 55270 71361 56590
rect 70039 55269 71361 55270
rect 66642 55202 66738 55218
rect 66642 54932 66738 54948
rect 65049 54880 66371 54881
rect 63120 54310 63260 54340
rect 63120 54250 63150 54310
rect 61732 54240 63150 54250
rect 63230 54240 63260 54310
rect 61732 54200 63260 54240
rect 61732 54190 63150 54200
rect 61732 53508 61748 54190
rect 63120 54130 63150 54190
rect 63230 54130 63260 54200
rect 63120 54090 63260 54130
rect 65049 53560 65050 54880
rect 66370 53560 66371 54880
rect 65049 53559 66371 53560
rect 61652 53492 61748 53508
rect 61652 53222 61748 53238
rect 60059 53170 61381 53171
rect 58130 52600 58270 52630
rect 58130 52540 58160 52600
rect 56742 52530 58160 52540
rect 58240 52530 58270 52600
rect 56742 52490 58270 52530
rect 56742 52480 58160 52490
rect 56742 51798 56758 52480
rect 58130 52420 58160 52480
rect 58240 52420 58270 52490
rect 58130 52380 58270 52420
rect 60059 51850 60060 53170
rect 61380 51850 61381 53170
rect 60059 51849 61381 51850
rect 56662 51782 56758 51798
rect 56662 51512 56758 51528
rect 55069 51460 56391 51461
rect 53140 50890 53280 50920
rect 53140 50830 53170 50890
rect 51752 50820 53170 50830
rect 53250 50820 53280 50890
rect 51752 50780 53280 50820
rect 51752 50770 53170 50780
rect 51752 50088 51768 50770
rect 53140 50710 53170 50770
rect 53250 50710 53280 50780
rect 53140 50670 53280 50710
rect 55069 50140 55070 51460
rect 56390 50140 56391 51460
rect 55069 50139 56391 50140
rect 51672 50072 51768 50088
rect 51672 49802 51768 49818
rect 50079 49750 51401 49751
rect 48150 49180 48290 49210
rect 48150 49120 48180 49180
rect 46762 49110 48180 49120
rect 48260 49110 48290 49180
rect 46762 49070 48290 49110
rect 46762 49060 48180 49070
rect 46762 48378 46778 49060
rect 48150 49000 48180 49060
rect 48260 49000 48290 49070
rect 48980 49060 49670 49120
rect 48150 48960 48290 49000
rect 50079 48430 50080 49750
rect 51400 48430 51401 49750
rect 50079 48429 51401 48430
rect 46682 48362 46778 48378
rect 46682 48092 46778 48108
rect 45089 48040 46411 48041
rect 43160 47470 43300 47500
rect 43160 47410 43190 47470
rect 41772 47400 43190 47410
rect 43270 47400 43300 47470
rect 41772 47360 43300 47400
rect 41772 47350 43190 47360
rect 41772 46668 41788 47350
rect 43160 47290 43190 47350
rect 43270 47290 43300 47360
rect 43160 47250 43300 47290
rect 45089 46720 45090 48040
rect 46410 46720 46411 48040
rect 45089 46719 46411 46720
rect 41692 46652 41788 46668
rect 41692 46382 41788 46398
rect 40099 46330 41421 46331
rect 38170 45760 38310 45790
rect 38170 45700 38200 45760
rect 36782 45690 38200 45700
rect 38280 45690 38310 45760
rect 36782 45650 38310 45690
rect 36782 45640 38200 45650
rect 36782 44958 36798 45640
rect 38170 45580 38200 45640
rect 38280 45580 38310 45650
rect 38170 45540 38310 45580
rect 40099 45010 40100 46330
rect 41420 45010 41421 46330
rect 40099 45009 41421 45010
rect 36702 44942 36798 44958
rect 36702 44672 36798 44688
rect 35109 44620 36431 44621
rect 33180 44050 33320 44080
rect 33180 43990 33210 44050
rect 31792 43980 33210 43990
rect 33290 43980 33320 44050
rect 31792 43940 33320 43980
rect 31792 43930 33210 43940
rect 31792 43248 31808 43930
rect 33180 43870 33210 43930
rect 33290 43870 33320 43940
rect 34010 43930 34700 43990
rect 33180 43830 33320 43870
rect 35109 43300 35110 44620
rect 36430 43300 36431 44620
rect 35109 43299 36431 43300
rect 31712 43232 31808 43248
rect 31712 42962 31808 42978
rect 30119 42910 31441 42911
rect 28190 42340 28330 42370
rect 28190 42280 28220 42340
rect 26802 42270 28220 42280
rect 28300 42270 28330 42340
rect 26802 42230 28330 42270
rect 26802 42220 28220 42230
rect 26802 41538 26818 42220
rect 28190 42160 28220 42220
rect 28300 42160 28330 42230
rect 28190 42120 28330 42160
rect 30119 41590 30120 42910
rect 31440 41590 31441 42910
rect 30119 41589 31441 41590
rect 26722 41522 26818 41538
rect 26722 41252 26818 41268
rect 25129 41200 26451 41201
rect 23200 40630 23340 40660
rect 23200 40570 23230 40630
rect 21812 40560 23230 40570
rect 23310 40560 23340 40630
rect 21812 40520 23340 40560
rect 21812 40510 23230 40520
rect 21812 39828 21828 40510
rect 23200 40450 23230 40510
rect 23310 40450 23340 40520
rect 23200 40410 23340 40450
rect 25129 39880 25130 41200
rect 26450 39880 26451 41200
rect 25129 39879 26451 39880
rect 21732 39812 21828 39828
rect 25130 39690 25190 39879
rect 26722 39828 26738 41252
rect 26802 40570 26818 41252
rect 30120 41201 30180 41589
rect 31712 41538 31728 42962
rect 31792 42280 31808 42962
rect 35110 42911 35170 43299
rect 36702 43248 36718 44672
rect 36782 43990 36798 44672
rect 40100 44621 40160 45009
rect 41692 44958 41708 46382
rect 41772 45700 41788 46382
rect 45090 46331 45150 46719
rect 46682 46668 46698 48092
rect 46762 47410 46778 48092
rect 50080 48041 50140 48429
rect 51672 48378 51688 49802
rect 51752 49120 51768 49802
rect 55070 49751 55130 50139
rect 56662 50088 56678 51512
rect 56742 50830 56758 51512
rect 60060 51461 60120 51849
rect 61652 51798 61668 53222
rect 61732 52540 61748 53222
rect 65050 53171 65110 53559
rect 66642 53508 66658 54932
rect 66722 54250 66738 54932
rect 70040 54881 70100 55269
rect 71632 55218 71648 56642
rect 71712 55960 71728 56642
rect 75030 56591 75090 56979
rect 76622 56928 76638 58352
rect 76702 57670 76718 58352
rect 78090 57730 78230 57760
rect 78090 57670 78120 57730
rect 76702 57660 78120 57670
rect 78200 57660 78230 57730
rect 76702 57620 78230 57660
rect 76702 57610 78120 57620
rect 76702 56928 76718 57610
rect 78090 57550 78120 57610
rect 78200 57550 78230 57620
rect 78090 57510 78230 57550
rect 76622 56912 76718 56928
rect 76622 56642 76718 56658
rect 75029 56590 76351 56591
rect 73100 56020 73240 56050
rect 73100 55960 73130 56020
rect 71712 55950 73130 55960
rect 73210 55950 73240 56020
rect 71712 55910 73240 55950
rect 71712 55900 73130 55910
rect 71712 55218 71728 55900
rect 73100 55840 73130 55900
rect 73210 55840 73240 55910
rect 73100 55800 73240 55840
rect 75029 55270 75030 56590
rect 76350 55270 76351 56590
rect 75029 55269 76351 55270
rect 71632 55202 71728 55218
rect 71632 54932 71728 54948
rect 70039 54880 71361 54881
rect 68110 54310 68250 54340
rect 68110 54250 68140 54310
rect 66722 54240 68140 54250
rect 68220 54240 68250 54310
rect 66722 54200 68250 54240
rect 66722 54190 68140 54200
rect 66722 53508 66738 54190
rect 68110 54130 68140 54190
rect 68220 54130 68250 54200
rect 68110 54090 68250 54130
rect 70039 53560 70040 54880
rect 71360 53560 71361 54880
rect 70039 53559 71361 53560
rect 66642 53492 66738 53508
rect 66642 53222 66738 53238
rect 65049 53170 66371 53171
rect 63120 52600 63260 52630
rect 63120 52540 63150 52600
rect 61732 52530 63150 52540
rect 63230 52530 63260 52600
rect 61732 52490 63260 52530
rect 61732 52480 63150 52490
rect 61732 51798 61748 52480
rect 63120 52420 63150 52480
rect 63230 52420 63260 52490
rect 63120 52380 63260 52420
rect 65049 51850 65050 53170
rect 66370 51850 66371 53170
rect 65049 51849 66371 51850
rect 61652 51782 61748 51798
rect 61652 51512 61748 51528
rect 60059 51460 61381 51461
rect 58130 50890 58270 50920
rect 58130 50830 58160 50890
rect 56742 50820 58160 50830
rect 58240 50820 58270 50890
rect 56742 50780 58270 50820
rect 56742 50770 58160 50780
rect 56742 50088 56758 50770
rect 58130 50710 58160 50770
rect 58240 50710 58270 50780
rect 58130 50670 58270 50710
rect 60059 50140 60060 51460
rect 61380 50140 61381 51460
rect 60059 50139 61381 50140
rect 56662 50072 56758 50088
rect 56662 49802 56758 49818
rect 55069 49750 56391 49751
rect 53140 49180 53280 49210
rect 53140 49120 53170 49180
rect 51752 49110 53170 49120
rect 53250 49110 53280 49180
rect 51752 49070 53280 49110
rect 51752 49060 53170 49070
rect 51752 48378 51768 49060
rect 53140 49000 53170 49060
rect 53250 49000 53280 49070
rect 53140 48960 53280 49000
rect 55069 48430 55070 49750
rect 56390 48430 56391 49750
rect 55069 48429 56391 48430
rect 51672 48362 51768 48378
rect 51672 48092 51768 48108
rect 50079 48040 51401 48041
rect 48150 47470 48290 47500
rect 48150 47410 48180 47470
rect 46762 47400 48180 47410
rect 48260 47400 48290 47470
rect 46762 47360 48290 47400
rect 46762 47350 48180 47360
rect 46762 46668 46778 47350
rect 48150 47290 48180 47350
rect 48260 47290 48290 47360
rect 48980 47350 49670 47410
rect 48150 47250 48290 47290
rect 50079 46720 50080 48040
rect 51400 46720 51401 48040
rect 50079 46719 51401 46720
rect 46682 46652 46778 46668
rect 46682 46382 46778 46398
rect 45089 46330 46411 46331
rect 43160 45760 43300 45790
rect 43160 45700 43190 45760
rect 41772 45690 43190 45700
rect 43270 45690 43300 45760
rect 41772 45650 43300 45690
rect 41772 45640 43190 45650
rect 41772 44958 41788 45640
rect 43160 45580 43190 45640
rect 43270 45580 43300 45650
rect 43160 45540 43300 45580
rect 45089 45010 45090 46330
rect 46410 45010 46411 46330
rect 45089 45009 46411 45010
rect 41692 44942 41788 44958
rect 41692 44672 41788 44688
rect 40099 44620 41421 44621
rect 38170 44050 38310 44080
rect 38170 43990 38200 44050
rect 36782 43980 38200 43990
rect 38280 43980 38310 44050
rect 36782 43940 38310 43980
rect 36782 43930 38200 43940
rect 36782 43248 36798 43930
rect 38170 43870 38200 43930
rect 38280 43870 38310 43940
rect 38170 43830 38310 43870
rect 40099 43300 40100 44620
rect 41420 43300 41421 44620
rect 40099 43299 41421 43300
rect 36702 43232 36798 43248
rect 36702 42962 36798 42978
rect 35109 42910 36431 42911
rect 33180 42340 33320 42370
rect 33180 42280 33210 42340
rect 31792 42270 33210 42280
rect 33290 42270 33320 42340
rect 31792 42230 33320 42270
rect 31792 42220 33210 42230
rect 31792 41538 31808 42220
rect 33180 42160 33210 42220
rect 33290 42160 33320 42230
rect 34010 42220 34700 42280
rect 33180 42120 33320 42160
rect 35109 41590 35110 42910
rect 36430 41590 36431 42910
rect 35109 41589 36431 41590
rect 31712 41522 31808 41538
rect 31712 41252 31808 41268
rect 30119 41200 31441 41201
rect 28190 40630 28330 40660
rect 28190 40570 28220 40630
rect 26802 40560 28220 40570
rect 28300 40560 28330 40630
rect 26802 40520 28330 40560
rect 26802 40510 28220 40520
rect 26802 39828 26818 40510
rect 28190 40450 28220 40510
rect 28300 40450 28330 40520
rect 28190 40410 28330 40450
rect 30119 39880 30120 41200
rect 31440 39880 31441 41200
rect 30119 39879 31441 39880
rect 26722 39812 26818 39828
rect 30120 39690 30180 39879
rect 31712 39828 31728 41252
rect 31792 40570 31808 41252
rect 35110 41201 35170 41589
rect 36702 41538 36718 42962
rect 36782 42280 36798 42962
rect 40100 42911 40160 43299
rect 41692 43248 41708 44672
rect 41772 43990 41788 44672
rect 45090 44621 45150 45009
rect 46682 44958 46698 46382
rect 46762 45700 46778 46382
rect 50080 46331 50140 46719
rect 51672 46668 51688 48092
rect 51752 47410 51768 48092
rect 55070 48041 55130 48429
rect 56662 48378 56678 49802
rect 56742 49120 56758 49802
rect 60060 49751 60120 50139
rect 61652 50088 61668 51512
rect 61732 50830 61748 51512
rect 65050 51461 65110 51849
rect 66642 51798 66658 53222
rect 66722 52540 66738 53222
rect 70040 53171 70100 53559
rect 71632 53508 71648 54932
rect 71712 54250 71728 54932
rect 75030 54881 75090 55269
rect 76622 55218 76638 56642
rect 76702 55960 76718 56642
rect 78090 56020 78230 56050
rect 78090 55960 78120 56020
rect 76702 55950 78120 55960
rect 78200 55950 78230 56020
rect 76702 55910 78230 55950
rect 76702 55900 78120 55910
rect 76702 55218 76718 55900
rect 78090 55840 78120 55900
rect 78200 55840 78230 55910
rect 78090 55800 78230 55840
rect 76622 55202 76718 55218
rect 76622 54932 76718 54948
rect 75029 54880 76351 54881
rect 73100 54310 73240 54340
rect 73100 54250 73130 54310
rect 71712 54240 73130 54250
rect 73210 54240 73240 54310
rect 71712 54200 73240 54240
rect 71712 54190 73130 54200
rect 71712 53508 71728 54190
rect 73100 54130 73130 54190
rect 73210 54130 73240 54200
rect 73100 54090 73240 54130
rect 75029 53560 75030 54880
rect 76350 53560 76351 54880
rect 75029 53559 76351 53560
rect 71632 53492 71728 53508
rect 71632 53222 71728 53238
rect 70039 53170 71361 53171
rect 68110 52600 68250 52630
rect 68110 52540 68140 52600
rect 66722 52530 68140 52540
rect 68220 52530 68250 52600
rect 66722 52490 68250 52530
rect 66722 52480 68140 52490
rect 66722 51798 66738 52480
rect 68110 52420 68140 52480
rect 68220 52420 68250 52490
rect 68110 52380 68250 52420
rect 70039 51850 70040 53170
rect 71360 51850 71361 53170
rect 70039 51849 71361 51850
rect 66642 51782 66738 51798
rect 66642 51512 66738 51528
rect 65049 51460 66371 51461
rect 63120 50890 63260 50920
rect 63120 50830 63150 50890
rect 61732 50820 63150 50830
rect 63230 50820 63260 50890
rect 61732 50780 63260 50820
rect 61732 50770 63150 50780
rect 61732 50088 61748 50770
rect 63120 50710 63150 50770
rect 63230 50710 63260 50780
rect 63120 50670 63260 50710
rect 65049 50140 65050 51460
rect 66370 50140 66371 51460
rect 65049 50139 66371 50140
rect 61652 50072 61748 50088
rect 61652 49802 61748 49818
rect 60059 49750 61381 49751
rect 58130 49180 58270 49210
rect 58130 49120 58160 49180
rect 56742 49110 58160 49120
rect 58240 49110 58270 49180
rect 56742 49070 58270 49110
rect 56742 49060 58160 49070
rect 56742 48378 56758 49060
rect 58130 49000 58160 49060
rect 58240 49000 58270 49070
rect 58130 48960 58270 49000
rect 60059 48430 60060 49750
rect 61380 48430 61381 49750
rect 60059 48429 61381 48430
rect 56662 48362 56758 48378
rect 56662 48092 56758 48108
rect 55069 48040 56391 48041
rect 53140 47470 53280 47500
rect 53140 47410 53170 47470
rect 51752 47400 53170 47410
rect 53250 47400 53280 47470
rect 51752 47360 53280 47400
rect 51752 47350 53170 47360
rect 51752 46668 51768 47350
rect 53140 47290 53170 47350
rect 53250 47290 53280 47360
rect 53140 47250 53280 47290
rect 55069 46720 55070 48040
rect 56390 46720 56391 48040
rect 55069 46719 56391 46720
rect 51672 46652 51768 46668
rect 51672 46382 51768 46398
rect 50079 46330 51401 46331
rect 48150 45760 48290 45790
rect 48150 45700 48180 45760
rect 46762 45690 48180 45700
rect 48260 45690 48290 45760
rect 46762 45650 48290 45690
rect 46762 45640 48180 45650
rect 46762 44958 46778 45640
rect 48150 45580 48180 45640
rect 48260 45580 48290 45650
rect 48980 45640 49670 45700
rect 48150 45540 48290 45580
rect 50079 45010 50080 46330
rect 51400 45010 51401 46330
rect 50079 45009 51401 45010
rect 46682 44942 46778 44958
rect 46682 44672 46778 44688
rect 45089 44620 46411 44621
rect 43160 44050 43300 44080
rect 43160 43990 43190 44050
rect 41772 43980 43190 43990
rect 43270 43980 43300 44050
rect 41772 43940 43300 43980
rect 41772 43930 43190 43940
rect 41772 43248 41788 43930
rect 43160 43870 43190 43930
rect 43270 43870 43300 43940
rect 43160 43830 43300 43870
rect 45089 43300 45090 44620
rect 46410 43300 46411 44620
rect 45089 43299 46411 43300
rect 41692 43232 41788 43248
rect 41692 42962 41788 42978
rect 40099 42910 41421 42911
rect 38170 42340 38310 42370
rect 38170 42280 38200 42340
rect 36782 42270 38200 42280
rect 38280 42270 38310 42340
rect 36782 42230 38310 42270
rect 36782 42220 38200 42230
rect 36782 41538 36798 42220
rect 38170 42160 38200 42220
rect 38280 42160 38310 42230
rect 38170 42120 38310 42160
rect 40099 41590 40100 42910
rect 41420 41590 41421 42910
rect 40099 41589 41421 41590
rect 36702 41522 36798 41538
rect 36702 41252 36798 41268
rect 35109 41200 36431 41201
rect 33180 40630 33320 40660
rect 33180 40570 33210 40630
rect 31792 40560 33210 40570
rect 33290 40560 33320 40630
rect 31792 40520 33320 40560
rect 31792 40510 33210 40520
rect 31792 39828 31808 40510
rect 33180 40450 33210 40510
rect 33290 40450 33320 40520
rect 34010 40510 34700 40570
rect 33180 40410 33320 40450
rect 35109 39880 35110 41200
rect 36430 39880 36431 41200
rect 35109 39879 36431 39880
rect 31712 39812 31808 39828
rect 35110 39690 35170 39879
rect 36702 39828 36718 41252
rect 36782 40570 36798 41252
rect 40100 41201 40160 41589
rect 41692 41538 41708 42962
rect 41772 42280 41788 42962
rect 45090 42911 45150 43299
rect 46682 43248 46698 44672
rect 46762 43990 46778 44672
rect 50080 44621 50140 45009
rect 51672 44958 51688 46382
rect 51752 45700 51768 46382
rect 55070 46331 55130 46719
rect 56662 46668 56678 48092
rect 56742 47410 56758 48092
rect 60060 48041 60120 48429
rect 61652 48378 61668 49802
rect 61732 49120 61748 49802
rect 65050 49751 65110 50139
rect 66642 50088 66658 51512
rect 66722 50830 66738 51512
rect 70040 51461 70100 51849
rect 71632 51798 71648 53222
rect 71712 52540 71728 53222
rect 75030 53171 75090 53559
rect 76622 53508 76638 54932
rect 76702 54250 76718 54932
rect 78090 54310 78230 54340
rect 78090 54250 78120 54310
rect 76702 54240 78120 54250
rect 78200 54240 78230 54310
rect 76702 54200 78230 54240
rect 76702 54190 78120 54200
rect 76702 53508 76718 54190
rect 78090 54130 78120 54190
rect 78200 54130 78230 54200
rect 78090 54090 78230 54130
rect 76622 53492 76718 53508
rect 76622 53222 76718 53238
rect 75029 53170 76351 53171
rect 73100 52600 73240 52630
rect 73100 52540 73130 52600
rect 71712 52530 73130 52540
rect 73210 52530 73240 52600
rect 71712 52490 73240 52530
rect 71712 52480 73130 52490
rect 71712 51798 71728 52480
rect 73100 52420 73130 52480
rect 73210 52420 73240 52490
rect 73100 52380 73240 52420
rect 75029 51850 75030 53170
rect 76350 51850 76351 53170
rect 75029 51849 76351 51850
rect 71632 51782 71728 51798
rect 71632 51512 71728 51528
rect 70039 51460 71361 51461
rect 68110 50890 68250 50920
rect 68110 50830 68140 50890
rect 66722 50820 68140 50830
rect 68220 50820 68250 50890
rect 66722 50780 68250 50820
rect 66722 50770 68140 50780
rect 66722 50088 66738 50770
rect 68110 50710 68140 50770
rect 68220 50710 68250 50780
rect 68110 50670 68250 50710
rect 70039 50140 70040 51460
rect 71360 50140 71361 51460
rect 70039 50139 71361 50140
rect 66642 50072 66738 50088
rect 66642 49802 66738 49818
rect 65049 49750 66371 49751
rect 63120 49180 63260 49210
rect 63120 49120 63150 49180
rect 61732 49110 63150 49120
rect 63230 49110 63260 49180
rect 61732 49070 63260 49110
rect 61732 49060 63150 49070
rect 61732 48378 61748 49060
rect 63120 49000 63150 49060
rect 63230 49000 63260 49070
rect 63120 48960 63260 49000
rect 65049 48430 65050 49750
rect 66370 48430 66371 49750
rect 65049 48429 66371 48430
rect 61652 48362 61748 48378
rect 61652 48092 61748 48108
rect 60059 48040 61381 48041
rect 58130 47470 58270 47500
rect 58130 47410 58160 47470
rect 56742 47400 58160 47410
rect 58240 47400 58270 47470
rect 56742 47360 58270 47400
rect 56742 47350 58160 47360
rect 56742 46668 56758 47350
rect 58130 47290 58160 47350
rect 58240 47290 58270 47360
rect 58130 47250 58270 47290
rect 60059 46720 60060 48040
rect 61380 46720 61381 48040
rect 60059 46719 61381 46720
rect 56662 46652 56758 46668
rect 56662 46382 56758 46398
rect 55069 46330 56391 46331
rect 53140 45760 53280 45790
rect 53140 45700 53170 45760
rect 51752 45690 53170 45700
rect 53250 45690 53280 45760
rect 51752 45650 53280 45690
rect 51752 45640 53170 45650
rect 51752 44958 51768 45640
rect 53140 45580 53170 45640
rect 53250 45580 53280 45650
rect 53140 45540 53280 45580
rect 55069 45010 55070 46330
rect 56390 45010 56391 46330
rect 55069 45009 56391 45010
rect 51672 44942 51768 44958
rect 51672 44672 51768 44688
rect 50079 44620 51401 44621
rect 48150 44050 48290 44080
rect 48150 43990 48180 44050
rect 46762 43980 48180 43990
rect 48260 43980 48290 44050
rect 46762 43940 48290 43980
rect 46762 43930 48180 43940
rect 46762 43248 46778 43930
rect 48150 43870 48180 43930
rect 48260 43870 48290 43940
rect 48980 43930 49670 43990
rect 48150 43830 48290 43870
rect 50079 43300 50080 44620
rect 51400 43300 51401 44620
rect 50079 43299 51401 43300
rect 46682 43232 46778 43248
rect 46682 42962 46778 42978
rect 45089 42910 46411 42911
rect 43160 42340 43300 42370
rect 43160 42280 43190 42340
rect 41772 42270 43190 42280
rect 43270 42270 43300 42340
rect 41772 42230 43300 42270
rect 41772 42220 43190 42230
rect 41772 41538 41788 42220
rect 43160 42160 43190 42220
rect 43270 42160 43300 42230
rect 43160 42120 43300 42160
rect 45089 41590 45090 42910
rect 46410 41590 46411 42910
rect 45089 41589 46411 41590
rect 41692 41522 41788 41538
rect 41692 41252 41788 41268
rect 40099 41200 41421 41201
rect 38170 40630 38310 40660
rect 38170 40570 38200 40630
rect 36782 40560 38200 40570
rect 38280 40560 38310 40630
rect 36782 40520 38310 40560
rect 36782 40510 38200 40520
rect 36782 39828 36798 40510
rect 38170 40450 38200 40510
rect 38280 40450 38310 40520
rect 38170 40410 38310 40450
rect 40099 39880 40100 41200
rect 41420 39880 41421 41200
rect 40099 39879 41421 39880
rect 36702 39812 36798 39828
rect 40100 39690 40160 39879
rect 41692 39828 41708 41252
rect 41772 40570 41788 41252
rect 45090 41201 45150 41589
rect 46682 41538 46698 42962
rect 46762 42280 46778 42962
rect 50080 42911 50140 43299
rect 51672 43248 51688 44672
rect 51752 43990 51768 44672
rect 55070 44621 55130 45009
rect 56662 44958 56678 46382
rect 56742 45700 56758 46382
rect 60060 46331 60120 46719
rect 61652 46668 61668 48092
rect 61732 47410 61748 48092
rect 65050 48041 65110 48429
rect 66642 48378 66658 49802
rect 66722 49120 66738 49802
rect 70040 49751 70100 50139
rect 71632 50088 71648 51512
rect 71712 50830 71728 51512
rect 75030 51461 75090 51849
rect 76622 51798 76638 53222
rect 76702 52540 76718 53222
rect 78090 52600 78230 52630
rect 78090 52540 78120 52600
rect 76702 52530 78120 52540
rect 78200 52530 78230 52600
rect 76702 52490 78230 52530
rect 76702 52480 78120 52490
rect 76702 51798 76718 52480
rect 78090 52420 78120 52480
rect 78200 52420 78230 52490
rect 78090 52380 78230 52420
rect 76622 51782 76718 51798
rect 76622 51512 76718 51528
rect 75029 51460 76351 51461
rect 73100 50890 73240 50920
rect 73100 50830 73130 50890
rect 71712 50820 73130 50830
rect 73210 50820 73240 50890
rect 71712 50780 73240 50820
rect 71712 50770 73130 50780
rect 71712 50088 71728 50770
rect 73100 50710 73130 50770
rect 73210 50710 73240 50780
rect 73100 50670 73240 50710
rect 75029 50140 75030 51460
rect 76350 50140 76351 51460
rect 75029 50139 76351 50140
rect 71632 50072 71728 50088
rect 71632 49802 71728 49818
rect 70039 49750 71361 49751
rect 68110 49180 68250 49210
rect 68110 49120 68140 49180
rect 66722 49110 68140 49120
rect 68220 49110 68250 49180
rect 66722 49070 68250 49110
rect 66722 49060 68140 49070
rect 66722 48378 66738 49060
rect 68110 49000 68140 49060
rect 68220 49000 68250 49070
rect 68110 48960 68250 49000
rect 70039 48430 70040 49750
rect 71360 48430 71361 49750
rect 70039 48429 71361 48430
rect 66642 48362 66738 48378
rect 66642 48092 66738 48108
rect 65049 48040 66371 48041
rect 63120 47470 63260 47500
rect 63120 47410 63150 47470
rect 61732 47400 63150 47410
rect 63230 47400 63260 47470
rect 61732 47360 63260 47400
rect 61732 47350 63150 47360
rect 61732 46668 61748 47350
rect 63120 47290 63150 47350
rect 63230 47290 63260 47360
rect 63120 47250 63260 47290
rect 65049 46720 65050 48040
rect 66370 46720 66371 48040
rect 65049 46719 66371 46720
rect 61652 46652 61748 46668
rect 61652 46382 61748 46398
rect 60059 46330 61381 46331
rect 58130 45760 58270 45790
rect 58130 45700 58160 45760
rect 56742 45690 58160 45700
rect 58240 45690 58270 45760
rect 56742 45650 58270 45690
rect 56742 45640 58160 45650
rect 56742 44958 56758 45640
rect 58130 45580 58160 45640
rect 58240 45580 58270 45650
rect 58130 45540 58270 45580
rect 60059 45010 60060 46330
rect 61380 45010 61381 46330
rect 60059 45009 61381 45010
rect 56662 44942 56758 44958
rect 56662 44672 56758 44688
rect 55069 44620 56391 44621
rect 53140 44050 53280 44080
rect 53140 43990 53170 44050
rect 51752 43980 53170 43990
rect 53250 43980 53280 44050
rect 51752 43940 53280 43980
rect 51752 43930 53170 43940
rect 51752 43248 51768 43930
rect 53140 43870 53170 43930
rect 53250 43870 53280 43940
rect 53140 43830 53280 43870
rect 55069 43300 55070 44620
rect 56390 43300 56391 44620
rect 55069 43299 56391 43300
rect 51672 43232 51768 43248
rect 51672 42962 51768 42978
rect 50079 42910 51401 42911
rect 48150 42340 48290 42370
rect 48150 42280 48180 42340
rect 46762 42270 48180 42280
rect 48260 42270 48290 42340
rect 46762 42230 48290 42270
rect 46762 42220 48180 42230
rect 46762 41538 46778 42220
rect 48150 42160 48180 42220
rect 48260 42160 48290 42230
rect 48980 42220 49670 42280
rect 48150 42120 48290 42160
rect 50079 41590 50080 42910
rect 51400 41590 51401 42910
rect 50079 41589 51401 41590
rect 46682 41522 46778 41538
rect 46682 41252 46778 41268
rect 45089 41200 46411 41201
rect 43160 40630 43300 40660
rect 43160 40570 43190 40630
rect 41772 40560 43190 40570
rect 43270 40560 43300 40630
rect 41772 40520 43300 40560
rect 41772 40510 43190 40520
rect 41772 39828 41788 40510
rect 43160 40450 43190 40510
rect 43270 40450 43300 40520
rect 43160 40410 43300 40450
rect 45089 39880 45090 41200
rect 46410 39880 46411 41200
rect 45089 39879 46411 39880
rect 41692 39812 41788 39828
rect 45090 39690 45150 39879
rect 46682 39828 46698 41252
rect 46762 40570 46778 41252
rect 50080 41201 50140 41589
rect 51672 41538 51688 42962
rect 51752 42280 51768 42962
rect 55070 42911 55130 43299
rect 56662 43248 56678 44672
rect 56742 43990 56758 44672
rect 60060 44621 60120 45009
rect 61652 44958 61668 46382
rect 61732 45700 61748 46382
rect 65050 46331 65110 46719
rect 66642 46668 66658 48092
rect 66722 47410 66738 48092
rect 70040 48041 70100 48429
rect 71632 48378 71648 49802
rect 71712 49120 71728 49802
rect 75030 49751 75090 50139
rect 76622 50088 76638 51512
rect 76702 50830 76718 51512
rect 78090 50890 78230 50920
rect 78090 50830 78120 50890
rect 76702 50820 78120 50830
rect 78200 50820 78230 50890
rect 76702 50780 78230 50820
rect 76702 50770 78120 50780
rect 76702 50088 76718 50770
rect 78090 50710 78120 50770
rect 78200 50710 78230 50780
rect 78090 50670 78230 50710
rect 76622 50072 76718 50088
rect 76622 49802 76718 49818
rect 75029 49750 76351 49751
rect 73100 49180 73240 49210
rect 73100 49120 73130 49180
rect 71712 49110 73130 49120
rect 73210 49110 73240 49180
rect 71712 49070 73240 49110
rect 71712 49060 73130 49070
rect 71712 48378 71728 49060
rect 73100 49000 73130 49060
rect 73210 49000 73240 49070
rect 73100 48960 73240 49000
rect 75029 48430 75030 49750
rect 76350 48430 76351 49750
rect 75029 48429 76351 48430
rect 71632 48362 71728 48378
rect 71632 48092 71728 48108
rect 70039 48040 71361 48041
rect 68110 47470 68250 47500
rect 68110 47410 68140 47470
rect 66722 47400 68140 47410
rect 68220 47400 68250 47470
rect 66722 47360 68250 47400
rect 66722 47350 68140 47360
rect 66722 46668 66738 47350
rect 68110 47290 68140 47350
rect 68220 47290 68250 47360
rect 68110 47250 68250 47290
rect 70039 46720 70040 48040
rect 71360 46720 71361 48040
rect 70039 46719 71361 46720
rect 66642 46652 66738 46668
rect 66642 46382 66738 46398
rect 65049 46330 66371 46331
rect 63120 45760 63260 45790
rect 63120 45700 63150 45760
rect 61732 45690 63150 45700
rect 63230 45690 63260 45760
rect 61732 45650 63260 45690
rect 61732 45640 63150 45650
rect 61732 44958 61748 45640
rect 63120 45580 63150 45640
rect 63230 45580 63260 45650
rect 63120 45540 63260 45580
rect 65049 45010 65050 46330
rect 66370 45010 66371 46330
rect 65049 45009 66371 45010
rect 61652 44942 61748 44958
rect 61652 44672 61748 44688
rect 60059 44620 61381 44621
rect 58130 44050 58270 44080
rect 58130 43990 58160 44050
rect 56742 43980 58160 43990
rect 58240 43980 58270 44050
rect 56742 43940 58270 43980
rect 56742 43930 58160 43940
rect 56742 43248 56758 43930
rect 58130 43870 58160 43930
rect 58240 43870 58270 43940
rect 58130 43830 58270 43870
rect 60059 43300 60060 44620
rect 61380 43300 61381 44620
rect 60059 43299 61381 43300
rect 56662 43232 56758 43248
rect 56662 42962 56758 42978
rect 55069 42910 56391 42911
rect 53140 42340 53280 42370
rect 53140 42280 53170 42340
rect 51752 42270 53170 42280
rect 53250 42270 53280 42340
rect 51752 42230 53280 42270
rect 51752 42220 53170 42230
rect 51752 41538 51768 42220
rect 53140 42160 53170 42220
rect 53250 42160 53280 42230
rect 53140 42120 53280 42160
rect 55069 41590 55070 42910
rect 56390 41590 56391 42910
rect 55069 41589 56391 41590
rect 51672 41522 51768 41538
rect 51672 41252 51768 41268
rect 50079 41200 51401 41201
rect 48150 40630 48290 40660
rect 48150 40570 48180 40630
rect 46762 40560 48180 40570
rect 48260 40560 48290 40630
rect 46762 40520 48290 40560
rect 46762 40510 48180 40520
rect 46762 39828 46778 40510
rect 48150 40450 48180 40510
rect 48260 40450 48290 40520
rect 48980 40510 49670 40570
rect 48150 40410 48290 40450
rect 50079 39880 50080 41200
rect 51400 39880 51401 41200
rect 50079 39879 51401 39880
rect 46682 39812 46778 39828
rect 50080 39690 50140 39879
rect 51672 39828 51688 41252
rect 51752 40570 51768 41252
rect 55070 41201 55130 41589
rect 56662 41538 56678 42962
rect 56742 42280 56758 42962
rect 60060 42911 60120 43299
rect 61652 43248 61668 44672
rect 61732 43990 61748 44672
rect 65050 44621 65110 45009
rect 66642 44958 66658 46382
rect 66722 45700 66738 46382
rect 70040 46331 70100 46719
rect 71632 46668 71648 48092
rect 71712 47410 71728 48092
rect 75030 48041 75090 48429
rect 76622 48378 76638 49802
rect 76702 49120 76718 49802
rect 78090 49180 78230 49210
rect 78090 49120 78120 49180
rect 76702 49110 78120 49120
rect 78200 49110 78230 49180
rect 76702 49070 78230 49110
rect 76702 49060 78120 49070
rect 76702 48378 76718 49060
rect 78090 49000 78120 49060
rect 78200 49000 78230 49070
rect 78090 48960 78230 49000
rect 76622 48362 76718 48378
rect 76622 48092 76718 48108
rect 75029 48040 76351 48041
rect 73100 47470 73240 47500
rect 73100 47410 73130 47470
rect 71712 47400 73130 47410
rect 73210 47400 73240 47470
rect 71712 47360 73240 47400
rect 71712 47350 73130 47360
rect 71712 46668 71728 47350
rect 73100 47290 73130 47350
rect 73210 47290 73240 47360
rect 73100 47250 73240 47290
rect 75029 46720 75030 48040
rect 76350 46720 76351 48040
rect 75029 46719 76351 46720
rect 71632 46652 71728 46668
rect 71632 46382 71728 46398
rect 70039 46330 71361 46331
rect 68110 45760 68250 45790
rect 68110 45700 68140 45760
rect 66722 45690 68140 45700
rect 68220 45690 68250 45760
rect 66722 45650 68250 45690
rect 66722 45640 68140 45650
rect 66722 44958 66738 45640
rect 68110 45580 68140 45640
rect 68220 45580 68250 45650
rect 68110 45540 68250 45580
rect 70039 45010 70040 46330
rect 71360 45010 71361 46330
rect 70039 45009 71361 45010
rect 66642 44942 66738 44958
rect 66642 44672 66738 44688
rect 65049 44620 66371 44621
rect 63120 44050 63260 44080
rect 63120 43990 63150 44050
rect 61732 43980 63150 43990
rect 63230 43980 63260 44050
rect 61732 43940 63260 43980
rect 61732 43930 63150 43940
rect 61732 43248 61748 43930
rect 63120 43870 63150 43930
rect 63230 43870 63260 43940
rect 63120 43830 63260 43870
rect 65049 43300 65050 44620
rect 66370 43300 66371 44620
rect 65049 43299 66371 43300
rect 61652 43232 61748 43248
rect 61652 42962 61748 42978
rect 60059 42910 61381 42911
rect 58130 42340 58270 42370
rect 58130 42280 58160 42340
rect 56742 42270 58160 42280
rect 58240 42270 58270 42340
rect 56742 42230 58270 42270
rect 56742 42220 58160 42230
rect 56742 41538 56758 42220
rect 58130 42160 58160 42220
rect 58240 42160 58270 42230
rect 58130 42120 58270 42160
rect 60059 41590 60060 42910
rect 61380 41590 61381 42910
rect 60059 41589 61381 41590
rect 56662 41522 56758 41538
rect 56662 41252 56758 41268
rect 55069 41200 56391 41201
rect 53140 40630 53280 40660
rect 53140 40570 53170 40630
rect 51752 40560 53170 40570
rect 53250 40560 53280 40630
rect 51752 40520 53280 40560
rect 51752 40510 53170 40520
rect 51752 39828 51768 40510
rect 53140 40450 53170 40510
rect 53250 40450 53280 40520
rect 53140 40410 53280 40450
rect 55069 39880 55070 41200
rect 56390 39880 56391 41200
rect 55069 39879 56391 39880
rect 51672 39812 51768 39828
rect 55070 39690 55130 39879
rect 56662 39828 56678 41252
rect 56742 40570 56758 41252
rect 60060 41201 60120 41589
rect 61652 41538 61668 42962
rect 61732 42280 61748 42962
rect 65050 42911 65110 43299
rect 66642 43248 66658 44672
rect 66722 43990 66738 44672
rect 70040 44621 70100 45009
rect 71632 44958 71648 46382
rect 71712 45700 71728 46382
rect 75030 46331 75090 46719
rect 76622 46668 76638 48092
rect 76702 47410 76718 48092
rect 78090 47470 78230 47500
rect 78090 47410 78120 47470
rect 76702 47400 78120 47410
rect 78200 47400 78230 47470
rect 76702 47360 78230 47400
rect 76702 47350 78120 47360
rect 76702 46668 76718 47350
rect 78090 47290 78120 47350
rect 78200 47290 78230 47360
rect 78090 47250 78230 47290
rect 76622 46652 76718 46668
rect 76622 46382 76718 46398
rect 75029 46330 76351 46331
rect 73100 45760 73240 45790
rect 73100 45700 73130 45760
rect 71712 45690 73130 45700
rect 73210 45690 73240 45760
rect 71712 45650 73240 45690
rect 71712 45640 73130 45650
rect 71712 44958 71728 45640
rect 73100 45580 73130 45640
rect 73210 45580 73240 45650
rect 73100 45540 73240 45580
rect 75029 45010 75030 46330
rect 76350 45010 76351 46330
rect 75029 45009 76351 45010
rect 71632 44942 71728 44958
rect 71632 44672 71728 44688
rect 70039 44620 71361 44621
rect 68110 44050 68250 44080
rect 68110 43990 68140 44050
rect 66722 43980 68140 43990
rect 68220 43980 68250 44050
rect 66722 43940 68250 43980
rect 66722 43930 68140 43940
rect 66722 43248 66738 43930
rect 68110 43870 68140 43930
rect 68220 43870 68250 43940
rect 68110 43830 68250 43870
rect 70039 43300 70040 44620
rect 71360 43300 71361 44620
rect 70039 43299 71361 43300
rect 66642 43232 66738 43248
rect 66642 42962 66738 42978
rect 65049 42910 66371 42911
rect 63120 42340 63260 42370
rect 63120 42280 63150 42340
rect 61732 42270 63150 42280
rect 63230 42270 63260 42340
rect 61732 42230 63260 42270
rect 61732 42220 63150 42230
rect 61732 41538 61748 42220
rect 63120 42160 63150 42220
rect 63230 42160 63260 42230
rect 63120 42120 63260 42160
rect 65049 41590 65050 42910
rect 66370 41590 66371 42910
rect 65049 41589 66371 41590
rect 61652 41522 61748 41538
rect 61652 41252 61748 41268
rect 60059 41200 61381 41201
rect 58130 40630 58270 40660
rect 58130 40570 58160 40630
rect 56742 40560 58160 40570
rect 58240 40560 58270 40630
rect 56742 40520 58270 40560
rect 56742 40510 58160 40520
rect 56742 39828 56758 40510
rect 58130 40450 58160 40510
rect 58240 40450 58270 40520
rect 58130 40410 58270 40450
rect 60059 39880 60060 41200
rect 61380 39880 61381 41200
rect 60059 39879 61381 39880
rect 56662 39812 56758 39828
rect 60060 39690 60120 39879
rect 61652 39828 61668 41252
rect 61732 40570 61748 41252
rect 65050 41201 65110 41589
rect 66642 41538 66658 42962
rect 66722 42280 66738 42962
rect 70040 42911 70100 43299
rect 71632 43248 71648 44672
rect 71712 43990 71728 44672
rect 75030 44621 75090 45009
rect 76622 44958 76638 46382
rect 76702 45700 76718 46382
rect 78090 45760 78230 45790
rect 78090 45700 78120 45760
rect 76702 45690 78120 45700
rect 78200 45690 78230 45760
rect 76702 45650 78230 45690
rect 76702 45640 78120 45650
rect 76702 44958 76718 45640
rect 78090 45580 78120 45640
rect 78200 45580 78230 45650
rect 78090 45540 78230 45580
rect 76622 44942 76718 44958
rect 76622 44672 76718 44688
rect 75029 44620 76351 44621
rect 73100 44050 73240 44080
rect 73100 43990 73130 44050
rect 71712 43980 73130 43990
rect 73210 43980 73240 44050
rect 71712 43940 73240 43980
rect 71712 43930 73130 43940
rect 71712 43248 71728 43930
rect 73100 43870 73130 43930
rect 73210 43870 73240 43940
rect 73100 43830 73240 43870
rect 75029 43300 75030 44620
rect 76350 43300 76351 44620
rect 75029 43299 76351 43300
rect 71632 43232 71728 43248
rect 71632 42962 71728 42978
rect 70039 42910 71361 42911
rect 68110 42340 68250 42370
rect 68110 42280 68140 42340
rect 66722 42270 68140 42280
rect 68220 42270 68250 42340
rect 66722 42230 68250 42270
rect 66722 42220 68140 42230
rect 66722 41538 66738 42220
rect 68110 42160 68140 42220
rect 68220 42160 68250 42230
rect 68110 42120 68250 42160
rect 70039 41590 70040 42910
rect 71360 41590 71361 42910
rect 70039 41589 71361 41590
rect 66642 41522 66738 41538
rect 66642 41252 66738 41268
rect 65049 41200 66371 41201
rect 63120 40630 63260 40660
rect 63120 40570 63150 40630
rect 61732 40560 63150 40570
rect 63230 40560 63260 40630
rect 61732 40520 63260 40560
rect 61732 40510 63150 40520
rect 61732 39828 61748 40510
rect 63120 40450 63150 40510
rect 63230 40450 63260 40520
rect 63120 40410 63260 40450
rect 65049 39880 65050 41200
rect 66370 39880 66371 41200
rect 65049 39879 66371 39880
rect 61652 39812 61748 39828
rect 65050 39690 65110 39879
rect 66642 39828 66658 41252
rect 66722 40570 66738 41252
rect 70040 41201 70100 41589
rect 71632 41538 71648 42962
rect 71712 42280 71728 42962
rect 75030 42911 75090 43299
rect 76622 43248 76638 44672
rect 76702 43990 76718 44672
rect 78090 44050 78230 44080
rect 78090 43990 78120 44050
rect 76702 43980 78120 43990
rect 78200 43980 78230 44050
rect 76702 43940 78230 43980
rect 76702 43930 78120 43940
rect 76702 43248 76718 43930
rect 78090 43870 78120 43930
rect 78200 43870 78230 43940
rect 78090 43830 78230 43870
rect 76622 43232 76718 43248
rect 76622 42962 76718 42978
rect 75029 42910 76351 42911
rect 73100 42340 73240 42370
rect 73100 42280 73130 42340
rect 71712 42270 73130 42280
rect 73210 42270 73240 42340
rect 71712 42230 73240 42270
rect 71712 42220 73130 42230
rect 71712 41538 71728 42220
rect 73100 42160 73130 42220
rect 73210 42160 73240 42230
rect 73100 42120 73240 42160
rect 75029 41590 75030 42910
rect 76350 41590 76351 42910
rect 75029 41589 76351 41590
rect 71632 41522 71728 41538
rect 71632 41252 71728 41268
rect 70039 41200 71361 41201
rect 68110 40630 68250 40660
rect 68110 40570 68140 40630
rect 66722 40560 68140 40570
rect 68220 40560 68250 40630
rect 66722 40520 68250 40560
rect 66722 40510 68140 40520
rect 66722 39828 66738 40510
rect 68110 40450 68140 40510
rect 68220 40450 68250 40520
rect 68110 40410 68250 40450
rect 70039 39880 70040 41200
rect 71360 39880 71361 41200
rect 70039 39879 71361 39880
rect 66642 39812 66738 39828
rect 70040 39690 70100 39879
rect 71632 39828 71648 41252
rect 71712 40570 71728 41252
rect 75030 41201 75090 41589
rect 76622 41538 76638 42962
rect 76702 42280 76718 42962
rect 78090 42340 78230 42370
rect 78090 42280 78120 42340
rect 76702 42270 78120 42280
rect 78200 42270 78230 42340
rect 76702 42230 78230 42270
rect 76702 42220 78120 42230
rect 76702 41538 76718 42220
rect 78090 42160 78120 42220
rect 78200 42160 78230 42230
rect 78090 42120 78230 42160
rect 76622 41522 76718 41538
rect 76622 41252 76718 41268
rect 75029 41200 76351 41201
rect 73100 40630 73240 40660
rect 73100 40570 73130 40630
rect 71712 40560 73130 40570
rect 73210 40560 73240 40630
rect 71712 40520 73240 40560
rect 71712 40510 73130 40520
rect 71712 39828 71728 40510
rect 73100 40450 73130 40510
rect 73210 40450 73240 40520
rect 73100 40410 73240 40450
rect 75029 39880 75030 41200
rect 76350 39880 76351 41200
rect 75029 39879 76351 39880
rect 71632 39812 71728 39828
rect 75030 39690 75090 39879
rect 76622 39828 76638 41252
rect 76702 40570 76718 41252
rect 78090 40630 78230 40660
rect 78090 40570 78120 40630
rect 76702 40560 78120 40570
rect 78200 40560 78230 40630
rect 76702 40520 78230 40560
rect 76702 40510 78120 40520
rect 76702 39828 76718 40510
rect 78090 40450 78120 40510
rect 78200 40450 78230 40520
rect 78090 40410 78230 40450
rect 76622 39812 76718 39828
rect 80 -60 140 0
rect 5070 -60 5130 0
rect 10060 -60 10120 0
rect 15050 -60 15110 0
rect 20040 -60 20100 0
rect 25030 -60 25090 0
rect 30020 -60 30080 0
rect 35010 -60 35070 0
rect 40000 -60 40060 0
rect 44990 -60 45050 0
rect 49980 -60 50040 0
rect 54970 -60 55030 0
rect 59960 -60 60020 0
rect 64950 -60 65010 0
rect 69940 -60 70000 0
rect 74930 -60 74990 0
rect 0 -120 79570 -60
use end  end_0 ~/dac_layout
timestamp 1729689530
transform 0 1 0 -1 0 27360
box 0 0 27360 4720
use end  end_1
timestamp 1729689530
transform 0 1 4990 -1 0 27360
box 0 0 27360 4720
use end  end_2
timestamp 1729689530
transform 0 1 69860 -1 0 27360
box 0 0 27360 4720
use end  end_3
timestamp 1729689530
transform 0 1 74850 -1 0 27360
box 0 0 27360 4720
use mid_2  mid_2_0 ~/dac_layout
timestamp 1729709358
transform 1 0 34930 0 1 13680
box 0 -13680 9800 13680
use mid_2to4_  mid_2to4__0 ~/dac_layout
timestamp 1729683266
transform 0 1 29940 -1 0 27360
box 0 0 27360 4720
use mid_2to4_  mid_2to4__1
timestamp 1729683266
transform 0 1 44910 -1 0 27360
box 0 0 27360 4720
use mid_4to8  mid_4to8_0 ~/dac_layout
timestamp 1729685583
transform 0 1 19960 -1 0 27360
box 0 0 27360 4720
use mid_4to8  mid_4to8_1
timestamp 1729685583
transform 0 1 24950 -1 0 27360
box 0 0 27360 4720
use mid_4to8  mid_4to8_2
timestamp 1729685583
transform 0 1 49900 -1 0 27360
box 0 0 27360 4720
use mid_4to8  mid_4to8_3
timestamp 1729685583
transform 0 1 54890 -1 0 27360
box 0 0 27360 4720
use mid_6to8  mid_6to8_0 ~/dac_layout
timestamp 1729688460
transform 0 1 9980 -1 0 27360
box 0 0 27360 4720
use mid_6to8  mid_6to8_1
timestamp 1729688460
transform 0 1 14970 -1 0 27360
box 0 0 27360 4720
use mid_6to8  mid_6to8_2
timestamp 1729688460
transform 0 1 59880 -1 0 27360
box 0 0 27360 4720
use mid_6to8  mid_6to8_3
timestamp 1729688460
transform 0 1 64870 -1 0 27360
box 0 0 27360 4720
<< labels >>
flabel metal1 2750 64130 2810 64190 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 3820 64130 3880 64190 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 3820 64460 3880 64510 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 3282 64222 3342 64282 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 3282 64672 3342 64732 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 3698 64288 3700 64348 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 3760 64594 3762 64654 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 2860 64290 2920 64350 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 2860 64600 2920 64660 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 2750 64440 2810 64500 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 220 63850 280 63910 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 2750 62420 2810 62480 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 3820 62420 3880 62480 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 3820 62750 3880 62800 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 3282 62512 3342 62572 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 3282 62962 3342 63022 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 3698 62578 3700 62638 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 3760 62884 3762 62944 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 2860 62580 2920 62640 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 2860 62890 2920 62950 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 2750 62730 2810 62790 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 220 62140 280 62200 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 2750 60710 2810 60770 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 3820 60710 3880 60770 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 3820 61040 3880 61090 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 3282 60802 3342 60862 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 3282 61252 3342 61312 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 3698 60868 3700 60928 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 3760 61174 3762 61234 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 2860 60870 2920 60930 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 2860 61180 2920 61240 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 2750 61020 2810 61080 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 220 60430 280 60490 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 2750 59000 2810 59060 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 3820 59000 3880 59060 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 3820 59330 3880 59380 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 3282 59092 3342 59152 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 3282 59542 3342 59602 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 3698 59158 3700 59218 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 3760 59464 3762 59524 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 2860 59160 2920 59220 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 2860 59470 2920 59530 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 2750 59310 2810 59370 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 220 58720 280 58780 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 2750 57290 2810 57350 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 3820 57290 3880 57350 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 3820 57620 3880 57670 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 3282 57382 3342 57442 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 3282 57832 3342 57892 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 3698 57448 3700 57508 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 3760 57754 3762 57814 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 2860 57450 2920 57510 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 2860 57760 2920 57820 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 2750 57600 2810 57660 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 220 57010 280 57070 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 2750 55580 2810 55640 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 3820 55580 3880 55640 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 3820 55910 3880 55960 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 3282 55672 3342 55732 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 3282 56122 3342 56182 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 3698 55738 3700 55798 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 3760 56044 3762 56104 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 2860 55740 2920 55800 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 2860 56050 2920 56110 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 2750 55890 2810 55950 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 220 55300 280 55360 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 2750 65840 2810 65900 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 3820 65840 3880 65900 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 3820 66170 3880 66220 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 3282 65932 3342 65992 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 3282 66382 3342 66442 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 3698 65998 3700 66058 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 3760 66304 3762 66364 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 2860 66000 2920 66060 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 2860 66310 2920 66370 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 2750 66150 2810 66210 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 220 65560 280 65620 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 2750 53870 2810 53930 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 3820 53870 3880 53930 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 3820 54200 3880 54250 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 3282 53962 3342 54022 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 3282 54412 3342 54472 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 3698 54028 3700 54088 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 3760 54334 3762 54394 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 2860 54030 2920 54090 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 2860 54340 2920 54400 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 2750 54180 2810 54240 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 220 53590 280 53650 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 2750 50450 2810 50510 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 3820 50450 3880 50510 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 3820 50780 3880 50830 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 3282 50542 3342 50602 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 3282 50992 3342 51052 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 3698 50608 3700 50668 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 3760 50914 3762 50974 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 2860 50610 2920 50670 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 2860 50920 2920 50980 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 2750 50760 2810 50820 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 220 50170 280 50230 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 2750 48740 2810 48800 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 3820 48740 3880 48800 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 3820 49070 3880 49120 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 3282 48832 3342 48892 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 3282 49282 3342 49342 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 3698 48898 3700 48958 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 3760 49204 3762 49264 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 2860 48900 2920 48960 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 2860 49210 2920 49270 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 2750 49050 2810 49110 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 220 48460 280 48520 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 2750 47030 2810 47090 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 3820 47030 3880 47090 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 3820 47360 3880 47410 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 3282 47122 3342 47182 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 3282 47572 3342 47632 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 3698 47188 3700 47248 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 3760 47494 3762 47554 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 2860 47190 2920 47250 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 2860 47500 2920 47560 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 2750 47340 2810 47400 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 220 46750 280 46810 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 2750 45320 2810 45380 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 3820 45320 3880 45380 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 3820 45650 3880 45700 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 3282 45412 3342 45472 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 3282 45862 3342 45922 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 3698 45478 3700 45538 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 3760 45784 3762 45844 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 2860 45480 2920 45540 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 2860 45790 2920 45850 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 2750 45630 2810 45690 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 220 45040 280 45100 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 2750 43610 2810 43670 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 3820 43610 3880 43670 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 3820 43940 3880 43990 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 3282 43702 3342 43762 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 3282 44152 3342 44212 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 3698 43768 3700 43828 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 3760 44074 3762 44134 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 2860 43770 2920 43830 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 2860 44080 2920 44140 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 2750 43920 2810 43980 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 220 43330 280 43390 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 2750 41900 2810 41960 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 3820 41900 3880 41960 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 3820 42230 3880 42280 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 3282 41992 3342 42052 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 3282 42442 3342 42502 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 3698 42058 3700 42118 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 3760 42364 3762 42424 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 2860 42060 2920 42120 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 2860 42370 2920 42430 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 2750 42210 2810 42270 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 220 41620 280 41680 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 2750 52160 2810 52220 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 3820 52160 3880 52220 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 3820 52490 3880 52540 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 3282 52252 3342 52312 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 3282 52702 3342 52762 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 3698 52318 3700 52378 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 3760 52624 3762 52684 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 2860 52320 2920 52380 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 2860 52630 2920 52690 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 2750 52470 2810 52530 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 220 51880 280 51940 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 2750 40190 2810 40250 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 3820 40190 3880 40250 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 3820 40520 3880 40570 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 3282 40282 3342 40342 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 3282 40732 3342 40792 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 3698 40348 3700 40408 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 3760 40654 3762 40714 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 2860 40350 2920 40410 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 2860 40660 2920 40720 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 2750 40500 2810 40560 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 220 39910 280 39970 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 7740 64130 7800 64190 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 8810 64130 8870 64190 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 8810 64460 8870 64510 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 8272 64222 8332 64282 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 8272 64672 8332 64732 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 8688 64288 8690 64348 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 8750 64594 8752 64654 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 7850 64290 7910 64350 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 7850 64600 7910 64660 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 7740 64440 7800 64500 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 5210 63850 5270 63910 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 7740 62420 7800 62480 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 8810 62420 8870 62480 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 8810 62750 8870 62800 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 8272 62512 8332 62572 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 8272 62962 8332 63022 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 8688 62578 8690 62638 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 8750 62884 8752 62944 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 7850 62580 7910 62640 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 7850 62890 7910 62950 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 7740 62730 7800 62790 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 5210 62140 5270 62200 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 7740 60710 7800 60770 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 8810 60710 8870 60770 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 8810 61040 8870 61090 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 8272 60802 8332 60862 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 8272 61252 8332 61312 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 8688 60868 8690 60928 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 8750 61174 8752 61234 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 7850 60870 7910 60930 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 7850 61180 7910 61240 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 7740 61020 7800 61080 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 5210 60430 5270 60490 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 7740 59000 7800 59060 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 8810 59000 8870 59060 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 8810 59330 8870 59380 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 8272 59092 8332 59152 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 8272 59542 8332 59602 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 8688 59158 8690 59218 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 8750 59464 8752 59524 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 7850 59160 7910 59220 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 7850 59470 7910 59530 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 7740 59310 7800 59370 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 5210 58720 5270 58780 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 7740 57290 7800 57350 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 8810 57290 8870 57350 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 8810 57620 8870 57670 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 8272 57382 8332 57442 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 8272 57832 8332 57892 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 8688 57448 8690 57508 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 8750 57754 8752 57814 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 7850 57450 7910 57510 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 7850 57760 7910 57820 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 7740 57600 7800 57660 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 5210 57010 5270 57070 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 7740 55580 7800 55640 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 8810 55580 8870 55640 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 8810 55910 8870 55960 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 8272 55672 8332 55732 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 8272 56122 8332 56182 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 8688 55738 8690 55798 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 8750 56044 8752 56104 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 7850 55740 7910 55800 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 7850 56050 7910 56110 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 7740 55890 7800 55950 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 5210 55300 5270 55360 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 7740 65840 7800 65900 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 8810 65840 8870 65900 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 8810 66170 8870 66220 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 8272 65932 8332 65992 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 8272 66382 8332 66442 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 8688 65998 8690 66058 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 8750 66304 8752 66364 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 7850 66000 7910 66060 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 7850 66310 7910 66370 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 7740 66150 7800 66210 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 5210 65560 5270 65620 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 7740 53870 7800 53930 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 8810 53870 8870 53930 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 8810 54200 8870 54250 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 8272 53962 8332 54022 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 8272 54412 8332 54472 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 8688 54028 8690 54088 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 8750 54334 8752 54394 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 7850 54030 7910 54090 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 7850 54340 7910 54400 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 7740 54180 7800 54240 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 5210 53590 5270 53650 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 7740 50450 7800 50510 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 8810 50450 8870 50510 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 8810 50780 8870 50830 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 8272 50542 8332 50602 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 8272 50992 8332 51052 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 8688 50608 8690 50668 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 8750 50914 8752 50974 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 7850 50610 7910 50670 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 7850 50920 7910 50980 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 7740 50760 7800 50820 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 5210 50170 5270 50230 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 7740 48740 7800 48800 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 8810 48740 8870 48800 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 8810 49070 8870 49120 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 8272 48832 8332 48892 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 8272 49282 8332 49342 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 8688 48898 8690 48958 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 8750 49204 8752 49264 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 7850 48900 7910 48960 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 7850 49210 7910 49270 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 7740 49050 7800 49110 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 5210 48460 5270 48520 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 7740 47030 7800 47090 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 8810 47030 8870 47090 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 8810 47360 8870 47410 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 8272 47122 8332 47182 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 8272 47572 8332 47632 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 8688 47188 8690 47248 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 8750 47494 8752 47554 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 7850 47190 7910 47250 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 7850 47500 7910 47560 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 7740 47340 7800 47400 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 5210 46750 5270 46810 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 7740 45320 7800 45380 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 8810 45320 8870 45380 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 8810 45650 8870 45700 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 8272 45412 8332 45472 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 8272 45862 8332 45922 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 8688 45478 8690 45538 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 8750 45784 8752 45844 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 7850 45480 7910 45540 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 7850 45790 7910 45850 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 7740 45630 7800 45690 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 5210 45040 5270 45100 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 7740 43610 7800 43670 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 8810 43610 8870 43670 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 8810 43940 8870 43990 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 8272 43702 8332 43762 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 8272 44152 8332 44212 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 8688 43768 8690 43828 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 8750 44074 8752 44134 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 7850 43770 7910 43830 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 7850 44080 7910 44140 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 7740 43920 7800 43980 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 5210 43330 5270 43390 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 7740 41900 7800 41960 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 8810 41900 8870 41960 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 8810 42230 8870 42280 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 8272 41992 8332 42052 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 8272 42442 8332 42502 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 8688 42058 8690 42118 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 8750 42364 8752 42424 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 7850 42060 7910 42120 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 7850 42370 7910 42430 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 7740 42210 7800 42270 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 5210 41620 5270 41680 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 7740 52160 7800 52220 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 8810 52160 8870 52220 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 8810 52490 8870 52540 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 8272 52252 8332 52312 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 8272 52702 8332 52762 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 8688 52318 8690 52378 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 8750 52624 8752 52684 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 7850 52320 7910 52380 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 7850 52630 7910 52690 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 7740 52470 7800 52530 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 5210 51880 5270 51940 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 7740 40190 7800 40250 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 8810 40190 8870 40250 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 8810 40520 8870 40570 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 8272 40282 8332 40342 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 8272 40732 8332 40792 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 8688 40348 8690 40408 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 8750 40654 8752 40714 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 7850 40350 7910 40410 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 7850 40660 7910 40720 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 7740 40500 7800 40560 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 5210 39910 5270 39970 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 12730 64130 12790 64190 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 13800 64130 13860 64190 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 13800 64460 13860 64510 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 13262 64222 13322 64282 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 13262 64672 13322 64732 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 13678 64288 13680 64348 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 13740 64594 13742 64654 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 12840 64290 12900 64350 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 12840 64600 12900 64660 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 12730 64440 12790 64500 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 10200 63850 10260 63910 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 12730 62420 12790 62480 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 13800 62420 13860 62480 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 13800 62750 13860 62800 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 13262 62512 13322 62572 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 13262 62962 13322 63022 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 13678 62578 13680 62638 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 13740 62884 13742 62944 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 12840 62580 12900 62640 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 12840 62890 12900 62950 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 12730 62730 12790 62790 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 10200 62140 10260 62200 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 12730 60710 12790 60770 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 13800 60710 13860 60770 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 13800 61040 13860 61090 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 13262 60802 13322 60862 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 13262 61252 13322 61312 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 13678 60868 13680 60928 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 13740 61174 13742 61234 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 12840 60870 12900 60930 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 12840 61180 12900 61240 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 12730 61020 12790 61080 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 10200 60430 10260 60490 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 12730 59000 12790 59060 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 13800 59000 13860 59060 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 13800 59330 13860 59380 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 13262 59092 13322 59152 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 13262 59542 13322 59602 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 13678 59158 13680 59218 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 13740 59464 13742 59524 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 12840 59160 12900 59220 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 12840 59470 12900 59530 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 12730 59310 12790 59370 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 10200 58720 10260 58780 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 12730 57290 12790 57350 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 13800 57290 13860 57350 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 13800 57620 13860 57670 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 13262 57382 13322 57442 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 13262 57832 13322 57892 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 13678 57448 13680 57508 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 13740 57754 13742 57814 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 12840 57450 12900 57510 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 12840 57760 12900 57820 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 12730 57600 12790 57660 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 10200 57010 10260 57070 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 12730 55580 12790 55640 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 13800 55580 13860 55640 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 13800 55910 13860 55960 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 13262 55672 13322 55732 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 13262 56122 13322 56182 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 13678 55738 13680 55798 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 13740 56044 13742 56104 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 12840 55740 12900 55800 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 12840 56050 12900 56110 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 12730 55890 12790 55950 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 10200 55300 10260 55360 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 12730 65840 12790 65900 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 13800 65840 13860 65900 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 13800 66170 13860 66220 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 13262 65932 13322 65992 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 13262 66382 13322 66442 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 13678 65998 13680 66058 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 13740 66304 13742 66364 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 12840 66000 12900 66060 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 12840 66310 12900 66370 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 12730 66150 12790 66210 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 10200 65560 10260 65620 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 12730 53870 12790 53930 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 13800 53870 13860 53930 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 13800 54200 13860 54250 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 13262 53962 13322 54022 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 13262 54412 13322 54472 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 13678 54028 13680 54088 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 13740 54334 13742 54394 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 12840 54030 12900 54090 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 12840 54340 12900 54400 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 12730 54180 12790 54240 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 10200 53590 10260 53650 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 12730 50450 12790 50510 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 13800 50450 13860 50510 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 13800 50780 13860 50830 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 13262 50542 13322 50602 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 13262 50992 13322 51052 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 13678 50608 13680 50668 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 13740 50914 13742 50974 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 12840 50610 12900 50670 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 12840 50920 12900 50980 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 12730 50760 12790 50820 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 10200 50170 10260 50230 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 12730 48740 12790 48800 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 13800 48740 13860 48800 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 13800 49070 13860 49120 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 13262 48832 13322 48892 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 13262 49282 13322 49342 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 13678 48898 13680 48958 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 13740 49204 13742 49264 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 12840 48900 12900 48960 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 12840 49210 12900 49270 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 12730 49050 12790 49110 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 10200 48460 10260 48520 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 12730 47030 12790 47090 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 13800 47030 13860 47090 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 13800 47360 13860 47410 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 13262 47122 13322 47182 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 13262 47572 13322 47632 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 13678 47188 13680 47248 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 13740 47494 13742 47554 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 12840 47190 12900 47250 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 12840 47500 12900 47560 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 12730 47340 12790 47400 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 10200 46750 10260 46810 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 12730 45320 12790 45380 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 13800 45320 13860 45380 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 13800 45650 13860 45700 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 13262 45412 13322 45472 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 13262 45862 13322 45922 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 13678 45478 13680 45538 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 13740 45784 13742 45844 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 12840 45480 12900 45540 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 12840 45790 12900 45850 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 12730 45630 12790 45690 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 10200 45040 10260 45100 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 12730 43610 12790 43670 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 13800 43610 13860 43670 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 13800 43940 13860 43990 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 13262 43702 13322 43762 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 13262 44152 13322 44212 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 13678 43768 13680 43828 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 13740 44074 13742 44134 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 12840 43770 12900 43830 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 12840 44080 12900 44140 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 12730 43920 12790 43980 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 10200 43330 10260 43390 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 12730 41900 12790 41960 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 13800 41900 13860 41960 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 13800 42230 13860 42280 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 13262 41992 13322 42052 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 13262 42442 13322 42502 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 13678 42058 13680 42118 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 13740 42364 13742 42424 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 12840 42060 12900 42120 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 12840 42370 12900 42430 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 12730 42210 12790 42270 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 10200 41620 10260 41680 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 12730 52160 12790 52220 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 13800 52160 13860 52220 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 13800 52490 13860 52540 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 13262 52252 13322 52312 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 13262 52702 13322 52762 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 13678 52318 13680 52378 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 13740 52624 13742 52684 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 12840 52320 12900 52380 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 12840 52630 12900 52690 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 12730 52470 12790 52530 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 10200 51880 10260 51940 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 12730 40190 12790 40250 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 13800 40190 13860 40250 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 13800 40520 13860 40570 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 13262 40282 13322 40342 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 13262 40732 13322 40792 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 13678 40348 13680 40408 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 13740 40654 13742 40714 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 12840 40350 12900 40410 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 12840 40660 12900 40720 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 12730 40500 12790 40560 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 10200 39910 10260 39970 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 17720 64130 17780 64190 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 18790 64130 18850 64190 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 18790 64460 18850 64510 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 18252 64222 18312 64282 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 18252 64672 18312 64732 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 18668 64288 18670 64348 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 18730 64594 18732 64654 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 17830 64290 17890 64350 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 17830 64600 17890 64660 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 17720 64440 17780 64500 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 15190 63850 15250 63910 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 17720 62420 17780 62480 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 18790 62420 18850 62480 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 18790 62750 18850 62800 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 18252 62512 18312 62572 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 18252 62962 18312 63022 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 18668 62578 18670 62638 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 18730 62884 18732 62944 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 17830 62580 17890 62640 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 17830 62890 17890 62950 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 17720 62730 17780 62790 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 15190 62140 15250 62200 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 17720 60710 17780 60770 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 18790 60710 18850 60770 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 18790 61040 18850 61090 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 18252 60802 18312 60862 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 18252 61252 18312 61312 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 18668 60868 18670 60928 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 18730 61174 18732 61234 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 17830 60870 17890 60930 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 17830 61180 17890 61240 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 17720 61020 17780 61080 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 15190 60430 15250 60490 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 17720 59000 17780 59060 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 18790 59000 18850 59060 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 18790 59330 18850 59380 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 18252 59092 18312 59152 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 18252 59542 18312 59602 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 18668 59158 18670 59218 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 18730 59464 18732 59524 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 17830 59160 17890 59220 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 17830 59470 17890 59530 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 17720 59310 17780 59370 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 15190 58720 15250 58780 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 17720 57290 17780 57350 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 18790 57290 18850 57350 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 18790 57620 18850 57670 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 18252 57382 18312 57442 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 18252 57832 18312 57892 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 18668 57448 18670 57508 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 18730 57754 18732 57814 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 17830 57450 17890 57510 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 17830 57760 17890 57820 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 17720 57600 17780 57660 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 15190 57010 15250 57070 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 17720 55580 17780 55640 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 18790 55580 18850 55640 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 18790 55910 18850 55960 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 18252 55672 18312 55732 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 18252 56122 18312 56182 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 18668 55738 18670 55798 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 18730 56044 18732 56104 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 17830 55740 17890 55800 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 17830 56050 17890 56110 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 17720 55890 17780 55950 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 15190 55300 15250 55360 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 17720 65840 17780 65900 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 18790 65840 18850 65900 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 18790 66170 18850 66220 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 18252 65932 18312 65992 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 18252 66382 18312 66442 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 18668 65998 18670 66058 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 18730 66304 18732 66364 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 17830 66000 17890 66060 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 17830 66310 17890 66370 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 17720 66150 17780 66210 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 15190 65560 15250 65620 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 17720 53870 17780 53930 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 18790 53870 18850 53930 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 18790 54200 18850 54250 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 18252 53962 18312 54022 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 18252 54412 18312 54472 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 18668 54028 18670 54088 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 18730 54334 18732 54394 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 17830 54030 17890 54090 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 17830 54340 17890 54400 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 17720 54180 17780 54240 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 15190 53590 15250 53650 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 17720 50450 17780 50510 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 18790 50450 18850 50510 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 18790 50780 18850 50830 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 18252 50542 18312 50602 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 18252 50992 18312 51052 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 18668 50608 18670 50668 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 18730 50914 18732 50974 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 17830 50610 17890 50670 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 17830 50920 17890 50980 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 17720 50760 17780 50820 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 15190 50170 15250 50230 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 17720 48740 17780 48800 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 18790 48740 18850 48800 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 18790 49070 18850 49120 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 18252 48832 18312 48892 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 18252 49282 18312 49342 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 18668 48898 18670 48958 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 18730 49204 18732 49264 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 17830 48900 17890 48960 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 17830 49210 17890 49270 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 17720 49050 17780 49110 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 15190 48460 15250 48520 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 17720 47030 17780 47090 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 18790 47030 18850 47090 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 18790 47360 18850 47410 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 18252 47122 18312 47182 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 18252 47572 18312 47632 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 18668 47188 18670 47248 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 18730 47494 18732 47554 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 17830 47190 17890 47250 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 17830 47500 17890 47560 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 17720 47340 17780 47400 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 15190 46750 15250 46810 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 17720 45320 17780 45380 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 18790 45320 18850 45380 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 18790 45650 18850 45700 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 18252 45412 18312 45472 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 18252 45862 18312 45922 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 18668 45478 18670 45538 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 18730 45784 18732 45844 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 17830 45480 17890 45540 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 17830 45790 17890 45850 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 17720 45630 17780 45690 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 15190 45040 15250 45100 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 17720 43610 17780 43670 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 18790 43610 18850 43670 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 18790 43940 18850 43990 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 18252 43702 18312 43762 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 18252 44152 18312 44212 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 18668 43768 18670 43828 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 18730 44074 18732 44134 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 17830 43770 17890 43830 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 17830 44080 17890 44140 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 17720 43920 17780 43980 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 15190 43330 15250 43390 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 17720 41900 17780 41960 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 18790 41900 18850 41960 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 18790 42230 18850 42280 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 18252 41992 18312 42052 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 18252 42442 18312 42502 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 18668 42058 18670 42118 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 18730 42364 18732 42424 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 17830 42060 17890 42120 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 17830 42370 17890 42430 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 17720 42210 17780 42270 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 15190 41620 15250 41680 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 17720 52160 17780 52220 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 18790 52160 18850 52220 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 18790 52490 18850 52540 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 18252 52252 18312 52312 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 18252 52702 18312 52762 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 18668 52318 18670 52378 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 18730 52624 18732 52684 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 17830 52320 17890 52380 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 17830 52630 17890 52690 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 17720 52470 17780 52530 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 15190 51880 15250 51940 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 17720 40190 17780 40250 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 18790 40190 18850 40250 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 18790 40520 18850 40570 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 18252 40282 18312 40342 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 18252 40732 18312 40792 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 18668 40348 18670 40408 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 18730 40654 18732 40714 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 17830 40350 17890 40410 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 17830 40660 17890 40720 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 17720 40500 17780 40560 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 15190 39910 15250 39970 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 22710 64130 22770 64190 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 23780 64130 23840 64190 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 23780 64460 23840 64510 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 23242 64222 23302 64282 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 23242 64672 23302 64732 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 23658 64288 23660 64348 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 23720 64594 23722 64654 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 22820 64290 22880 64350 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 22820 64600 22880 64660 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 22710 64440 22770 64500 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 20180 63850 20240 63910 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 22710 62420 22770 62480 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 23780 62420 23840 62480 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 23780 62750 23840 62800 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 23242 62512 23302 62572 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 23242 62962 23302 63022 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 23658 62578 23660 62638 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 23720 62884 23722 62944 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 22820 62580 22880 62640 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 22820 62890 22880 62950 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 22710 62730 22770 62790 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 20180 62140 20240 62200 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 22710 60710 22770 60770 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 23780 60710 23840 60770 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 23780 61040 23840 61090 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 23242 60802 23302 60862 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 23242 61252 23302 61312 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 23658 60868 23660 60928 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 23720 61174 23722 61234 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 22820 60870 22880 60930 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 22820 61180 22880 61240 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 22710 61020 22770 61080 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 20180 60430 20240 60490 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 22710 59000 22770 59060 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 23780 59000 23840 59060 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 23780 59330 23840 59380 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 23242 59092 23302 59152 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 23242 59542 23302 59602 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 23658 59158 23660 59218 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 23720 59464 23722 59524 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 22820 59160 22880 59220 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 22820 59470 22880 59530 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 22710 59310 22770 59370 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 20180 58720 20240 58780 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 22710 57290 22770 57350 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 23780 57290 23840 57350 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 23780 57620 23840 57670 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 23242 57382 23302 57442 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 23242 57832 23302 57892 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 23658 57448 23660 57508 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 23720 57754 23722 57814 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 22820 57450 22880 57510 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 22820 57760 22880 57820 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 22710 57600 22770 57660 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 20180 57010 20240 57070 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 22710 55580 22770 55640 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 23780 55580 23840 55640 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 23780 55910 23840 55960 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 23242 55672 23302 55732 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 23242 56122 23302 56182 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 23658 55738 23660 55798 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 23720 56044 23722 56104 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 22820 55740 22880 55800 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 22820 56050 22880 56110 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 22710 55890 22770 55950 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 20180 55300 20240 55360 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 22710 65840 22770 65900 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 23780 65840 23840 65900 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 23780 66170 23840 66220 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 23242 65932 23302 65992 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 23242 66382 23302 66442 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 23658 65998 23660 66058 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 23720 66304 23722 66364 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 22820 66000 22880 66060 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 22820 66310 22880 66370 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 22710 66150 22770 66210 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 20180 65560 20240 65620 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 22710 53870 22770 53930 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 23780 53870 23840 53930 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 23780 54200 23840 54250 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 23242 53962 23302 54022 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 23242 54412 23302 54472 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 23658 54028 23660 54088 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 23720 54334 23722 54394 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 22820 54030 22880 54090 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 22820 54340 22880 54400 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 22710 54180 22770 54240 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 20180 53590 20240 53650 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 22710 50450 22770 50510 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 23780 50450 23840 50510 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 23780 50780 23840 50830 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 23242 50542 23302 50602 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 23242 50992 23302 51052 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 23658 50608 23660 50668 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 23720 50914 23722 50974 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 22820 50610 22880 50670 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 22820 50920 22880 50980 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 22710 50760 22770 50820 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 20180 50170 20240 50230 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 22710 48740 22770 48800 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 23780 48740 23840 48800 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 23780 49070 23840 49120 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 23242 48832 23302 48892 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 23242 49282 23302 49342 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 23658 48898 23660 48958 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 23720 49204 23722 49264 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 22820 48900 22880 48960 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 22820 49210 22880 49270 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 22710 49050 22770 49110 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 20180 48460 20240 48520 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 22710 47030 22770 47090 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 23780 47030 23840 47090 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 23780 47360 23840 47410 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 23242 47122 23302 47182 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 23242 47572 23302 47632 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 23658 47188 23660 47248 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 23720 47494 23722 47554 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 22820 47190 22880 47250 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 22820 47500 22880 47560 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 22710 47340 22770 47400 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 20180 46750 20240 46810 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 22710 45320 22770 45380 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 23780 45320 23840 45380 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 23780 45650 23840 45700 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 23242 45412 23302 45472 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 23242 45862 23302 45922 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 23658 45478 23660 45538 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 23720 45784 23722 45844 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 22820 45480 22880 45540 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 22820 45790 22880 45850 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 22710 45630 22770 45690 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 20180 45040 20240 45100 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 22710 43610 22770 43670 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 23780 43610 23840 43670 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 23780 43940 23840 43990 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 23242 43702 23302 43762 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 23242 44152 23302 44212 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 23658 43768 23660 43828 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 23720 44074 23722 44134 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 22820 43770 22880 43830 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 22820 44080 22880 44140 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 22710 43920 22770 43980 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 20180 43330 20240 43390 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 22710 41900 22770 41960 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 23780 41900 23840 41960 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 23780 42230 23840 42280 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 23242 41992 23302 42052 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 23242 42442 23302 42502 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 23658 42058 23660 42118 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 23720 42364 23722 42424 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 22820 42060 22880 42120 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 22820 42370 22880 42430 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 22710 42210 22770 42270 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 20180 41620 20240 41680 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 22710 52160 22770 52220 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 23780 52160 23840 52220 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 23780 52490 23840 52540 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 23242 52252 23302 52312 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 23242 52702 23302 52762 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 23658 52318 23660 52378 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 23720 52624 23722 52684 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 22820 52320 22880 52380 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 22820 52630 22880 52690 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 22710 52470 22770 52530 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 20180 51880 20240 51940 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 22710 40190 22770 40250 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 23780 40190 23840 40250 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 23780 40520 23840 40570 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 23242 40282 23302 40342 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 23242 40732 23302 40792 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 23658 40348 23660 40408 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 23720 40654 23722 40714 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 22820 40350 22880 40410 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 22820 40660 22880 40720 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 22710 40500 22770 40560 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 20180 39910 20240 39970 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 27700 64130 27760 64190 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 28770 64130 28830 64190 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 28770 64460 28830 64510 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 28232 64222 28292 64282 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 28232 64672 28292 64732 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 28648 64288 28650 64348 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 28710 64594 28712 64654 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 27810 64290 27870 64350 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 27810 64600 27870 64660 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 27700 64440 27760 64500 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 25170 63850 25230 63910 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 27700 62420 27760 62480 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 28770 62420 28830 62480 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 28770 62750 28830 62800 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 28232 62512 28292 62572 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 28232 62962 28292 63022 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 28648 62578 28650 62638 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 28710 62884 28712 62944 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 27810 62580 27870 62640 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 27810 62890 27870 62950 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 27700 62730 27760 62790 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 25170 62140 25230 62200 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 27700 60710 27760 60770 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 28770 60710 28830 60770 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 28770 61040 28830 61090 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 28232 60802 28292 60862 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 28232 61252 28292 61312 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 28648 60868 28650 60928 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 28710 61174 28712 61234 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 27810 60870 27870 60930 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 27810 61180 27870 61240 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 27700 61020 27760 61080 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 25170 60430 25230 60490 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 27700 59000 27760 59060 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 28770 59000 28830 59060 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 28770 59330 28830 59380 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 28232 59092 28292 59152 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 28232 59542 28292 59602 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 28648 59158 28650 59218 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 28710 59464 28712 59524 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 27810 59160 27870 59220 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 27810 59470 27870 59530 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 27700 59310 27760 59370 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 25170 58720 25230 58780 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 27700 57290 27760 57350 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 28770 57290 28830 57350 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 28770 57620 28830 57670 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 28232 57382 28292 57442 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 28232 57832 28292 57892 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 28648 57448 28650 57508 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 28710 57754 28712 57814 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 27810 57450 27870 57510 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 27810 57760 27870 57820 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 27700 57600 27760 57660 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 25170 57010 25230 57070 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 27700 55580 27760 55640 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 28770 55580 28830 55640 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 28770 55910 28830 55960 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 28232 55672 28292 55732 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 28232 56122 28292 56182 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 28648 55738 28650 55798 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 28710 56044 28712 56104 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 27810 55740 27870 55800 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 27810 56050 27870 56110 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 27700 55890 27760 55950 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 25170 55300 25230 55360 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 27700 65840 27760 65900 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 28770 65840 28830 65900 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 28770 66170 28830 66220 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 28232 65932 28292 65992 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 28232 66382 28292 66442 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 28648 65998 28650 66058 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 28710 66304 28712 66364 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 27810 66000 27870 66060 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 27810 66310 27870 66370 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 27700 66150 27760 66210 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 25170 65560 25230 65620 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 27700 53870 27760 53930 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 28770 53870 28830 53930 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 28770 54200 28830 54250 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 28232 53962 28292 54022 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 28232 54412 28292 54472 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 28648 54028 28650 54088 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 28710 54334 28712 54394 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 27810 54030 27870 54090 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 27810 54340 27870 54400 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 27700 54180 27760 54240 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 25170 53590 25230 53650 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 27700 50450 27760 50510 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 28770 50450 28830 50510 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 28770 50780 28830 50830 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 28232 50542 28292 50602 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 28232 50992 28292 51052 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 28648 50608 28650 50668 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 28710 50914 28712 50974 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 27810 50610 27870 50670 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 27810 50920 27870 50980 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 27700 50760 27760 50820 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 25170 50170 25230 50230 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 27700 48740 27760 48800 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 28770 48740 28830 48800 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 28770 49070 28830 49120 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 28232 48832 28292 48892 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 28232 49282 28292 49342 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 28648 48898 28650 48958 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 28710 49204 28712 49264 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 27810 48900 27870 48960 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 27810 49210 27870 49270 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 27700 49050 27760 49110 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 25170 48460 25230 48520 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 27700 47030 27760 47090 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 28770 47030 28830 47090 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 28770 47360 28830 47410 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 28232 47122 28292 47182 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 28232 47572 28292 47632 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 28648 47188 28650 47248 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 28710 47494 28712 47554 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 27810 47190 27870 47250 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 27810 47500 27870 47560 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 27700 47340 27760 47400 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 25170 46750 25230 46810 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 27700 45320 27760 45380 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 28770 45320 28830 45380 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 28770 45650 28830 45700 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 28232 45412 28292 45472 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 28232 45862 28292 45922 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 28648 45478 28650 45538 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 28710 45784 28712 45844 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 27810 45480 27870 45540 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 27810 45790 27870 45850 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 27700 45630 27760 45690 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 25170 45040 25230 45100 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 27700 43610 27760 43670 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 28770 43610 28830 43670 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 28770 43940 28830 43990 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 28232 43702 28292 43762 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 28232 44152 28292 44212 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 28648 43768 28650 43828 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 28710 44074 28712 44134 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 27810 43770 27870 43830 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 27810 44080 27870 44140 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 27700 43920 27760 43980 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 25170 43330 25230 43390 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 27700 41900 27760 41960 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 28770 41900 28830 41960 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 28770 42230 28830 42280 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 28232 41992 28292 42052 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 28232 42442 28292 42502 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 28648 42058 28650 42118 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 28710 42364 28712 42424 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 27810 42060 27870 42120 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 27810 42370 27870 42430 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 27700 42210 27760 42270 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 25170 41620 25230 41680 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 27700 52160 27760 52220 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 28770 52160 28830 52220 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 28770 52490 28830 52540 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 28232 52252 28292 52312 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 28232 52702 28292 52762 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 28648 52318 28650 52378 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 28710 52624 28712 52684 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 27810 52320 27870 52380 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 27810 52630 27870 52690 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 27700 52470 27760 52530 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 25170 51880 25230 51940 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 27700 40190 27760 40250 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 28770 40190 28830 40250 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 28770 40520 28830 40570 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 28232 40282 28292 40342 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 28232 40732 28292 40792 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 28648 40348 28650 40408 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 28710 40654 28712 40714 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 27810 40350 27870 40410 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 27810 40660 27870 40720 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 27700 40500 27760 40560 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 25170 39910 25230 39970 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 42670 50450 42730 50510 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 43740 50450 43800 50510 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 43740 50780 43800 50830 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 43202 50542 43262 50602 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 43202 50992 43262 51052 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 43618 50608 43620 50668 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 43680 50914 43682 50974 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 42780 50610 42840 50670 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 42780 50920 42840 50980 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 42670 50760 42730 50820 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 40140 50170 40200 50230 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 42670 48740 42730 48800 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 43740 48740 43800 48800 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 43740 49070 43800 49120 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 43202 48832 43262 48892 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 43202 49282 43262 49342 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 43618 48898 43620 48958 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 43680 49204 43682 49264 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 42780 48900 42840 48960 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 42780 49210 42840 49270 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 42670 49050 42730 49110 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 40140 48460 40200 48520 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 42670 47030 42730 47090 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 43740 47030 43800 47090 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 43740 47360 43800 47410 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 43202 47122 43262 47182 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 43202 47572 43262 47632 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 43618 47188 43620 47248 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 43680 47494 43682 47554 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 42780 47190 42840 47250 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 42780 47500 42840 47560 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 42670 47340 42730 47400 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 40140 46750 40200 46810 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 42670 45320 42730 45380 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 43740 45320 43800 45380 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 43740 45650 43800 45700 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 43202 45412 43262 45472 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 43202 45862 43262 45922 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 43618 45478 43620 45538 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 43680 45784 43682 45844 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 42780 45480 42840 45540 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 42780 45790 42840 45850 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 42670 45630 42730 45690 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 40140 45040 40200 45100 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 42670 43610 42730 43670 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 43740 43610 43800 43670 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 43740 43940 43800 43990 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 43202 43702 43262 43762 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 43202 44152 43262 44212 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 43618 43768 43620 43828 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 43680 44074 43682 44134 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 42780 43770 42840 43830 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 42780 44080 42840 44140 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 42670 43920 42730 43980 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 40140 43330 40200 43390 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 42670 41900 42730 41960 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 43740 41900 43800 41960 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 43740 42230 43800 42280 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 43202 41992 43262 42052 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 43202 42442 43262 42502 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 43618 42058 43620 42118 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 43680 42364 43682 42424 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 42780 42060 42840 42120 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 42780 42370 42840 42430 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 42670 42210 42730 42270 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 40140 41620 40200 41680 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 42670 52160 42730 52220 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 43740 52160 43800 52220 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 43740 52490 43800 52540 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 43202 52252 43262 52312 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 43202 52702 43262 52762 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 43618 52318 43620 52378 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 43680 52624 43682 52684 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 42780 52320 42840 52380 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 42780 52630 42840 52690 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 42670 52470 42730 52530 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 40140 51880 40200 51940 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 42670 40190 42730 40250 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 43740 40190 43800 40250 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 43740 40520 43800 40570 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 43202 40282 43262 40342 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 43202 40732 43262 40792 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 43618 40348 43620 40408 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 43680 40654 43682 40714 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 42780 40350 42840 40410 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 42780 40660 42840 40720 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 42670 40500 42730 40560 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 40140 39910 40200 39970 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 37680 50450 37740 50510 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 38750 50450 38810 50510 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 38750 50780 38810 50830 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 38212 50542 38272 50602 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 38212 50992 38272 51052 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 38628 50608 38630 50668 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 38690 50914 38692 50974 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 37790 50610 37850 50670 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 37790 50920 37850 50980 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 37680 50760 37740 50820 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 35150 50170 35210 50230 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 37680 48740 37740 48800 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 38750 48740 38810 48800 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 38750 49070 38810 49120 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 38212 48832 38272 48892 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 38212 49282 38272 49342 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 38628 48898 38630 48958 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 38690 49204 38692 49264 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 37790 48900 37850 48960 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 37790 49210 37850 49270 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 37680 49050 37740 49110 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 35150 48460 35210 48520 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 37680 47030 37740 47090 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 38750 47030 38810 47090 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 38750 47360 38810 47410 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 38212 47122 38272 47182 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 38212 47572 38272 47632 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 38628 47188 38630 47248 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 38690 47494 38692 47554 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 37790 47190 37850 47250 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 37790 47500 37850 47560 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 37680 47340 37740 47400 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 35150 46750 35210 46810 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 37680 45320 37740 45380 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 38750 45320 38810 45380 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 38750 45650 38810 45700 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 38212 45412 38272 45472 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 38212 45862 38272 45922 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 38628 45478 38630 45538 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 38690 45784 38692 45844 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 37790 45480 37850 45540 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 37790 45790 37850 45850 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 37680 45630 37740 45690 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 35150 45040 35210 45100 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 37680 43610 37740 43670 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 38750 43610 38810 43670 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 38750 43940 38810 43990 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 38212 43702 38272 43762 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 38212 44152 38272 44212 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 38628 43768 38630 43828 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 38690 44074 38692 44134 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 37790 43770 37850 43830 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 37790 44080 37850 44140 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 37680 43920 37740 43980 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 35150 43330 35210 43390 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 37680 41900 37740 41960 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 38750 41900 38810 41960 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 38750 42230 38810 42280 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 38212 41992 38272 42052 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 38212 42442 38272 42502 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 38628 42058 38630 42118 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 38690 42364 38692 42424 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 37790 42060 37850 42120 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 37790 42370 37850 42430 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 37680 42210 37740 42270 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 35150 41620 35210 41680 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 37680 52160 37740 52220 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 38750 52160 38810 52220 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 38750 52490 38810 52540 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 38212 52252 38272 52312 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 38212 52702 38272 52762 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 38628 52318 38630 52378 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 38690 52624 38692 52684 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 37790 52320 37850 52380 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 37790 52630 37850 52690 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 37680 52470 37740 52530 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 35150 51880 35210 51940 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 37680 40190 37740 40250 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 38750 40190 38810 40250 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 38750 40520 38810 40570 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 38212 40282 38272 40342 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 38212 40732 38272 40792 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 38628 40348 38630 40408 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 38690 40654 38692 40714 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 37790 40350 37850 40410 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 37790 40660 37850 40720 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 37680 40500 37740 40560 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 35150 39910 35210 39970 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 42670 64130 42730 64190 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 43740 64130 43800 64190 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 43740 64460 43800 64510 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 43202 64222 43262 64282 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 43202 64672 43262 64732 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 43618 64288 43620 64348 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 43680 64594 43682 64654 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 42780 64290 42840 64350 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 42780 64600 42840 64660 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 42670 64440 42730 64500 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 40140 63850 40200 63910 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 42670 62420 42730 62480 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 43740 62420 43800 62480 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 43740 62750 43800 62800 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 43202 62512 43262 62572 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 43202 62962 43262 63022 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 43618 62578 43620 62638 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 43680 62884 43682 62944 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 42780 62580 42840 62640 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 42780 62890 42840 62950 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 42670 62730 42730 62790 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 40140 62140 40200 62200 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 42670 60710 42730 60770 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 43740 60710 43800 60770 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 43740 61040 43800 61090 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 43202 60802 43262 60862 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 43202 61252 43262 61312 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 43618 60868 43620 60928 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 43680 61174 43682 61234 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 42780 60870 42840 60930 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 42780 61180 42840 61240 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 42670 61020 42730 61080 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 40140 60430 40200 60490 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 42670 59000 42730 59060 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 43740 59000 43800 59060 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 43740 59330 43800 59380 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 43202 59092 43262 59152 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 43202 59542 43262 59602 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 43618 59158 43620 59218 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 43680 59464 43682 59524 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 42780 59160 42840 59220 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 42780 59470 42840 59530 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 42670 59310 42730 59370 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 40140 58720 40200 58780 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 42670 57290 42730 57350 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 43740 57290 43800 57350 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 43740 57620 43800 57670 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 43202 57382 43262 57442 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 43202 57832 43262 57892 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 43618 57448 43620 57508 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 43680 57754 43682 57814 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 42780 57450 42840 57510 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 42780 57760 42840 57820 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 42670 57600 42730 57660 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 40140 57010 40200 57070 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 42670 55580 42730 55640 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 43740 55580 43800 55640 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 43740 55910 43800 55960 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 43202 55672 43262 55732 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 43202 56122 43262 56182 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 43618 55738 43620 55798 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 43680 56044 43682 56104 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 42780 55740 42840 55800 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 42780 56050 42840 56110 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 42670 55890 42730 55950 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 40140 55300 40200 55360 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 42670 65840 42730 65900 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 43740 65840 43800 65900 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 43740 66170 43800 66220 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 43202 65932 43262 65992 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 43202 66382 43262 66442 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 43618 65998 43620 66058 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 43680 66304 43682 66364 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 42780 66000 42840 66060 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 42780 66310 42840 66370 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 42670 66150 42730 66210 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 40140 65560 40200 65620 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 42670 53870 42730 53930 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 43740 53870 43800 53930 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 43740 54200 43800 54250 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 43202 53962 43262 54022 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 43202 54412 43262 54472 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 43618 54028 43620 54088 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 43680 54334 43682 54394 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 42780 54030 42840 54090 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 42780 54340 42840 54400 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 42670 54180 42730 54240 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 40140 53590 40200 53650 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 37680 64130 37740 64190 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 38750 64130 38810 64190 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 38750 64460 38810 64510 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 38212 64222 38272 64282 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 38212 64672 38272 64732 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 38628 64288 38630 64348 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 38690 64594 38692 64654 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 37790 64290 37850 64350 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 37790 64600 37850 64660 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 37680 64440 37740 64500 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 35150 63850 35210 63910 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 37680 62420 37740 62480 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 38750 62420 38810 62480 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 38750 62750 38810 62800 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 38212 62512 38272 62572 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 38212 62962 38272 63022 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 38628 62578 38630 62638 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 38690 62884 38692 62944 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 37790 62580 37850 62640 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 37790 62890 37850 62950 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 37680 62730 37740 62790 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 35150 62140 35210 62200 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 37680 60710 37740 60770 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 38750 60710 38810 60770 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 38750 61040 38810 61090 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 38212 60802 38272 60862 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 38212 61252 38272 61312 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 38628 60868 38630 60928 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 38690 61174 38692 61234 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 37790 60870 37850 60930 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 37790 61180 37850 61240 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 37680 61020 37740 61080 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 35150 60430 35210 60490 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 37680 59000 37740 59060 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 38750 59000 38810 59060 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 38750 59330 38810 59380 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 38212 59092 38272 59152 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 38212 59542 38272 59602 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 38628 59158 38630 59218 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 38690 59464 38692 59524 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 37790 59160 37850 59220 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 37790 59470 37850 59530 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 37680 59310 37740 59370 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 35150 58720 35210 58780 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 37680 57290 37740 57350 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 38750 57290 38810 57350 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 38750 57620 38810 57670 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 38212 57382 38272 57442 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 38212 57832 38272 57892 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 38628 57448 38630 57508 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 38690 57754 38692 57814 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 37790 57450 37850 57510 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 37790 57760 37850 57820 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 37680 57600 37740 57660 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 35150 57010 35210 57070 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 37680 55580 37740 55640 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 38750 55580 38810 55640 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 38750 55910 38810 55960 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 38212 55672 38272 55732 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 38212 56122 38272 56182 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 38628 55738 38630 55798 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 38690 56044 38692 56104 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 37790 55740 37850 55800 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 37790 56050 37850 56110 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 37680 55890 37740 55950 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 35150 55300 35210 55360 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 37680 65840 37740 65900 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 38750 65840 38810 65900 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 38750 66170 38810 66220 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 38212 65932 38272 65992 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 38212 66382 38272 66442 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 38628 65998 38630 66058 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 38690 66304 38692 66364 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 37790 66000 37850 66060 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 37790 66310 37850 66370 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 37680 66150 37740 66210 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 35150 65560 35210 65620 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 37680 53870 37740 53930 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 38750 53870 38810 53930 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 38750 54200 38810 54250 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 38212 53962 38272 54022 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 38212 54412 38272 54472 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 38628 54028 38630 54088 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 38690 54334 38692 54394 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 37790 54030 37850 54090 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 37790 54340 37850 54400 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 37680 54180 37740 54240 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 35150 53590 35210 53650 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 32690 64130 32750 64190 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 33760 64130 33820 64190 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 33760 64460 33820 64510 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 33222 64222 33282 64282 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 33222 64672 33282 64732 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 33638 64288 33640 64348 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 33700 64594 33702 64654 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 32800 64290 32860 64350 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 32800 64600 32860 64660 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 32690 64440 32750 64500 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 30160 63850 30220 63910 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 32690 62420 32750 62480 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 33760 62420 33820 62480 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 33760 62750 33820 62800 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 33222 62512 33282 62572 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 33222 62962 33282 63022 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 33638 62578 33640 62638 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 33700 62884 33702 62944 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 32800 62580 32860 62640 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 32800 62890 32860 62950 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 32690 62730 32750 62790 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 30160 62140 30220 62200 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 32690 60710 32750 60770 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 33760 60710 33820 60770 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 33760 61040 33820 61090 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 33222 60802 33282 60862 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 33222 61252 33282 61312 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 33638 60868 33640 60928 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 33700 61174 33702 61234 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 32800 60870 32860 60930 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 32800 61180 32860 61240 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 32690 61020 32750 61080 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 30160 60430 30220 60490 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 32690 59000 32750 59060 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 33760 59000 33820 59060 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 33760 59330 33820 59380 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 33222 59092 33282 59152 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 33222 59542 33282 59602 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 33638 59158 33640 59218 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 33700 59464 33702 59524 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 32800 59160 32860 59220 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 32800 59470 32860 59530 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 32690 59310 32750 59370 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 30160 58720 30220 58780 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 32690 57290 32750 57350 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 33760 57290 33820 57350 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 33760 57620 33820 57670 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 33222 57382 33282 57442 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 33222 57832 33282 57892 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 33638 57448 33640 57508 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 33700 57754 33702 57814 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 32800 57450 32860 57510 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 32800 57760 32860 57820 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 32690 57600 32750 57660 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 30160 57010 30220 57070 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 32690 55580 32750 55640 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 33760 55580 33820 55640 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 33760 55910 33820 55960 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 33222 55672 33282 55732 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 33222 56122 33282 56182 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 33638 55738 33640 55798 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 33700 56044 33702 56104 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 32800 55740 32860 55800 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 32800 56050 32860 56110 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 32690 55890 32750 55950 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 30160 55300 30220 55360 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 32690 65840 32750 65900 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 33760 65840 33820 65900 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 33760 66170 33820 66220 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 33222 65932 33282 65992 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 33222 66382 33282 66442 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 33638 65998 33640 66058 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 33700 66304 33702 66364 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 32800 66000 32860 66060 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 32800 66310 32860 66370 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 32690 66150 32750 66210 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 30160 65560 30220 65620 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 32690 53870 32750 53930 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 33760 53870 33820 53930 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 33760 54200 33820 54250 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 33222 53962 33282 54022 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 33222 54412 33282 54472 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 33638 54028 33640 54088 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 33700 54334 33702 54394 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 32800 54030 32860 54090 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 32800 54340 32860 54400 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 32690 54180 32750 54240 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 30160 53590 30220 53650 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 32690 50450 32750 50510 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 33760 50450 33820 50510 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 33760 50780 33820 50830 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 33222 50542 33282 50602 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 33222 50992 33282 51052 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 33638 50608 33640 50668 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 33700 50914 33702 50974 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 32800 50610 32860 50670 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 32800 50920 32860 50980 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 32690 50760 32750 50820 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 30160 50170 30220 50230 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 32690 48740 32750 48800 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 33760 48740 33820 48800 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 33760 49070 33820 49120 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 33222 48832 33282 48892 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 33222 49282 33282 49342 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 33638 48898 33640 48958 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 33700 49204 33702 49264 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 32800 48900 32860 48960 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 32800 49210 32860 49270 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 32690 49050 32750 49110 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 30160 48460 30220 48520 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 32690 47030 32750 47090 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 33760 47030 33820 47090 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 33760 47360 33820 47410 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 33222 47122 33282 47182 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 33222 47572 33282 47632 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 33638 47188 33640 47248 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 33700 47494 33702 47554 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 32800 47190 32860 47250 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 32800 47500 32860 47560 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 32690 47340 32750 47400 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 30160 46750 30220 46810 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 32690 45320 32750 45380 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 33760 45320 33820 45380 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 33760 45650 33820 45700 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 33222 45412 33282 45472 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 33222 45862 33282 45922 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 33638 45478 33640 45538 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 33700 45784 33702 45844 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 32800 45480 32860 45540 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 32800 45790 32860 45850 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 32690 45630 32750 45690 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 30160 45040 30220 45100 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 32690 43610 32750 43670 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 33760 43610 33820 43670 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 33760 43940 33820 43990 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 33222 43702 33282 43762 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 33222 44152 33282 44212 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 33638 43768 33640 43828 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 33700 44074 33702 44134 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 32800 43770 32860 43830 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 32800 44080 32860 44140 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 32690 43920 32750 43980 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 30160 43330 30220 43390 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 32690 41900 32750 41960 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 33760 41900 33820 41960 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 33760 42230 33820 42280 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 33222 41992 33282 42052 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 33222 42442 33282 42502 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 33638 42058 33640 42118 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 33700 42364 33702 42424 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 32800 42060 32860 42120 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 32800 42370 32860 42430 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 32690 42210 32750 42270 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 30160 41620 30220 41680 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 32690 52160 32750 52220 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 33760 52160 33820 52220 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 33760 52490 33820 52540 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 33222 52252 33282 52312 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 33222 52702 33282 52762 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 33638 52318 33640 52378 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 33700 52624 33702 52684 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 32800 52320 32860 52380 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 32800 52630 32860 52690 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 32690 52470 32750 52530 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 30160 51880 30220 51940 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 32690 40190 32750 40250 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 33760 40190 33820 40250 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 33760 40520 33820 40570 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 33222 40282 33282 40342 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 33222 40732 33282 40792 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 33638 40348 33640 40408 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 33700 40654 33702 40714 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 32800 40350 32860 40410 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 32800 40660 32860 40720 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 32690 40500 32750 40560 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 30160 39910 30220 39970 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 47660 64130 47720 64190 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 48730 64130 48790 64190 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 48730 64460 48790 64510 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 48192 64222 48252 64282 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 48192 64672 48252 64732 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 48608 64288 48610 64348 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 48670 64594 48672 64654 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 47770 64290 47830 64350 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 47770 64600 47830 64660 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 47660 64440 47720 64500 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 45130 63850 45190 63910 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 47660 62420 47720 62480 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 48730 62420 48790 62480 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 48730 62750 48790 62800 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 48192 62512 48252 62572 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 48192 62962 48252 63022 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 48608 62578 48610 62638 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 48670 62884 48672 62944 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 47770 62580 47830 62640 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 47770 62890 47830 62950 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 47660 62730 47720 62790 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 45130 62140 45190 62200 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 47660 60710 47720 60770 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 48730 60710 48790 60770 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 48730 61040 48790 61090 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 48192 60802 48252 60862 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 48192 61252 48252 61312 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 48608 60868 48610 60928 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 48670 61174 48672 61234 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 47770 60870 47830 60930 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 47770 61180 47830 61240 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 47660 61020 47720 61080 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 45130 60430 45190 60490 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 47660 59000 47720 59060 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 48730 59000 48790 59060 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 48730 59330 48790 59380 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 48192 59092 48252 59152 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 48192 59542 48252 59602 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 48608 59158 48610 59218 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 48670 59464 48672 59524 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 47770 59160 47830 59220 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 47770 59470 47830 59530 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 47660 59310 47720 59370 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 45130 58720 45190 58780 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 47660 57290 47720 57350 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 48730 57290 48790 57350 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 48730 57620 48790 57670 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 48192 57382 48252 57442 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 48192 57832 48252 57892 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 48608 57448 48610 57508 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 48670 57754 48672 57814 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 47770 57450 47830 57510 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 47770 57760 47830 57820 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 47660 57600 47720 57660 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 45130 57010 45190 57070 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 47660 55580 47720 55640 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 48730 55580 48790 55640 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 48730 55910 48790 55960 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 48192 55672 48252 55732 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 48192 56122 48252 56182 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 48608 55738 48610 55798 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 48670 56044 48672 56104 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 47770 55740 47830 55800 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 47770 56050 47830 56110 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 47660 55890 47720 55950 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 45130 55300 45190 55360 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 47660 65840 47720 65900 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 48730 65840 48790 65900 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 48730 66170 48790 66220 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 48192 65932 48252 65992 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 48192 66382 48252 66442 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 48608 65998 48610 66058 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 48670 66304 48672 66364 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 47770 66000 47830 66060 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 47770 66310 47830 66370 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 47660 66150 47720 66210 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 45130 65560 45190 65620 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 47660 53870 47720 53930 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 48730 53870 48790 53930 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 48730 54200 48790 54250 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 48192 53962 48252 54022 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 48192 54412 48252 54472 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 48608 54028 48610 54088 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 48670 54334 48672 54394 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 47770 54030 47830 54090 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 47770 54340 47830 54400 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 47660 54180 47720 54240 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 45130 53590 45190 53650 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 47660 50450 47720 50510 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 48730 50450 48790 50510 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 48730 50780 48790 50830 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 48192 50542 48252 50602 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 48192 50992 48252 51052 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 48608 50608 48610 50668 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 48670 50914 48672 50974 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 47770 50610 47830 50670 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 47770 50920 47830 50980 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 47660 50760 47720 50820 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 45130 50170 45190 50230 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 47660 48740 47720 48800 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 48730 48740 48790 48800 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 48730 49070 48790 49120 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 48192 48832 48252 48892 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 48192 49282 48252 49342 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 48608 48898 48610 48958 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 48670 49204 48672 49264 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 47770 48900 47830 48960 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 47770 49210 47830 49270 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 47660 49050 47720 49110 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 45130 48460 45190 48520 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 47660 47030 47720 47090 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 48730 47030 48790 47090 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 48730 47360 48790 47410 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 48192 47122 48252 47182 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 48192 47572 48252 47632 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 48608 47188 48610 47248 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 48670 47494 48672 47554 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 47770 47190 47830 47250 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 47770 47500 47830 47560 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 47660 47340 47720 47400 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 45130 46750 45190 46810 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 47660 45320 47720 45380 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 48730 45320 48790 45380 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 48730 45650 48790 45700 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 48192 45412 48252 45472 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 48192 45862 48252 45922 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 48608 45478 48610 45538 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 48670 45784 48672 45844 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 47770 45480 47830 45540 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 47770 45790 47830 45850 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 47660 45630 47720 45690 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 45130 45040 45190 45100 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 47660 43610 47720 43670 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 48730 43610 48790 43670 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 48730 43940 48790 43990 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 48192 43702 48252 43762 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 48192 44152 48252 44212 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 48608 43768 48610 43828 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 48670 44074 48672 44134 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 47770 43770 47830 43830 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 47770 44080 47830 44140 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 47660 43920 47720 43980 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 45130 43330 45190 43390 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 47660 41900 47720 41960 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 48730 41900 48790 41960 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 48730 42230 48790 42280 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 48192 41992 48252 42052 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 48192 42442 48252 42502 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 48608 42058 48610 42118 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 48670 42364 48672 42424 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 47770 42060 47830 42120 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 47770 42370 47830 42430 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 47660 42210 47720 42270 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 45130 41620 45190 41680 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 47660 52160 47720 52220 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 48730 52160 48790 52220 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 48730 52490 48790 52540 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 48192 52252 48252 52312 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 48192 52702 48252 52762 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 48608 52318 48610 52378 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 48670 52624 48672 52684 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 47770 52320 47830 52380 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 47770 52630 47830 52690 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 47660 52470 47720 52530 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 45130 51880 45190 51940 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 47660 40190 47720 40250 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 48730 40190 48790 40250 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 48730 40520 48790 40570 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 48192 40282 48252 40342 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 48192 40732 48252 40792 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 48608 40348 48610 40408 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 48670 40654 48672 40714 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 47770 40350 47830 40410 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 47770 40660 47830 40720 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 47660 40500 47720 40560 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 45130 39910 45190 39970 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 52650 64130 52710 64190 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 53720 64130 53780 64190 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 53720 64460 53780 64510 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 53182 64222 53242 64282 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 53182 64672 53242 64732 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 53598 64288 53600 64348 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 53660 64594 53662 64654 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 52760 64290 52820 64350 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 52760 64600 52820 64660 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 52650 64440 52710 64500 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 50120 63850 50180 63910 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 52650 62420 52710 62480 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 53720 62420 53780 62480 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 53720 62750 53780 62800 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 53182 62512 53242 62572 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 53182 62962 53242 63022 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 53598 62578 53600 62638 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 53660 62884 53662 62944 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 52760 62580 52820 62640 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 52760 62890 52820 62950 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 52650 62730 52710 62790 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 50120 62140 50180 62200 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 52650 60710 52710 60770 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 53720 60710 53780 60770 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 53720 61040 53780 61090 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 53182 60802 53242 60862 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 53182 61252 53242 61312 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 53598 60868 53600 60928 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 53660 61174 53662 61234 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 52760 60870 52820 60930 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 52760 61180 52820 61240 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 52650 61020 52710 61080 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 50120 60430 50180 60490 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 52650 59000 52710 59060 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 53720 59000 53780 59060 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 53720 59330 53780 59380 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 53182 59092 53242 59152 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 53182 59542 53242 59602 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 53598 59158 53600 59218 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 53660 59464 53662 59524 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 52760 59160 52820 59220 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 52760 59470 52820 59530 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 52650 59310 52710 59370 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 50120 58720 50180 58780 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 52650 57290 52710 57350 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 53720 57290 53780 57350 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 53720 57620 53780 57670 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 53182 57382 53242 57442 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 53182 57832 53242 57892 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 53598 57448 53600 57508 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 53660 57754 53662 57814 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 52760 57450 52820 57510 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 52760 57760 52820 57820 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 52650 57600 52710 57660 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 50120 57010 50180 57070 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 52650 55580 52710 55640 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 53720 55580 53780 55640 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 53720 55910 53780 55960 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 53182 55672 53242 55732 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 53182 56122 53242 56182 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 53598 55738 53600 55798 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 53660 56044 53662 56104 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 52760 55740 52820 55800 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 52760 56050 52820 56110 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 52650 55890 52710 55950 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 50120 55300 50180 55360 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 52650 65840 52710 65900 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 53720 65840 53780 65900 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 53720 66170 53780 66220 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 53182 65932 53242 65992 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 53182 66382 53242 66442 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 53598 65998 53600 66058 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 53660 66304 53662 66364 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 52760 66000 52820 66060 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 52760 66310 52820 66370 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 52650 66150 52710 66210 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 50120 65560 50180 65620 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 52650 53870 52710 53930 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 53720 53870 53780 53930 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 53720 54200 53780 54250 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 53182 53962 53242 54022 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 53182 54412 53242 54472 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 53598 54028 53600 54088 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 53660 54334 53662 54394 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 52760 54030 52820 54090 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 52760 54340 52820 54400 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 52650 54180 52710 54240 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 50120 53590 50180 53650 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 52650 50450 52710 50510 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 53720 50450 53780 50510 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 53720 50780 53780 50830 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 53182 50542 53242 50602 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 53182 50992 53242 51052 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 53598 50608 53600 50668 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 53660 50914 53662 50974 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 52760 50610 52820 50670 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 52760 50920 52820 50980 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 52650 50760 52710 50820 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 50120 50170 50180 50230 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 52650 48740 52710 48800 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 53720 48740 53780 48800 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 53720 49070 53780 49120 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 53182 48832 53242 48892 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 53182 49282 53242 49342 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 53598 48898 53600 48958 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 53660 49204 53662 49264 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 52760 48900 52820 48960 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 52760 49210 52820 49270 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 52650 49050 52710 49110 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 50120 48460 50180 48520 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 52650 47030 52710 47090 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 53720 47030 53780 47090 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 53720 47360 53780 47410 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 53182 47122 53242 47182 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 53182 47572 53242 47632 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 53598 47188 53600 47248 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 53660 47494 53662 47554 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 52760 47190 52820 47250 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 52760 47500 52820 47560 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 52650 47340 52710 47400 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 50120 46750 50180 46810 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 52650 45320 52710 45380 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 53720 45320 53780 45380 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 53720 45650 53780 45700 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 53182 45412 53242 45472 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 53182 45862 53242 45922 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 53598 45478 53600 45538 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 53660 45784 53662 45844 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 52760 45480 52820 45540 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 52760 45790 52820 45850 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 52650 45630 52710 45690 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 50120 45040 50180 45100 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 52650 43610 52710 43670 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 53720 43610 53780 43670 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 53720 43940 53780 43990 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 53182 43702 53242 43762 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 53182 44152 53242 44212 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 53598 43768 53600 43828 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 53660 44074 53662 44134 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 52760 43770 52820 43830 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 52760 44080 52820 44140 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 52650 43920 52710 43980 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 50120 43330 50180 43390 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 52650 41900 52710 41960 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 53720 41900 53780 41960 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 53720 42230 53780 42280 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 53182 41992 53242 42052 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 53182 42442 53242 42502 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 53598 42058 53600 42118 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 53660 42364 53662 42424 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 52760 42060 52820 42120 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 52760 42370 52820 42430 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 52650 42210 52710 42270 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 50120 41620 50180 41680 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 52650 52160 52710 52220 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 53720 52160 53780 52220 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 53720 52490 53780 52540 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 53182 52252 53242 52312 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 53182 52702 53242 52762 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 53598 52318 53600 52378 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 53660 52624 53662 52684 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 52760 52320 52820 52380 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 52760 52630 52820 52690 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 52650 52470 52710 52530 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 50120 51880 50180 51940 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 52650 40190 52710 40250 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 53720 40190 53780 40250 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 53720 40520 53780 40570 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 53182 40282 53242 40342 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 53182 40732 53242 40792 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 53598 40348 53600 40408 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 53660 40654 53662 40714 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 52760 40350 52820 40410 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 52760 40660 52820 40720 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 52650 40500 52710 40560 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 50120 39910 50180 39970 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 57640 64130 57700 64190 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 58710 64130 58770 64190 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 58710 64460 58770 64510 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 58172 64222 58232 64282 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 58172 64672 58232 64732 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 58588 64288 58590 64348 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 58650 64594 58652 64654 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 57750 64290 57810 64350 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 57750 64600 57810 64660 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 57640 64440 57700 64500 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 55110 63850 55170 63910 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 57640 62420 57700 62480 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 58710 62420 58770 62480 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 58710 62750 58770 62800 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 58172 62512 58232 62572 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 58172 62962 58232 63022 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 58588 62578 58590 62638 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 58650 62884 58652 62944 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 57750 62580 57810 62640 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 57750 62890 57810 62950 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 57640 62730 57700 62790 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 55110 62140 55170 62200 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 57640 60710 57700 60770 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 58710 60710 58770 60770 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 58710 61040 58770 61090 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 58172 60802 58232 60862 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 58172 61252 58232 61312 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 58588 60868 58590 60928 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 58650 61174 58652 61234 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 57750 60870 57810 60930 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 57750 61180 57810 61240 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 57640 61020 57700 61080 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 55110 60430 55170 60490 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 57640 59000 57700 59060 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 58710 59000 58770 59060 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 58710 59330 58770 59380 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 58172 59092 58232 59152 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 58172 59542 58232 59602 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 58588 59158 58590 59218 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 58650 59464 58652 59524 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 57750 59160 57810 59220 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 57750 59470 57810 59530 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 57640 59310 57700 59370 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 55110 58720 55170 58780 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 57640 57290 57700 57350 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 58710 57290 58770 57350 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 58710 57620 58770 57670 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 58172 57382 58232 57442 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 58172 57832 58232 57892 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 58588 57448 58590 57508 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 58650 57754 58652 57814 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 57750 57450 57810 57510 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 57750 57760 57810 57820 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 57640 57600 57700 57660 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 55110 57010 55170 57070 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 57640 55580 57700 55640 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 58710 55580 58770 55640 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 58710 55910 58770 55960 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 58172 55672 58232 55732 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 58172 56122 58232 56182 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 58588 55738 58590 55798 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 58650 56044 58652 56104 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 57750 55740 57810 55800 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 57750 56050 57810 56110 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 57640 55890 57700 55950 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 55110 55300 55170 55360 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 57640 65840 57700 65900 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 58710 65840 58770 65900 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 58710 66170 58770 66220 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 58172 65932 58232 65992 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 58172 66382 58232 66442 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 58588 65998 58590 66058 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 58650 66304 58652 66364 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 57750 66000 57810 66060 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 57750 66310 57810 66370 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 57640 66150 57700 66210 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 55110 65560 55170 65620 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 57640 53870 57700 53930 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 58710 53870 58770 53930 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 58710 54200 58770 54250 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 58172 53962 58232 54022 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 58172 54412 58232 54472 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 58588 54028 58590 54088 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 58650 54334 58652 54394 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 57750 54030 57810 54090 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 57750 54340 57810 54400 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 57640 54180 57700 54240 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 55110 53590 55170 53650 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 57640 50450 57700 50510 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 58710 50450 58770 50510 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 58710 50780 58770 50830 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 58172 50542 58232 50602 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 58172 50992 58232 51052 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 58588 50608 58590 50668 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 58650 50914 58652 50974 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 57750 50610 57810 50670 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 57750 50920 57810 50980 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 57640 50760 57700 50820 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 55110 50170 55170 50230 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 57640 48740 57700 48800 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 58710 48740 58770 48800 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 58710 49070 58770 49120 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 58172 48832 58232 48892 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 58172 49282 58232 49342 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 58588 48898 58590 48958 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 58650 49204 58652 49264 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 57750 48900 57810 48960 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 57750 49210 57810 49270 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 57640 49050 57700 49110 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 55110 48460 55170 48520 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 57640 47030 57700 47090 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 58710 47030 58770 47090 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 58710 47360 58770 47410 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 58172 47122 58232 47182 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 58172 47572 58232 47632 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 58588 47188 58590 47248 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 58650 47494 58652 47554 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 57750 47190 57810 47250 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 57750 47500 57810 47560 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 57640 47340 57700 47400 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 55110 46750 55170 46810 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 57640 45320 57700 45380 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 58710 45320 58770 45380 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 58710 45650 58770 45700 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 58172 45412 58232 45472 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 58172 45862 58232 45922 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 58588 45478 58590 45538 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 58650 45784 58652 45844 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 57750 45480 57810 45540 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 57750 45790 57810 45850 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 57640 45630 57700 45690 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 55110 45040 55170 45100 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 57640 43610 57700 43670 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 58710 43610 58770 43670 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 58710 43940 58770 43990 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 58172 43702 58232 43762 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 58172 44152 58232 44212 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 58588 43768 58590 43828 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 58650 44074 58652 44134 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 57750 43770 57810 43830 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 57750 44080 57810 44140 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 57640 43920 57700 43980 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 55110 43330 55170 43390 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 57640 41900 57700 41960 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 58710 41900 58770 41960 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 58710 42230 58770 42280 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 58172 41992 58232 42052 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 58172 42442 58232 42502 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 58588 42058 58590 42118 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 58650 42364 58652 42424 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 57750 42060 57810 42120 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 57750 42370 57810 42430 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 57640 42210 57700 42270 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 55110 41620 55170 41680 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 57640 52160 57700 52220 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 58710 52160 58770 52220 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 58710 52490 58770 52540 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 58172 52252 58232 52312 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 58172 52702 58232 52762 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 58588 52318 58590 52378 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 58650 52624 58652 52684 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 57750 52320 57810 52380 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 57750 52630 57810 52690 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 57640 52470 57700 52530 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 55110 51880 55170 51940 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 57640 40190 57700 40250 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 58710 40190 58770 40250 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 58710 40520 58770 40570 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 58172 40282 58232 40342 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 58172 40732 58232 40792 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 58588 40348 58590 40408 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 58650 40654 58652 40714 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 57750 40350 57810 40410 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 57750 40660 57810 40720 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 57640 40500 57700 40560 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 55110 39910 55170 39970 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 62630 64130 62690 64190 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 63700 64130 63760 64190 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 63700 64460 63760 64510 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 63162 64222 63222 64282 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 63162 64672 63222 64732 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 63578 64288 63580 64348 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 63640 64594 63642 64654 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 62740 64290 62800 64350 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 62740 64600 62800 64660 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 62630 64440 62690 64500 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 60100 63850 60160 63910 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 62630 62420 62690 62480 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 63700 62420 63760 62480 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 63700 62750 63760 62800 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 63162 62512 63222 62572 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 63162 62962 63222 63022 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 63578 62578 63580 62638 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 63640 62884 63642 62944 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 62740 62580 62800 62640 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 62740 62890 62800 62950 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 62630 62730 62690 62790 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 60100 62140 60160 62200 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 62630 60710 62690 60770 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 63700 60710 63760 60770 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 63700 61040 63760 61090 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 63162 60802 63222 60862 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 63162 61252 63222 61312 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 63578 60868 63580 60928 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 63640 61174 63642 61234 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 62740 60870 62800 60930 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 62740 61180 62800 61240 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 62630 61020 62690 61080 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 60100 60430 60160 60490 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 62630 59000 62690 59060 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 63700 59000 63760 59060 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 63700 59330 63760 59380 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 63162 59092 63222 59152 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 63162 59542 63222 59602 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 63578 59158 63580 59218 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 63640 59464 63642 59524 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 62740 59160 62800 59220 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 62740 59470 62800 59530 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 62630 59310 62690 59370 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 60100 58720 60160 58780 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 62630 57290 62690 57350 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 63700 57290 63760 57350 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 63700 57620 63760 57670 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 63162 57382 63222 57442 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 63162 57832 63222 57892 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 63578 57448 63580 57508 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 63640 57754 63642 57814 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 62740 57450 62800 57510 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 62740 57760 62800 57820 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 62630 57600 62690 57660 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 60100 57010 60160 57070 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 62630 55580 62690 55640 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 63700 55580 63760 55640 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 63700 55910 63760 55960 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 63162 55672 63222 55732 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 63162 56122 63222 56182 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 63578 55738 63580 55798 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 63640 56044 63642 56104 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 62740 55740 62800 55800 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 62740 56050 62800 56110 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 62630 55890 62690 55950 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 60100 55300 60160 55360 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 62630 65840 62690 65900 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 63700 65840 63760 65900 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 63700 66170 63760 66220 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 63162 65932 63222 65992 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 63162 66382 63222 66442 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 63578 65998 63580 66058 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 63640 66304 63642 66364 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 62740 66000 62800 66060 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 62740 66310 62800 66370 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 62630 66150 62690 66210 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 60100 65560 60160 65620 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 62630 53870 62690 53930 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 63700 53870 63760 53930 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 63700 54200 63760 54250 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 63162 53962 63222 54022 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 63162 54412 63222 54472 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 63578 54028 63580 54088 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 63640 54334 63642 54394 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 62740 54030 62800 54090 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 62740 54340 62800 54400 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 62630 54180 62690 54240 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 60100 53590 60160 53650 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 62630 50450 62690 50510 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 63700 50450 63760 50510 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 63700 50780 63760 50830 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 63162 50542 63222 50602 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 63162 50992 63222 51052 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 63578 50608 63580 50668 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 63640 50914 63642 50974 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 62740 50610 62800 50670 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 62740 50920 62800 50980 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 62630 50760 62690 50820 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 60100 50170 60160 50230 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 62630 48740 62690 48800 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 63700 48740 63760 48800 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 63700 49070 63760 49120 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 63162 48832 63222 48892 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 63162 49282 63222 49342 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 63578 48898 63580 48958 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 63640 49204 63642 49264 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 62740 48900 62800 48960 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 62740 49210 62800 49270 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 62630 49050 62690 49110 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 60100 48460 60160 48520 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 62630 47030 62690 47090 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 63700 47030 63760 47090 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 63700 47360 63760 47410 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 63162 47122 63222 47182 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 63162 47572 63222 47632 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 63578 47188 63580 47248 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 63640 47494 63642 47554 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 62740 47190 62800 47250 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 62740 47500 62800 47560 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 62630 47340 62690 47400 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 60100 46750 60160 46810 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 62630 45320 62690 45380 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 63700 45320 63760 45380 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 63700 45650 63760 45700 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 63162 45412 63222 45472 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 63162 45862 63222 45922 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 63578 45478 63580 45538 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 63640 45784 63642 45844 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 62740 45480 62800 45540 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 62740 45790 62800 45850 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 62630 45630 62690 45690 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 60100 45040 60160 45100 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 62630 43610 62690 43670 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 63700 43610 63760 43670 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 63700 43940 63760 43990 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 63162 43702 63222 43762 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 63162 44152 63222 44212 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 63578 43768 63580 43828 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 63640 44074 63642 44134 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 62740 43770 62800 43830 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 62740 44080 62800 44140 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 62630 43920 62690 43980 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 60100 43330 60160 43390 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 62630 41900 62690 41960 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 63700 41900 63760 41960 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 63700 42230 63760 42280 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 63162 41992 63222 42052 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 63162 42442 63222 42502 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 63578 42058 63580 42118 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 63640 42364 63642 42424 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 62740 42060 62800 42120 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 62740 42370 62800 42430 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 62630 42210 62690 42270 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 60100 41620 60160 41680 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 62630 52160 62690 52220 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 63700 52160 63760 52220 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 63700 52490 63760 52540 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 63162 52252 63222 52312 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 63162 52702 63222 52762 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 63578 52318 63580 52378 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 63640 52624 63642 52684 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 62740 52320 62800 52380 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 62740 52630 62800 52690 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 62630 52470 62690 52530 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 60100 51880 60160 51940 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 62630 40190 62690 40250 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 63700 40190 63760 40250 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 63700 40520 63760 40570 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 63162 40282 63222 40342 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 63162 40732 63222 40792 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 63578 40348 63580 40408 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 63640 40654 63642 40714 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 62740 40350 62800 40410 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 62740 40660 62800 40720 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 62630 40500 62690 40560 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 60100 39910 60160 39970 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 67620 64130 67680 64190 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 68690 64130 68750 64190 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 68690 64460 68750 64510 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 68152 64222 68212 64282 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 68152 64672 68212 64732 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 68568 64288 68570 64348 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 68630 64594 68632 64654 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 67730 64290 67790 64350 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 67730 64600 67790 64660 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 67620 64440 67680 64500 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 65090 63850 65150 63910 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 67620 62420 67680 62480 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 68690 62420 68750 62480 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 68690 62750 68750 62800 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 68152 62512 68212 62572 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 68152 62962 68212 63022 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 68568 62578 68570 62638 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 68630 62884 68632 62944 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 67730 62580 67790 62640 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 67730 62890 67790 62950 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 67620 62730 67680 62790 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 65090 62140 65150 62200 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 67620 60710 67680 60770 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 68690 60710 68750 60770 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 68690 61040 68750 61090 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 68152 60802 68212 60862 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 68152 61252 68212 61312 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 68568 60868 68570 60928 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 68630 61174 68632 61234 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 67730 60870 67790 60930 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 67730 61180 67790 61240 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 67620 61020 67680 61080 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 65090 60430 65150 60490 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 67620 59000 67680 59060 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 68690 59000 68750 59060 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 68690 59330 68750 59380 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 68152 59092 68212 59152 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 68152 59542 68212 59602 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 68568 59158 68570 59218 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 68630 59464 68632 59524 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 67730 59160 67790 59220 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 67730 59470 67790 59530 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 67620 59310 67680 59370 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 65090 58720 65150 58780 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 67620 57290 67680 57350 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 68690 57290 68750 57350 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 68690 57620 68750 57670 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 68152 57382 68212 57442 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 68152 57832 68212 57892 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 68568 57448 68570 57508 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 68630 57754 68632 57814 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 67730 57450 67790 57510 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 67730 57760 67790 57820 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 67620 57600 67680 57660 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 65090 57010 65150 57070 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 67620 55580 67680 55640 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 68690 55580 68750 55640 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 68690 55910 68750 55960 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 68152 55672 68212 55732 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 68152 56122 68212 56182 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 68568 55738 68570 55798 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 68630 56044 68632 56104 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 67730 55740 67790 55800 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 67730 56050 67790 56110 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 67620 55890 67680 55950 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 65090 55300 65150 55360 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 67620 65840 67680 65900 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 68690 65840 68750 65900 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 68690 66170 68750 66220 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 68152 65932 68212 65992 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 68152 66382 68212 66442 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 68568 65998 68570 66058 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 68630 66304 68632 66364 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 67730 66000 67790 66060 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 67730 66310 67790 66370 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 67620 66150 67680 66210 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 65090 65560 65150 65620 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 67620 53870 67680 53930 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 68690 53870 68750 53930 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 68690 54200 68750 54250 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 68152 53962 68212 54022 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 68152 54412 68212 54472 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 68568 54028 68570 54088 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 68630 54334 68632 54394 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 67730 54030 67790 54090 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 67730 54340 67790 54400 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 67620 54180 67680 54240 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 65090 53590 65150 53650 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 67620 50450 67680 50510 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 68690 50450 68750 50510 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 68690 50780 68750 50830 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 68152 50542 68212 50602 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 68152 50992 68212 51052 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 68568 50608 68570 50668 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 68630 50914 68632 50974 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 67730 50610 67790 50670 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 67730 50920 67790 50980 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 67620 50760 67680 50820 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 65090 50170 65150 50230 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 67620 48740 67680 48800 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 68690 48740 68750 48800 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 68690 49070 68750 49120 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 68152 48832 68212 48892 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 68152 49282 68212 49342 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 68568 48898 68570 48958 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 68630 49204 68632 49264 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 67730 48900 67790 48960 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 67730 49210 67790 49270 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 67620 49050 67680 49110 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 65090 48460 65150 48520 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 67620 47030 67680 47090 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 68690 47030 68750 47090 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 68690 47360 68750 47410 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 68152 47122 68212 47182 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 68152 47572 68212 47632 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 68568 47188 68570 47248 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 68630 47494 68632 47554 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 67730 47190 67790 47250 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 67730 47500 67790 47560 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 67620 47340 67680 47400 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 65090 46750 65150 46810 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 67620 45320 67680 45380 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 68690 45320 68750 45380 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 68690 45650 68750 45700 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 68152 45412 68212 45472 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 68152 45862 68212 45922 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 68568 45478 68570 45538 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 68630 45784 68632 45844 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 67730 45480 67790 45540 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 67730 45790 67790 45850 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 67620 45630 67680 45690 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 65090 45040 65150 45100 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 67620 43610 67680 43670 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 68690 43610 68750 43670 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 68690 43940 68750 43990 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 68152 43702 68212 43762 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 68152 44152 68212 44212 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 68568 43768 68570 43828 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 68630 44074 68632 44134 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 67730 43770 67790 43830 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 67730 44080 67790 44140 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 67620 43920 67680 43980 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 65090 43330 65150 43390 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 67620 41900 67680 41960 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 68690 41900 68750 41960 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 68690 42230 68750 42280 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 68152 41992 68212 42052 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 68152 42442 68212 42502 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 68568 42058 68570 42118 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 68630 42364 68632 42424 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 67730 42060 67790 42120 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 67730 42370 67790 42430 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 67620 42210 67680 42270 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 65090 41620 65150 41680 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 67620 52160 67680 52220 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 68690 52160 68750 52220 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 68690 52490 68750 52540 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 68152 52252 68212 52312 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 68152 52702 68212 52762 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 68568 52318 68570 52378 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 68630 52624 68632 52684 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 67730 52320 67790 52380 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 67730 52630 67790 52690 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 67620 52470 67680 52530 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 65090 51880 65150 51940 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 67620 40190 67680 40250 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 68690 40190 68750 40250 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 68690 40520 68750 40570 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 68152 40282 68212 40342 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 68152 40732 68212 40792 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 68568 40348 68570 40408 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 68630 40654 68632 40714 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 67730 40350 67790 40410 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 67730 40660 67790 40720 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 67620 40500 67680 40560 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 65090 39910 65150 39970 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 72610 64130 72670 64190 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 73680 64130 73740 64190 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 73680 64460 73740 64510 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 73142 64222 73202 64282 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 73142 64672 73202 64732 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 73558 64288 73560 64348 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 73620 64594 73622 64654 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 72720 64290 72780 64350 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 72720 64600 72780 64660 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 72610 64440 72670 64500 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 70080 63850 70140 63910 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 72610 62420 72670 62480 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 73680 62420 73740 62480 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 73680 62750 73740 62800 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 73142 62512 73202 62572 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 73142 62962 73202 63022 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 73558 62578 73560 62638 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 73620 62884 73622 62944 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 72720 62580 72780 62640 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 72720 62890 72780 62950 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 72610 62730 72670 62790 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 70080 62140 70140 62200 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 72610 60710 72670 60770 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 73680 60710 73740 60770 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 73680 61040 73740 61090 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 73142 60802 73202 60862 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 73142 61252 73202 61312 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 73558 60868 73560 60928 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 73620 61174 73622 61234 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 72720 60870 72780 60930 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 72720 61180 72780 61240 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 72610 61020 72670 61080 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 70080 60430 70140 60490 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 72610 59000 72670 59060 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 73680 59000 73740 59060 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 73680 59330 73740 59380 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 73142 59092 73202 59152 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 73142 59542 73202 59602 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 73558 59158 73560 59218 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 73620 59464 73622 59524 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 72720 59160 72780 59220 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 72720 59470 72780 59530 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 72610 59310 72670 59370 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 70080 58720 70140 58780 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 72610 57290 72670 57350 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 73680 57290 73740 57350 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 73680 57620 73740 57670 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 73142 57382 73202 57442 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 73142 57832 73202 57892 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 73558 57448 73560 57508 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 73620 57754 73622 57814 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 72720 57450 72780 57510 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 72720 57760 72780 57820 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 72610 57600 72670 57660 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 70080 57010 70140 57070 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 72610 55580 72670 55640 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 73680 55580 73740 55640 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 73680 55910 73740 55960 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 73142 55672 73202 55732 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 73142 56122 73202 56182 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 73558 55738 73560 55798 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 73620 56044 73622 56104 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 72720 55740 72780 55800 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 72720 56050 72780 56110 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 72610 55890 72670 55950 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 70080 55300 70140 55360 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 72610 65840 72670 65900 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 73680 65840 73740 65900 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 73680 66170 73740 66220 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 73142 65932 73202 65992 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 73142 66382 73202 66442 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 73558 65998 73560 66058 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 73620 66304 73622 66364 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 72720 66000 72780 66060 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 72720 66310 72780 66370 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 72610 66150 72670 66210 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 70080 65560 70140 65620 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 72610 53870 72670 53930 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 73680 53870 73740 53930 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 73680 54200 73740 54250 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 73142 53962 73202 54022 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 73142 54412 73202 54472 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 73558 54028 73560 54088 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 73620 54334 73622 54394 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 72720 54030 72780 54090 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 72720 54340 72780 54400 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 72610 54180 72670 54240 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 70080 53590 70140 53650 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 72610 50450 72670 50510 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 73680 50450 73740 50510 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 73680 50780 73740 50830 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 73142 50542 73202 50602 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 73142 50992 73202 51052 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 73558 50608 73560 50668 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 73620 50914 73622 50974 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 72720 50610 72780 50670 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 72720 50920 72780 50980 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 72610 50760 72670 50820 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 70080 50170 70140 50230 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 72610 48740 72670 48800 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 73680 48740 73740 48800 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 73680 49070 73740 49120 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 73142 48832 73202 48892 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 73142 49282 73202 49342 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 73558 48898 73560 48958 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 73620 49204 73622 49264 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 72720 48900 72780 48960 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 72720 49210 72780 49270 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 72610 49050 72670 49110 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 70080 48460 70140 48520 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 72610 47030 72670 47090 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 73680 47030 73740 47090 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 73680 47360 73740 47410 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 73142 47122 73202 47182 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 73142 47572 73202 47632 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 73558 47188 73560 47248 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 73620 47494 73622 47554 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 72720 47190 72780 47250 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 72720 47500 72780 47560 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 72610 47340 72670 47400 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 70080 46750 70140 46810 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 72610 45320 72670 45380 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 73680 45320 73740 45380 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 73680 45650 73740 45700 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 73142 45412 73202 45472 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 73142 45862 73202 45922 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 73558 45478 73560 45538 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 73620 45784 73622 45844 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 72720 45480 72780 45540 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 72720 45790 72780 45850 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 72610 45630 72670 45690 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 70080 45040 70140 45100 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 72610 43610 72670 43670 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 73680 43610 73740 43670 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 73680 43940 73740 43990 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 73142 43702 73202 43762 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 73142 44152 73202 44212 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 73558 43768 73560 43828 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 73620 44074 73622 44134 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 72720 43770 72780 43830 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 72720 44080 72780 44140 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 72610 43920 72670 43980 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 70080 43330 70140 43390 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 72610 41900 72670 41960 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 73680 41900 73740 41960 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 73680 42230 73740 42280 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 73142 41992 73202 42052 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 73142 42442 73202 42502 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 73558 42058 73560 42118 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 73620 42364 73622 42424 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 72720 42060 72780 42120 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 72720 42370 72780 42430 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 72610 42210 72670 42270 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 70080 41620 70140 41680 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 72610 52160 72670 52220 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 73680 52160 73740 52220 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 73680 52490 73740 52540 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 73142 52252 73202 52312 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 73142 52702 73202 52762 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 73558 52318 73560 52378 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 73620 52624 73622 52684 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 72720 52320 72780 52380 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 72720 52630 72780 52690 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 72610 52470 72670 52530 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 70080 51880 70140 51940 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 72610 40190 72670 40250 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 73680 40190 73740 40250 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 73680 40520 73740 40570 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 73142 40282 73202 40342 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 73142 40732 73202 40792 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 73558 40348 73560 40408 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 73620 40654 73622 40714 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 72720 40350 72780 40410 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 72720 40660 72780 40720 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 72610 40500 72670 40560 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 70080 39910 70140 39970 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 77600 64130 77660 64190 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 78670 64130 78730 64190 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 78670 64460 78730 64510 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 78132 64222 78192 64282 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 78132 64672 78192 64732 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 78548 64288 78550 64348 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 78610 64594 78612 64654 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 77710 64290 77770 64350 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 77710 64600 77770 64660 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 77600 64440 77660 64500 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 75070 63850 75130 63910 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 77600 62420 77660 62480 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 78670 62420 78730 62480 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 78670 62750 78730 62800 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 78132 62512 78192 62572 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 78132 62962 78192 63022 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 78548 62578 78550 62638 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 78610 62884 78612 62944 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 77710 62580 77770 62640 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 77710 62890 77770 62950 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 77600 62730 77660 62790 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 75070 62140 75130 62200 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 77600 60710 77660 60770 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 78670 60710 78730 60770 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 78670 61040 78730 61090 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 78132 60802 78192 60862 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 78132 61252 78192 61312 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 78548 60868 78550 60928 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 78610 61174 78612 61234 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 77710 60870 77770 60930 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 77710 61180 77770 61240 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 77600 61020 77660 61080 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 75070 60430 75130 60490 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 77600 59000 77660 59060 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 78670 59000 78730 59060 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 78670 59330 78730 59380 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 78132 59092 78192 59152 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 78132 59542 78192 59602 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 78548 59158 78550 59218 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 78610 59464 78612 59524 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 77710 59160 77770 59220 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 77710 59470 77770 59530 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 77600 59310 77660 59370 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 75070 58720 75130 58780 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 77600 57290 77660 57350 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 78670 57290 78730 57350 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 78670 57620 78730 57670 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 78132 57382 78192 57442 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 78132 57832 78192 57892 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 78548 57448 78550 57508 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 78610 57754 78612 57814 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 77710 57450 77770 57510 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 77710 57760 77770 57820 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 77600 57600 77660 57660 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 75070 57010 75130 57070 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 77600 55580 77660 55640 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 78670 55580 78730 55640 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 78670 55910 78730 55960 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 78132 55672 78192 55732 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 78132 56122 78192 56182 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 78548 55738 78550 55798 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 78610 56044 78612 56104 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 77710 55740 77770 55800 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 77710 56050 77770 56110 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 77600 55890 77660 55950 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 75070 55300 75130 55360 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 77600 65840 77660 65900 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 78670 65840 78730 65900 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 78670 66170 78730 66220 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 78132 65932 78192 65992 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 78132 66382 78192 66442 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 78548 65998 78550 66058 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 78610 66304 78612 66364 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 77710 66000 77770 66060 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 77710 66310 77770 66370 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 77600 66150 77660 66210 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 75070 65560 75130 65620 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 77600 53870 77660 53930 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 78670 53870 78730 53930 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 78670 54200 78730 54250 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 78132 53962 78192 54022 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 78132 54412 78192 54472 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 78548 54028 78550 54088 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 78610 54334 78612 54394 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 77710 54030 77770 54090 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 77710 54340 77770 54400 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 77600 54180 77660 54240 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 75070 53590 75130 53650 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 77600 50450 77660 50510 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 78670 50450 78730 50510 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 78670 50780 78730 50830 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 78132 50542 78192 50602 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 78132 50992 78192 51052 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 78548 50608 78550 50668 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 78610 50914 78612 50974 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 77710 50610 77770 50670 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 77710 50920 77770 50980 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 77600 50760 77660 50820 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 75070 50170 75130 50230 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 77600 48740 77660 48800 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 78670 48740 78730 48800 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 78670 49070 78730 49120 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 78132 48832 78192 48892 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 78132 49282 78192 49342 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 78548 48898 78550 48958 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 78610 49204 78612 49264 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 77710 48900 77770 48960 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 77710 49210 77770 49270 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 77600 49050 77660 49110 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 75070 48460 75130 48520 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 77600 47030 77660 47090 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 78670 47030 78730 47090 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 78670 47360 78730 47410 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 78132 47122 78192 47182 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 78132 47572 78192 47632 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 78548 47188 78550 47248 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 78610 47494 78612 47554 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 77710 47190 77770 47250 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 77710 47500 77770 47560 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 77600 47340 77660 47400 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 75070 46750 75130 46810 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 77600 45320 77660 45380 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 78670 45320 78730 45380 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 78670 45650 78730 45700 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 78132 45412 78192 45472 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 78132 45862 78192 45922 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 78548 45478 78550 45538 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 78610 45784 78612 45844 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 77710 45480 77770 45540 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 77710 45790 77770 45850 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 77600 45630 77660 45690 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 75070 45040 75130 45100 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 77600 43610 77660 43670 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 78670 43610 78730 43670 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 78670 43940 78730 43990 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 78132 43702 78192 43762 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 78132 44152 78192 44212 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 78548 43768 78550 43828 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 78610 44074 78612 44134 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 77710 43770 77770 43830 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 77710 44080 77770 44140 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 77600 43920 77660 43980 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 75070 43330 75130 43390 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 77600 41900 77660 41960 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 78670 41900 78730 41960 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 78670 42230 78730 42280 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 78132 41992 78192 42052 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 78132 42442 78192 42502 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 78548 42058 78550 42118 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 78610 42364 78612 42424 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 77710 42060 77770 42120 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 77710 42370 77770 42430 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 77600 42210 77660 42270 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 75070 41620 75130 41680 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 77600 52160 77660 52220 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 78670 52160 78730 52220 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 78670 52490 78730 52540 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 78132 52252 78192 52312 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 78132 52702 78192 52762 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 78548 52318 78550 52378 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 78610 52624 78612 52684 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 77710 52320 77770 52380 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 77710 52630 77770 52690 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 77600 52470 77660 52530 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 75070 51880 75130 51940 0 FreeSans 256 270 0 0 com_x
port 0 nsew
flabel metal1 77600 40190 77660 40250 0 FreeSans 256 270 0 0 sub
port 6 nsew
flabel metal1 78670 40190 78730 40250 0 FreeSans 256 270 0 0 Vdd
port 3 nsew
flabel metal1 78670 40520 78730 40570 0 FreeSans 256 270 0 0 Vdd
port 7 nsew
flabel metal1 78132 40282 78192 40342 0 FreeSans 256 270 0 0 Vin
port 5 nsew
flabel metal1 78132 40732 78192 40792 0 FreeSans 256 270 0 0 GND
port 9 nsew
flabel metal1 78548 40348 78550 40408 0 FreeSans 256 270 0 0 phi1_n
port 4 nsew
flabel metal1 78610 40654 78612 40714 0 FreeSans 256 270 0 0 phi2_n
port 10 nsew
flabel via1 77710 40350 77770 40410 0 FreeSans 256 270 0 0 phi1
port 2 nsew
flabel via1 77710 40660 77770 40720 0 FreeSans 256 270 0 0 phi2
port 8 nsew
flabel metal1 77600 40500 77660 40560 0 FreeSans 256 270 0 0 sub
port 1 nsew
flabel metal4 75070 39910 75130 39970 0 FreeSans 256 270 0 0 com_x
port 0 nsew
<< end >>
