magic
tech sky130A
timestamp 1730537705
<< metal1 >>
rect 2075 15450 2080 15465
rect -30 15435 2080 15450
rect 2110 15450 2115 15465
rect 4570 15450 4575 15465
rect 2110 15435 4575 15450
rect 4605 15450 4610 15465
rect 7065 15450 7070 15465
rect 4605 15435 7070 15450
rect 7100 15450 7105 15465
rect 9560 15450 9565 15465
rect 7100 15435 9565 15450
rect 9595 15450 9600 15465
rect 12055 15450 12060 15465
rect 9595 15435 12060 15450
rect 12090 15450 12095 15465
rect 14550 15450 14555 15465
rect 12090 15435 14555 15450
rect 14585 15450 14590 15465
rect 17045 15450 17050 15465
rect 14585 15435 17050 15450
rect 17080 15450 17085 15465
rect 19540 15450 19545 15465
rect 17080 15435 19545 15450
rect 19575 15450 19580 15465
rect 22035 15450 22040 15465
rect 19575 15435 22040 15450
rect 22070 15450 22075 15465
rect 24530 15450 24535 15465
rect 22070 15435 24535 15450
rect 24565 15450 24570 15465
rect 27025 15450 27030 15465
rect 24565 15435 27030 15450
rect 27060 15450 27065 15465
rect 29520 15450 29525 15465
rect 27060 15435 29525 15450
rect 29555 15450 29560 15465
rect 32015 15450 32020 15465
rect 29555 15435 32020 15450
rect 32050 15450 32055 15465
rect 34510 15450 34515 15465
rect 32050 15435 34515 15450
rect 34545 15450 34550 15465
rect 37005 15450 37010 15465
rect 34545 15435 37010 15450
rect 37040 15450 37045 15465
rect 39500 15450 39505 15465
rect 37040 15435 39505 15450
rect 39535 15450 39540 15465
rect 39535 15435 39850 15450
rect 64 15433 117 15435
rect 1210 15380 1240 15400
rect 2045 15380 2050 15395
rect -30 15365 2050 15380
rect 2080 15380 2085 15395
rect 3705 15380 3735 15400
rect 4540 15380 4545 15395
rect 2080 15365 4545 15380
rect 4575 15380 4580 15395
rect 6200 15380 6230 15400
rect 7035 15380 7040 15395
rect 4575 15365 7040 15380
rect 7070 15380 7075 15395
rect 8695 15380 8725 15400
rect 9530 15380 9535 15395
rect 7070 15365 9535 15380
rect 9565 15380 9570 15395
rect 11190 15380 11220 15400
rect 12025 15380 12030 15395
rect 9565 15365 12030 15380
rect 12060 15380 12065 15395
rect 13685 15380 13715 15400
rect 14520 15380 14525 15395
rect 12060 15365 14525 15380
rect 14555 15380 14560 15395
rect 16180 15380 16210 15400
rect 17015 15380 17020 15395
rect 14555 15365 17020 15380
rect 17050 15380 17055 15395
rect 18675 15380 18705 15400
rect 19510 15380 19515 15395
rect 17050 15365 19515 15380
rect 19545 15380 19550 15395
rect 21170 15380 21200 15400
rect 22005 15380 22010 15395
rect 19545 15365 22010 15380
rect 22040 15380 22045 15395
rect 23665 15380 23695 15400
rect 24500 15380 24505 15395
rect 22040 15365 24505 15380
rect 24535 15380 24540 15395
rect 26160 15380 26190 15400
rect 26995 15380 27000 15395
rect 24535 15365 27000 15380
rect 27030 15380 27035 15395
rect 28655 15380 28685 15400
rect 29490 15380 29495 15395
rect 27030 15365 29495 15380
rect 29525 15380 29530 15395
rect 31150 15380 31180 15400
rect 31985 15380 31990 15395
rect 29525 15365 31990 15380
rect 32020 15380 32025 15395
rect 33645 15380 33675 15400
rect 34480 15380 34485 15395
rect 32020 15365 34485 15380
rect 34515 15380 34520 15395
rect 36140 15380 36170 15400
rect 36975 15380 36980 15395
rect 34515 15365 36980 15380
rect 37010 15380 37015 15395
rect 38635 15380 38665 15400
rect 39470 15380 39475 15395
rect 37010 15365 39475 15380
rect 39505 15380 39510 15395
rect 39505 15365 39850 15380
rect 65 15364 118 15365
rect 7155 15310 7160 15325
rect -30 15295 7160 15310
rect 7190 15310 7195 15325
rect 9650 15310 9655 15325
rect 7190 15295 9655 15310
rect 9685 15310 9690 15325
rect 12145 15310 12150 15325
rect 9685 15295 12150 15310
rect 12180 15310 12185 15325
rect 14640 15310 14645 15325
rect 12180 15295 14645 15310
rect 14675 15310 14680 15325
rect 17135 15310 17140 15325
rect 14675 15295 17140 15310
rect 17170 15310 17175 15325
rect 19630 15310 19635 15325
rect 17170 15295 19635 15310
rect 19665 15310 19670 15325
rect 22125 15310 22130 15325
rect 19665 15295 22130 15310
rect 22160 15310 22165 15325
rect 24620 15310 24625 15325
rect 22160 15295 24625 15310
rect 24655 15310 24660 15325
rect 27115 15310 27120 15325
rect 24655 15295 27120 15310
rect 27150 15310 27155 15325
rect 29610 15310 29615 15325
rect 27150 15295 29615 15310
rect 29645 15310 29650 15325
rect 32105 15310 32110 15325
rect 29645 15295 32110 15310
rect 32140 15310 32145 15325
rect 34600 15310 34605 15325
rect 32140 15295 34605 15310
rect 34635 15310 34640 15325
rect 34635 15295 39850 15310
rect 63 15293 116 15295
rect 6110 15240 6140 15260
rect 7125 15240 7130 15255
rect -30 15225 7130 15240
rect 7160 15240 7165 15255
rect 8605 15240 8635 15260
rect 9620 15240 9625 15255
rect 7160 15225 9625 15240
rect 9655 15240 9660 15255
rect 11100 15240 11130 15260
rect 12115 15240 12120 15255
rect 9655 15225 12120 15240
rect 12150 15240 12155 15255
rect 13595 15240 13625 15260
rect 14610 15240 14615 15255
rect 12150 15225 14615 15240
rect 14645 15240 14650 15255
rect 16090 15240 16120 15260
rect 17105 15240 17110 15255
rect 14645 15225 17110 15240
rect 17140 15240 17145 15255
rect 18585 15240 18615 15260
rect 19600 15240 19605 15255
rect 17140 15225 19605 15240
rect 19635 15240 19640 15255
rect 21080 15240 21110 15260
rect 22095 15240 22100 15255
rect 19635 15225 22100 15240
rect 22130 15240 22135 15255
rect 23575 15240 23605 15260
rect 24590 15240 24595 15255
rect 22130 15225 24595 15240
rect 24625 15240 24630 15255
rect 26070 15240 26100 15260
rect 27085 15240 27090 15255
rect 24625 15225 27090 15240
rect 27120 15240 27125 15255
rect 28565 15240 28595 15260
rect 29580 15240 29585 15255
rect 27120 15225 29585 15240
rect 29615 15240 29620 15255
rect 31060 15240 31090 15260
rect 32075 15240 32080 15255
rect 29615 15225 32080 15240
rect 32110 15240 32115 15255
rect 33555 15240 33585 15260
rect 34570 15240 34575 15255
rect 32110 15225 34575 15240
rect 34605 15240 34610 15255
rect 34605 15225 39850 15240
rect 61 15223 114 15225
rect 12325 15170 12330 15185
rect -30 15155 12330 15170
rect 12360 15170 12365 15185
rect 14820 15170 14825 15185
rect 12360 15155 14825 15170
rect 14855 15170 14860 15185
rect 17225 15170 17230 15185
rect 14855 15155 17230 15170
rect 17260 15170 17265 15185
rect 19720 15170 19725 15185
rect 17260 15155 19725 15170
rect 19755 15170 19760 15185
rect 22215 15170 22220 15185
rect 19755 15155 22220 15170
rect 22250 15170 22255 15185
rect 24710 15170 24715 15185
rect 22250 15155 24715 15170
rect 24745 15170 24750 15185
rect 27295 15170 27300 15185
rect 24745 15155 27300 15170
rect 27330 15170 27335 15185
rect 29790 15170 29795 15185
rect 27330 15155 29795 15170
rect 29825 15170 29830 15185
rect 29825 15155 39850 15170
rect 59 15154 112 15155
rect 10920 15100 10950 15120
rect 12295 15100 12300 15115
rect -30 15085 12300 15100
rect 12330 15100 12335 15115
rect 13415 15100 13445 15120
rect 14790 15100 14795 15115
rect 12330 15085 14795 15100
rect 14825 15100 14830 15115
rect 16000 15100 16030 15120
rect 17195 15100 17200 15115
rect 14825 15085 17200 15100
rect 17230 15100 17235 15115
rect 18495 15100 18525 15120
rect 19690 15100 19695 15115
rect 17230 15085 19695 15100
rect 19725 15100 19730 15115
rect 20990 15100 21020 15120
rect 22185 15100 22190 15115
rect 19725 15085 22190 15100
rect 22220 15100 22225 15115
rect 23485 15100 23515 15120
rect 24680 15100 24685 15115
rect 22220 15085 24685 15100
rect 24715 15100 24720 15115
rect 25890 15100 25920 15120
rect 27265 15100 27270 15115
rect 24715 15085 27270 15100
rect 27300 15100 27305 15115
rect 28385 15100 28415 15120
rect 29760 15100 29765 15115
rect 27300 15085 29765 15100
rect 29795 15100 29800 15115
rect 29795 15085 39850 15100
rect 59 15084 112 15085
rect 12235 15030 12240 15045
rect -30 15015 12240 15030
rect 12270 15030 12275 15045
rect 14730 15030 14735 15045
rect 12270 15015 14735 15030
rect 14765 15030 14770 15045
rect 17315 15030 17320 15045
rect 14765 15015 17320 15030
rect 17350 15030 17355 15045
rect 19810 15030 19815 15045
rect 17350 15015 19815 15030
rect 19845 15030 19850 15045
rect 22305 15030 22310 15045
rect 19845 15015 22310 15030
rect 22340 15030 22345 15045
rect 24800 15030 24805 15045
rect 22340 15015 24805 15030
rect 24835 15030 24840 15045
rect 27205 15030 27210 15045
rect 24835 15015 27210 15030
rect 27240 15030 27245 15045
rect 29700 15030 29705 15045
rect 27240 15015 29705 15030
rect 29735 15030 29740 15045
rect 29735 15015 39850 15030
rect 58 15013 111 15015
rect 11010 14960 11040 14980
rect 12205 14960 12210 14975
rect -30 14945 12210 14960
rect 12240 14960 12245 14975
rect 13505 14960 13535 14980
rect 14700 14960 14705 14975
rect 12240 14945 14705 14960
rect 14735 14960 14740 14975
rect 15910 14960 15940 14980
rect 17285 14960 17290 14975
rect 14735 14945 17290 14960
rect 17320 14960 17325 14975
rect 18405 14960 18435 14980
rect 19780 14960 19785 14975
rect 17320 14945 19785 14960
rect 19815 14960 19820 14975
rect 20900 14960 20930 14980
rect 22275 14960 22280 14975
rect 19815 14945 22280 14960
rect 22310 14960 22315 14975
rect 23395 14960 23425 14980
rect 24770 14960 24775 14975
rect 22310 14945 24775 14960
rect 24805 14960 24810 14975
rect 25980 14960 26010 14980
rect 27175 14960 27180 14975
rect 24805 14945 27180 14960
rect 27210 14960 27215 14975
rect 28475 14960 28505 14980
rect 29670 14960 29675 14975
rect 27210 14945 29675 14960
rect 29705 14960 29710 14975
rect 29705 14945 39850 14960
rect 55 14943 108 14945
rect 17495 14890 17500 14905
rect -30 14875 17500 14890
rect 17530 14890 17535 14905
rect 19900 14890 19905 14905
rect 17530 14875 19905 14890
rect 19935 14890 19940 14905
rect 22395 14890 22400 14905
rect 19935 14875 22400 14890
rect 22430 14890 22435 14905
rect 24980 14890 24985 14905
rect 22430 14875 24985 14890
rect 25015 14890 25020 14905
rect 25015 14875 39850 14890
rect 58 14873 111 14875
rect 15730 14820 15760 14840
rect 17465 14820 17470 14835
rect -30 14805 17470 14820
rect 17500 14820 17505 14835
rect 18315 14820 18345 14840
rect 19870 14820 19875 14835
rect 17500 14805 19875 14820
rect 19905 14820 19910 14835
rect 20810 14820 20840 14840
rect 22365 14820 22370 14835
rect 19905 14805 22370 14820
rect 22400 14820 22405 14835
rect 23215 14820 23245 14840
rect 24950 14820 24955 14835
rect 22400 14805 24955 14820
rect 24985 14820 24990 14835
rect 24985 14805 39850 14820
rect 58 14804 111 14805
rect 17405 14750 17410 14765
rect -30 14735 17410 14750
rect 17440 14750 17445 14765
rect 24890 14750 24895 14765
rect 17440 14735 24895 14750
rect 24925 14750 24930 14765
rect 24925 14735 39850 14750
rect 61 14733 114 14735
rect 15820 14680 15850 14700
rect 17375 14680 17380 14695
rect -30 14665 17380 14680
rect 17410 14680 17415 14695
rect 23305 14680 23335 14700
rect 24860 14680 24865 14695
rect 17410 14665 24865 14680
rect 24895 14680 24900 14695
rect 24895 14665 39850 14680
rect 63 14664 116 14665
rect 19990 14610 19995 14625
rect -30 14595 19995 14610
rect 20025 14610 20030 14625
rect 22575 14610 22580 14625
rect 20025 14595 22580 14610
rect 22610 14610 22615 14625
rect 22610 14595 39850 14610
rect 58 14593 111 14595
rect 18225 14540 18255 14560
rect 19960 14540 19965 14555
rect -30 14525 19965 14540
rect 19995 14540 20000 14555
rect 22545 14540 22550 14555
rect 19995 14525 22550 14540
rect 22580 14540 22585 14555
rect 22580 14525 39850 14540
rect 62 14523 115 14525
rect 22500 14470 22505 14485
rect -30 14455 22505 14470
rect 22535 14470 22540 14485
rect 22535 14455 39850 14470
rect 65 14453 118 14455
rect 22455 14400 22460 14415
rect -30 14385 22460 14400
rect 22490 14400 22495 14415
rect 22490 14385 39850 14400
rect 68 14383 121 14385
rect 18105 14330 18135 14350
rect 20080 14330 20085 14345
rect -30 14315 20085 14330
rect 20115 14330 20120 14345
rect 20115 14315 39850 14330
rect 67 14314 120 14315
rect 18135 14260 18165 14280
rect 20045 14260 20050 14275
rect -30 14245 20050 14260
rect 20080 14260 20085 14275
rect 20080 14245 39850 14260
rect 67 14190 120 14191
rect 1930 14190 1935 14205
rect -30 14175 1935 14190
rect 1965 14190 1970 14205
rect 4425 14190 4430 14205
rect 1965 14175 4430 14190
rect 4460 14190 4465 14205
rect 6920 14190 6925 14205
rect 4460 14175 6925 14190
rect 6955 14190 6960 14205
rect 9415 14190 9420 14205
rect 6955 14175 9420 14190
rect 9450 14190 9455 14205
rect 11910 14190 11915 14205
rect 9450 14175 11915 14190
rect 11945 14190 11950 14205
rect 14405 14190 14410 14205
rect 11945 14175 14410 14190
rect 14440 14190 14445 14205
rect 16900 14190 16905 14205
rect 14440 14175 16905 14190
rect 16935 14190 16940 14205
rect 19395 14190 19400 14205
rect 16935 14175 19400 14190
rect 19430 14190 19435 14205
rect 21890 14190 21895 14205
rect 19430 14175 21895 14190
rect 21925 14190 21930 14205
rect 24385 14190 24390 14205
rect 21925 14175 24390 14190
rect 24420 14190 24425 14205
rect 26880 14190 26885 14205
rect 24420 14175 26885 14190
rect 26915 14190 26920 14205
rect 29375 14190 29380 14205
rect 26915 14175 29380 14190
rect 29410 14190 29415 14205
rect 31870 14190 31875 14205
rect 29410 14175 31875 14190
rect 31905 14190 31910 14205
rect 34365 14190 34370 14205
rect 31905 14175 34370 14190
rect 34400 14190 34405 14205
rect 36860 14190 36865 14205
rect 34400 14175 36865 14190
rect 36895 14190 36900 14205
rect 39355 14190 39360 14205
rect 36895 14175 39360 14190
rect 39390 14190 39395 14205
rect 39390 14175 39850 14190
rect 66 14174 119 14175
rect 67 14120 120 14121
rect -30 14105 39850 14120
rect 68 14103 121 14105
rect 1175 13940 1205 13945
rect 1205 13910 1305 13920
rect 1175 13905 1305 13910
rect 1290 13680 1305 13905
rect 1855 13715 1895 13720
rect 1320 13685 1325 13715
rect 1355 13685 1360 13715
rect 1320 13680 1360 13685
rect 1855 13685 1860 13715
rect 1890 13685 1895 13715
rect 1855 13680 1895 13685
rect 1910 13680 1925 14105
rect 2085 13940 2115 13945
rect 1985 13910 2085 13920
rect 1985 13905 2115 13910
rect 3670 13940 3700 13945
rect 3700 13910 3800 13920
rect 3670 13905 3800 13910
rect 1940 13715 1970 13720
rect 1940 13680 1970 13685
rect 1985 13680 2000 13905
rect 3785 13680 3800 13905
rect 4350 13715 4390 13720
rect 3815 13685 3820 13715
rect 3850 13685 3855 13715
rect 3815 13680 3855 13685
rect 4350 13685 4355 13715
rect 4385 13685 4390 13715
rect 4350 13680 4390 13685
rect 4405 13680 4420 14105
rect 4580 13940 4610 13945
rect 4480 13910 4580 13920
rect 6165 13940 6195 13945
rect 4480 13905 4610 13910
rect 6075 13910 6105 13915
rect 4435 13715 4465 13720
rect 4435 13680 4465 13685
rect 4480 13680 4495 13905
rect 6195 13910 6295 13920
rect 6165 13905 6295 13910
rect 6105 13880 6235 13890
rect 6075 13875 6235 13880
rect 6220 13680 6235 13875
rect 6280 13680 6295 13905
rect 6845 13715 6885 13720
rect 6310 13685 6315 13715
rect 6345 13685 6350 13715
rect 6310 13680 6350 13685
rect 6845 13685 6850 13715
rect 6880 13685 6885 13715
rect 6845 13680 6885 13685
rect 6900 13680 6915 14105
rect 7075 13940 7105 13945
rect 6975 13910 7075 13920
rect 8660 13940 8690 13945
rect 6975 13905 7105 13910
rect 7165 13910 7195 13915
rect 6930 13715 6960 13720
rect 6930 13680 6960 13685
rect 6975 13680 6990 13905
rect 7035 13880 7165 13890
rect 7035 13875 7195 13880
rect 8570 13910 8600 13915
rect 8690 13910 8790 13920
rect 8660 13905 8790 13910
rect 8600 13880 8730 13890
rect 8570 13875 8730 13880
rect 7035 13680 7050 13875
rect 8715 13680 8730 13875
rect 8775 13680 8790 13905
rect 9340 13715 9380 13720
rect 8805 13685 8810 13715
rect 8840 13685 8845 13715
rect 8805 13680 8845 13685
rect 9340 13685 9345 13715
rect 9375 13685 9380 13715
rect 9340 13680 9380 13685
rect 9395 13680 9410 14105
rect 9570 13940 9600 13945
rect 9470 13910 9570 13920
rect 11155 13940 11185 13945
rect 9470 13905 9600 13910
rect 9660 13910 9690 13915
rect 9425 13715 9455 13720
rect 9425 13680 9455 13685
rect 9470 13680 9485 13905
rect 9530 13880 9660 13890
rect 11065 13910 11095 13915
rect 9530 13875 9690 13880
rect 10975 13880 11005 13885
rect 9530 13680 9545 13875
rect 10885 13850 10915 13855
rect 11185 13910 11285 13920
rect 11155 13905 11285 13910
rect 11095 13880 11225 13890
rect 11065 13875 11225 13880
rect 11005 13850 11165 13860
rect 10975 13845 11165 13850
rect 10915 13820 11105 13830
rect 10885 13815 11105 13820
rect 11090 13680 11105 13815
rect 11150 13680 11165 13845
rect 11210 13680 11225 13875
rect 11270 13680 11285 13905
rect 11835 13715 11875 13720
rect 11300 13685 11305 13715
rect 11335 13685 11340 13715
rect 11300 13680 11340 13685
rect 11835 13685 11840 13715
rect 11870 13685 11875 13715
rect 11835 13680 11875 13685
rect 11890 13680 11905 14105
rect 12065 13940 12095 13945
rect 11965 13910 12065 13920
rect 13650 13940 13680 13945
rect 11965 13905 12095 13910
rect 12155 13910 12185 13915
rect 11920 13715 11950 13720
rect 11920 13680 11950 13685
rect 11965 13680 11980 13905
rect 12025 13880 12155 13890
rect 13560 13910 13590 13915
rect 12025 13875 12185 13880
rect 12245 13880 12275 13885
rect 12025 13680 12040 13875
rect 12085 13850 12245 13860
rect 13470 13880 13500 13885
rect 12085 13845 12275 13850
rect 12335 13850 12365 13855
rect 12085 13680 12100 13845
rect 12145 13820 12335 13830
rect 12145 13815 12365 13820
rect 13380 13850 13410 13855
rect 13680 13910 13780 13920
rect 13650 13905 13780 13910
rect 13590 13880 13720 13890
rect 13560 13875 13720 13880
rect 13500 13850 13660 13860
rect 13470 13845 13660 13850
rect 13410 13820 13600 13830
rect 13380 13815 13600 13820
rect 12145 13680 12160 13815
rect 13585 13680 13600 13815
rect 13645 13680 13660 13845
rect 13705 13680 13720 13875
rect 13765 13680 13780 13905
rect 14330 13715 14370 13720
rect 13795 13685 13800 13715
rect 13830 13685 13835 13715
rect 13795 13680 13835 13685
rect 14330 13685 14335 13715
rect 14365 13685 14370 13715
rect 14330 13680 14370 13685
rect 14385 13680 14400 14105
rect 14560 13940 14590 13945
rect 14460 13910 14560 13920
rect 16145 13940 16175 13945
rect 14460 13905 14590 13910
rect 14650 13910 14680 13915
rect 14415 13715 14445 13720
rect 14415 13680 14445 13685
rect 14460 13680 14475 13905
rect 14520 13880 14650 13890
rect 16055 13910 16085 13915
rect 14520 13875 14680 13880
rect 14740 13880 14770 13885
rect 14520 13680 14535 13875
rect 14580 13850 14740 13860
rect 15965 13880 15995 13885
rect 14580 13845 14770 13850
rect 14830 13850 14860 13855
rect 14580 13680 14595 13845
rect 14640 13820 14830 13830
rect 15875 13850 15905 13855
rect 14640 13815 14860 13820
rect 15785 13820 15815 13825
rect 14640 13680 14655 13815
rect 15695 13790 15725 13795
rect 16175 13910 16275 13920
rect 16145 13905 16275 13910
rect 16085 13880 16215 13890
rect 16055 13875 16215 13880
rect 15995 13850 16155 13860
rect 15965 13845 16155 13850
rect 15905 13820 16095 13830
rect 15875 13815 16095 13820
rect 15815 13790 16035 13800
rect 15785 13785 16035 13790
rect 15725 13760 15975 13770
rect 15695 13755 15975 13760
rect 15960 13680 15975 13755
rect 16020 13680 16035 13785
rect 16080 13680 16095 13815
rect 16140 13680 16155 13845
rect 16200 13680 16215 13875
rect 16260 13680 16275 13905
rect 16825 13715 16865 13720
rect 16290 13685 16295 13715
rect 16325 13685 16330 13715
rect 16290 13680 16330 13685
rect 16825 13685 16830 13715
rect 16860 13685 16865 13715
rect 16825 13680 16865 13685
rect 16880 13680 16895 14105
rect 17055 13940 17085 13945
rect 16955 13910 17055 13920
rect 18640 13940 18670 13945
rect 16955 13905 17085 13910
rect 17145 13910 17175 13915
rect 16910 13715 16940 13720
rect 16910 13680 16940 13685
rect 16955 13680 16970 13905
rect 17015 13880 17145 13890
rect 18550 13910 18580 13915
rect 17015 13875 17175 13880
rect 17235 13880 17265 13885
rect 17015 13680 17030 13875
rect 17075 13850 17235 13860
rect 18460 13880 18490 13885
rect 17075 13845 17265 13850
rect 17325 13850 17355 13855
rect 17075 13680 17090 13845
rect 17135 13820 17325 13830
rect 18370 13850 18400 13855
rect 17135 13815 17355 13820
rect 17415 13820 17445 13825
rect 17135 13680 17150 13815
rect 17195 13790 17415 13800
rect 18280 13820 18310 13825
rect 17195 13785 17445 13790
rect 17505 13790 17535 13795
rect 17195 13680 17210 13785
rect 17255 13760 17505 13770
rect 18190 13790 18220 13795
rect 17255 13755 17535 13760
rect 18100 13760 18130 13765
rect 17255 13680 17270 13755
rect 18670 13910 18770 13920
rect 18640 13905 18770 13910
rect 18580 13880 18710 13890
rect 18550 13875 18710 13880
rect 18490 13850 18650 13860
rect 18460 13845 18650 13850
rect 18400 13820 18590 13830
rect 18370 13815 18590 13820
rect 18310 13790 18530 13800
rect 18280 13785 18530 13790
rect 18220 13760 18470 13770
rect 18190 13755 18470 13760
rect 18130 13730 18410 13740
rect 18100 13725 18410 13730
rect 18395 13680 18410 13725
rect 18455 13680 18470 13755
rect 18515 13680 18530 13785
rect 18575 13680 18590 13815
rect 18635 13680 18650 13845
rect 18695 13680 18710 13875
rect 18755 13680 18770 13905
rect 19320 13715 19360 13720
rect 18785 13685 18790 13715
rect 18820 13685 18825 13715
rect 18785 13680 18825 13685
rect 19320 13685 19325 13715
rect 19355 13685 19360 13715
rect 19320 13680 19360 13685
rect 19375 13680 19390 14105
rect 19550 13940 19580 13945
rect 19450 13910 19550 13920
rect 21135 13940 21165 13945
rect 19450 13905 19580 13910
rect 19640 13910 19670 13915
rect 19405 13715 19435 13720
rect 19405 13680 19435 13685
rect 19450 13680 19465 13905
rect 19510 13880 19640 13890
rect 21045 13910 21075 13915
rect 19510 13875 19670 13880
rect 19730 13880 19760 13885
rect 19510 13680 19525 13875
rect 19570 13850 19730 13860
rect 20955 13880 20985 13885
rect 19570 13845 19760 13850
rect 19820 13850 19850 13855
rect 19570 13680 19585 13845
rect 19630 13820 19820 13830
rect 20865 13850 20895 13855
rect 19630 13815 19850 13820
rect 19910 13820 19940 13825
rect 19630 13680 19645 13815
rect 19690 13790 19910 13800
rect 20775 13820 20805 13825
rect 19690 13785 19940 13790
rect 20000 13790 20030 13795
rect 19690 13680 19705 13785
rect 19750 13760 20000 13770
rect 20685 13790 20715 13795
rect 19750 13755 20030 13760
rect 20090 13760 20120 13765
rect 19750 13680 19765 13755
rect 19810 13730 20090 13740
rect 19810 13725 20120 13730
rect 20595 13760 20625 13765
rect 21165 13910 21265 13920
rect 21135 13905 21265 13910
rect 21075 13880 21205 13890
rect 21045 13875 21205 13880
rect 20985 13850 21145 13860
rect 20955 13845 21145 13850
rect 20895 13820 21085 13830
rect 20865 13815 21085 13820
rect 20805 13790 21025 13800
rect 20775 13785 21025 13790
rect 20715 13760 20965 13770
rect 20685 13755 20965 13760
rect 20625 13730 20905 13740
rect 20595 13725 20905 13730
rect 19810 13680 19825 13725
rect 20890 13680 20905 13725
rect 20950 13680 20965 13755
rect 21010 13680 21025 13785
rect 21070 13680 21085 13815
rect 21130 13680 21145 13845
rect 21190 13680 21205 13875
rect 21250 13680 21265 13905
rect 21815 13715 21855 13720
rect 21280 13685 21285 13715
rect 21315 13685 21320 13715
rect 21280 13680 21320 13685
rect 21815 13685 21820 13715
rect 21850 13685 21855 13715
rect 21815 13680 21855 13685
rect 21870 13680 21885 14105
rect 22045 13940 22075 13945
rect 21945 13910 22045 13920
rect 23630 13940 23660 13945
rect 21945 13905 22075 13910
rect 22135 13910 22165 13915
rect 21900 13715 21930 13720
rect 21900 13680 21930 13685
rect 21945 13680 21960 13905
rect 22005 13880 22135 13890
rect 23540 13910 23570 13915
rect 22005 13875 22165 13880
rect 22225 13880 22255 13885
rect 22005 13680 22020 13875
rect 22065 13850 22225 13860
rect 23450 13880 23480 13885
rect 22065 13845 22255 13850
rect 22315 13850 22345 13855
rect 22065 13680 22080 13845
rect 22125 13820 22315 13830
rect 23360 13850 23390 13855
rect 22125 13815 22345 13820
rect 22405 13820 22435 13825
rect 22125 13680 22140 13815
rect 22185 13790 22405 13800
rect 23270 13820 23300 13825
rect 22185 13785 22435 13790
rect 22495 13790 22525 13795
rect 22185 13665 22200 13785
rect 22245 13760 22495 13770
rect 23180 13790 23210 13795
rect 22245 13755 22525 13760
rect 22585 13760 22615 13765
rect 22245 13680 22260 13755
rect 22305 13730 22585 13740
rect 23660 13910 23760 13920
rect 23630 13905 23760 13910
rect 23570 13880 23700 13890
rect 23540 13875 23700 13880
rect 23480 13850 23640 13860
rect 23450 13845 23640 13850
rect 23390 13820 23580 13830
rect 23360 13815 23580 13820
rect 23300 13790 23520 13800
rect 23270 13785 23520 13790
rect 23210 13760 23460 13770
rect 23180 13755 23460 13760
rect 22305 13725 22615 13730
rect 22305 13680 22320 13725
rect 23445 13680 23460 13755
rect 23505 13680 23520 13785
rect 23565 13680 23580 13815
rect 23625 13680 23640 13845
rect 23685 13680 23700 13875
rect 23745 13680 23760 13905
rect 24310 13715 24350 13720
rect 23775 13685 23780 13715
rect 23810 13685 23815 13715
rect 23775 13680 23815 13685
rect 24310 13685 24315 13715
rect 24345 13685 24350 13715
rect 24310 13680 24350 13685
rect 24365 13680 24380 14105
rect 24540 13940 24570 13945
rect 24440 13910 24540 13920
rect 26125 13940 26155 13945
rect 24440 13905 24570 13910
rect 24630 13910 24660 13915
rect 24395 13715 24425 13720
rect 24395 13680 24425 13685
rect 24440 13680 24455 13905
rect 24500 13880 24630 13890
rect 26035 13910 26065 13915
rect 24500 13875 24660 13880
rect 24720 13880 24750 13885
rect 24500 13680 24515 13875
rect 24560 13850 24720 13860
rect 25945 13880 25975 13885
rect 24560 13845 24750 13850
rect 24810 13850 24840 13855
rect 24560 13680 24575 13845
rect 24620 13820 24810 13830
rect 25855 13850 25885 13855
rect 24620 13815 24840 13820
rect 24900 13820 24930 13825
rect 24620 13680 24635 13815
rect 24680 13790 24900 13800
rect 26155 13910 26255 13920
rect 26125 13905 26255 13910
rect 26065 13880 26195 13890
rect 26035 13875 26195 13880
rect 25975 13850 26135 13860
rect 25945 13845 26135 13850
rect 25885 13820 26075 13830
rect 25855 13815 26075 13820
rect 24680 13785 24930 13790
rect 24990 13790 25020 13795
rect 24680 13680 24695 13785
rect 24740 13760 24990 13770
rect 24740 13755 25020 13760
rect 24740 13680 24755 13755
rect 26060 13680 26075 13815
rect 26120 13680 26135 13845
rect 26180 13680 26195 13875
rect 26240 13680 26255 13905
rect 26805 13715 26845 13720
rect 26270 13685 26275 13715
rect 26305 13685 26310 13715
rect 26270 13680 26310 13685
rect 26805 13685 26810 13715
rect 26840 13685 26845 13715
rect 26805 13680 26845 13685
rect 26860 13680 26875 14105
rect 27035 13940 27065 13945
rect 26935 13910 27035 13920
rect 28620 13940 28650 13945
rect 26935 13905 27065 13910
rect 27125 13910 27155 13915
rect 26890 13715 26920 13720
rect 26890 13680 26920 13685
rect 26935 13680 26950 13905
rect 26995 13880 27125 13890
rect 28530 13910 28560 13915
rect 26995 13875 27155 13880
rect 27215 13880 27245 13885
rect 26995 13680 27010 13875
rect 27055 13850 27215 13860
rect 28440 13880 28470 13885
rect 27055 13845 27245 13850
rect 27305 13850 27335 13855
rect 27055 13680 27070 13845
rect 27115 13820 27305 13830
rect 27115 13815 27335 13820
rect 28350 13850 28380 13855
rect 28650 13910 28750 13920
rect 28620 13905 28750 13910
rect 28560 13880 28690 13890
rect 28530 13875 28690 13880
rect 28470 13850 28630 13860
rect 28440 13845 28630 13850
rect 28380 13820 28570 13830
rect 28350 13815 28570 13820
rect 27115 13680 27130 13815
rect 28555 13680 28570 13815
rect 28615 13680 28630 13845
rect 28675 13680 28690 13875
rect 28735 13680 28750 13905
rect 29300 13715 29340 13720
rect 28765 13685 28770 13715
rect 28800 13685 28805 13715
rect 28765 13680 28805 13685
rect 29300 13685 29305 13715
rect 29335 13685 29340 13715
rect 29300 13680 29340 13685
rect 29355 13680 29370 14105
rect 29530 13940 29560 13945
rect 29430 13910 29530 13920
rect 31115 13940 31145 13945
rect 29430 13905 29560 13910
rect 29620 13910 29650 13915
rect 29385 13715 29415 13720
rect 29385 13680 29415 13685
rect 29430 13680 29445 13905
rect 29490 13880 29620 13890
rect 31025 13910 31055 13915
rect 29490 13875 29650 13880
rect 29710 13880 29740 13885
rect 29490 13680 29505 13875
rect 29550 13850 29710 13860
rect 31145 13910 31245 13920
rect 31115 13905 31245 13910
rect 31055 13880 31185 13890
rect 31025 13875 31185 13880
rect 29550 13845 29740 13850
rect 29800 13850 29830 13855
rect 29550 13680 29565 13845
rect 29610 13820 29800 13830
rect 29610 13815 29830 13820
rect 29610 13680 29625 13815
rect 31170 13680 31185 13875
rect 31230 13680 31245 13905
rect 31795 13715 31835 13720
rect 31260 13685 31265 13715
rect 31295 13685 31300 13715
rect 31260 13680 31300 13685
rect 31795 13685 31800 13715
rect 31830 13685 31835 13715
rect 31795 13680 31835 13685
rect 31850 13680 31865 14105
rect 32025 13940 32055 13945
rect 31925 13910 32025 13920
rect 33610 13940 33640 13945
rect 31925 13905 32055 13910
rect 32115 13910 32145 13915
rect 31880 13715 31910 13720
rect 31880 13680 31910 13685
rect 31925 13680 31940 13905
rect 31985 13880 32115 13890
rect 31985 13875 32145 13880
rect 33520 13910 33550 13915
rect 33640 13910 33740 13920
rect 33610 13905 33740 13910
rect 33550 13880 33680 13890
rect 33520 13875 33680 13880
rect 31985 13680 32000 13875
rect 33665 13680 33680 13875
rect 33725 13680 33740 13905
rect 34290 13715 34330 13720
rect 33755 13685 33760 13715
rect 33790 13685 33795 13715
rect 33755 13680 33795 13685
rect 34290 13685 34295 13715
rect 34325 13685 34330 13715
rect 34290 13680 34330 13685
rect 34345 13680 34360 14105
rect 34520 13940 34550 13945
rect 34420 13910 34520 13920
rect 36105 13940 36135 13945
rect 34420 13905 34550 13910
rect 34610 13910 34640 13915
rect 34375 13715 34405 13720
rect 34375 13680 34405 13685
rect 34420 13680 34435 13905
rect 34480 13880 34610 13890
rect 36135 13910 36235 13920
rect 36105 13905 36235 13910
rect 34480 13875 34640 13880
rect 34480 13680 34495 13875
rect 36220 13680 36235 13905
rect 36785 13715 36825 13720
rect 36250 13685 36255 13715
rect 36285 13685 36290 13715
rect 36250 13680 36290 13685
rect 36785 13685 36790 13715
rect 36820 13685 36825 13715
rect 36785 13680 36825 13685
rect 36840 13680 36855 14105
rect 37015 13940 37045 13945
rect 36915 13910 37015 13920
rect 36915 13905 37045 13910
rect 38600 13940 38630 13945
rect 38630 13910 38730 13920
rect 38600 13905 38730 13910
rect 36870 13715 36900 13720
rect 36870 13680 36900 13685
rect 36915 13680 36930 13905
rect 38715 13680 38730 13905
rect 39280 13715 39320 13720
rect 38745 13685 38750 13715
rect 38780 13685 38785 13715
rect 38745 13680 38785 13685
rect 39280 13685 39285 13715
rect 39315 13685 39320 13715
rect 39280 13680 39320 13685
rect 39335 13680 39350 14105
rect 39510 13940 39540 13945
rect 39410 13910 39510 13920
rect 39410 13905 39540 13910
rect 39365 13715 39395 13720
rect 39365 13680 39395 13685
rect 39410 13680 39425 13905
<< via1 >>
rect 2080 15435 2110 15465
rect 4575 15435 4605 15465
rect 7070 15435 7100 15465
rect 9565 15435 9595 15465
rect 12060 15435 12090 15465
rect 14555 15435 14585 15465
rect 17050 15435 17080 15465
rect 19545 15435 19575 15465
rect 22040 15435 22070 15465
rect 24535 15435 24565 15465
rect 27030 15435 27060 15465
rect 29525 15435 29555 15465
rect 32020 15435 32050 15465
rect 34515 15435 34545 15465
rect 37010 15435 37040 15465
rect 39505 15435 39535 15465
rect 2050 15365 2080 15395
rect 4545 15365 4575 15395
rect 7040 15365 7070 15395
rect 9535 15365 9565 15395
rect 12030 15365 12060 15395
rect 14525 15365 14555 15395
rect 17020 15365 17050 15395
rect 19515 15365 19545 15395
rect 22010 15365 22040 15395
rect 24505 15365 24535 15395
rect 27000 15365 27030 15395
rect 29495 15365 29525 15395
rect 31990 15365 32020 15395
rect 34485 15365 34515 15395
rect 36980 15365 37010 15395
rect 39475 15365 39505 15395
rect 7160 15295 7190 15325
rect 9655 15295 9685 15325
rect 12150 15295 12180 15325
rect 14645 15295 14675 15325
rect 17140 15295 17170 15325
rect 19635 15295 19665 15325
rect 22130 15295 22160 15325
rect 24625 15295 24655 15325
rect 27120 15295 27150 15325
rect 29615 15295 29645 15325
rect 32110 15295 32140 15325
rect 34605 15295 34635 15325
rect 7130 15225 7160 15255
rect 9625 15225 9655 15255
rect 12120 15225 12150 15255
rect 14615 15225 14645 15255
rect 17110 15225 17140 15255
rect 19605 15225 19635 15255
rect 22100 15225 22130 15255
rect 24595 15225 24625 15255
rect 27090 15225 27120 15255
rect 29585 15225 29615 15255
rect 32080 15225 32110 15255
rect 34575 15225 34605 15255
rect 12330 15155 12360 15185
rect 14825 15155 14855 15185
rect 17230 15155 17260 15185
rect 19725 15155 19755 15185
rect 22220 15155 22250 15185
rect 24715 15155 24745 15185
rect 27300 15155 27330 15185
rect 29795 15155 29825 15185
rect 12300 15085 12330 15115
rect 14795 15085 14825 15115
rect 17200 15085 17230 15115
rect 19695 15085 19725 15115
rect 22190 15085 22220 15115
rect 24685 15085 24715 15115
rect 27270 15085 27300 15115
rect 29765 15085 29795 15115
rect 12240 15015 12270 15045
rect 14735 15015 14765 15045
rect 17320 15015 17350 15045
rect 19815 15015 19845 15045
rect 22310 15015 22340 15045
rect 24805 15015 24835 15045
rect 27210 15015 27240 15045
rect 29705 15015 29735 15045
rect 12210 14945 12240 14975
rect 14705 14945 14735 14975
rect 17290 14945 17320 14975
rect 19785 14945 19815 14975
rect 22280 14945 22310 14975
rect 24775 14945 24805 14975
rect 27180 14945 27210 14975
rect 29675 14945 29705 14975
rect 17500 14875 17530 14905
rect 19905 14875 19935 14905
rect 22400 14875 22430 14905
rect 24985 14875 25015 14905
rect 17470 14805 17500 14835
rect 19875 14805 19905 14835
rect 22370 14805 22400 14835
rect 24955 14805 24985 14835
rect 17410 14735 17440 14765
rect 24895 14735 24925 14765
rect 17380 14665 17410 14695
rect 24865 14665 24895 14695
rect 19995 14595 20025 14625
rect 22580 14595 22610 14625
rect 19965 14525 19995 14555
rect 22550 14525 22580 14555
rect 22505 14455 22535 14485
rect 22460 14385 22490 14415
rect 20085 14315 20115 14345
rect 20050 14245 20080 14275
rect 1935 14175 1965 14205
rect 4430 14175 4460 14205
rect 6925 14175 6955 14205
rect 9420 14175 9450 14205
rect 11915 14175 11945 14205
rect 14410 14175 14440 14205
rect 16905 14175 16935 14205
rect 19400 14175 19430 14205
rect 21895 14175 21925 14205
rect 24390 14175 24420 14205
rect 26885 14175 26915 14205
rect 29380 14175 29410 14205
rect 31875 14175 31905 14205
rect 34370 14175 34400 14205
rect 36865 14175 36895 14205
rect 39360 14175 39390 14205
rect 1175 13910 1205 13940
rect 1325 13685 1355 13715
rect 1860 13685 1890 13715
rect 2085 13910 2115 13940
rect 3670 13910 3700 13940
rect 1940 13685 1970 13715
rect 3820 13685 3850 13715
rect 4355 13685 4385 13715
rect 4580 13910 4610 13940
rect 4435 13685 4465 13715
rect 6075 13880 6105 13910
rect 6165 13910 6195 13940
rect 6315 13685 6345 13715
rect 6850 13685 6880 13715
rect 7075 13910 7105 13940
rect 6930 13685 6960 13715
rect 7165 13880 7195 13910
rect 8570 13880 8600 13910
rect 8660 13910 8690 13940
rect 8810 13685 8840 13715
rect 9345 13685 9375 13715
rect 9570 13910 9600 13940
rect 9425 13685 9455 13715
rect 9660 13880 9690 13910
rect 10885 13820 10915 13850
rect 10975 13850 11005 13880
rect 11065 13880 11095 13910
rect 11155 13910 11185 13940
rect 11305 13685 11335 13715
rect 11840 13685 11870 13715
rect 12065 13910 12095 13940
rect 11920 13685 11950 13715
rect 12155 13880 12185 13910
rect 12245 13850 12275 13880
rect 12335 13820 12365 13850
rect 13380 13820 13410 13850
rect 13470 13850 13500 13880
rect 13560 13880 13590 13910
rect 13650 13910 13680 13940
rect 13800 13685 13830 13715
rect 14335 13685 14365 13715
rect 14560 13910 14590 13940
rect 14415 13685 14445 13715
rect 14650 13880 14680 13910
rect 14740 13850 14770 13880
rect 14830 13820 14860 13850
rect 15695 13760 15725 13790
rect 15785 13790 15815 13820
rect 15875 13820 15905 13850
rect 15965 13850 15995 13880
rect 16055 13880 16085 13910
rect 16145 13910 16175 13940
rect 16295 13685 16325 13715
rect 16830 13685 16860 13715
rect 17055 13910 17085 13940
rect 16910 13685 16940 13715
rect 17145 13880 17175 13910
rect 17235 13850 17265 13880
rect 17325 13820 17355 13850
rect 17415 13790 17445 13820
rect 17505 13760 17535 13790
rect 18100 13730 18130 13760
rect 18190 13760 18220 13790
rect 18280 13790 18310 13820
rect 18370 13820 18400 13850
rect 18460 13850 18490 13880
rect 18550 13880 18580 13910
rect 18640 13910 18670 13940
rect 18790 13685 18820 13715
rect 19325 13685 19355 13715
rect 19550 13910 19580 13940
rect 19405 13685 19435 13715
rect 19640 13880 19670 13910
rect 19730 13850 19760 13880
rect 19820 13820 19850 13850
rect 19910 13790 19940 13820
rect 20000 13760 20030 13790
rect 20090 13730 20120 13760
rect 20595 13730 20625 13760
rect 20685 13760 20715 13790
rect 20775 13790 20805 13820
rect 20865 13820 20895 13850
rect 20955 13850 20985 13880
rect 21045 13880 21075 13910
rect 21135 13910 21165 13940
rect 21285 13685 21315 13715
rect 21820 13685 21850 13715
rect 22045 13910 22075 13940
rect 21900 13685 21930 13715
rect 22135 13880 22165 13910
rect 22225 13850 22255 13880
rect 22315 13820 22345 13850
rect 22405 13790 22435 13820
rect 22495 13760 22525 13790
rect 22585 13730 22615 13760
rect 23180 13760 23210 13790
rect 23270 13790 23300 13820
rect 23360 13820 23390 13850
rect 23450 13850 23480 13880
rect 23540 13880 23570 13910
rect 23630 13910 23660 13940
rect 23780 13685 23810 13715
rect 24315 13685 24345 13715
rect 24540 13910 24570 13940
rect 24395 13685 24425 13715
rect 24630 13880 24660 13910
rect 24720 13850 24750 13880
rect 24810 13820 24840 13850
rect 24900 13790 24930 13820
rect 25855 13820 25885 13850
rect 25945 13850 25975 13880
rect 26035 13880 26065 13910
rect 26125 13910 26155 13940
rect 24990 13760 25020 13790
rect 26275 13685 26305 13715
rect 26810 13685 26840 13715
rect 27035 13910 27065 13940
rect 26890 13685 26920 13715
rect 27125 13880 27155 13910
rect 27215 13850 27245 13880
rect 27305 13820 27335 13850
rect 28350 13820 28380 13850
rect 28440 13850 28470 13880
rect 28530 13880 28560 13910
rect 28620 13910 28650 13940
rect 28770 13685 28800 13715
rect 29305 13685 29335 13715
rect 29530 13910 29560 13940
rect 29385 13685 29415 13715
rect 29620 13880 29650 13910
rect 29710 13850 29740 13880
rect 31025 13880 31055 13910
rect 31115 13910 31145 13940
rect 29800 13820 29830 13850
rect 31265 13685 31295 13715
rect 31800 13685 31830 13715
rect 32025 13910 32055 13940
rect 31880 13685 31910 13715
rect 32115 13880 32145 13910
rect 33520 13880 33550 13910
rect 33610 13910 33640 13940
rect 33760 13685 33790 13715
rect 34295 13685 34325 13715
rect 34520 13910 34550 13940
rect 34375 13685 34405 13715
rect 34610 13880 34640 13910
rect 36105 13910 36135 13940
rect 36255 13685 36285 13715
rect 36790 13685 36820 13715
rect 37015 13910 37045 13940
rect 38600 13910 38630 13940
rect 36870 13685 36900 13715
rect 38750 13685 38780 13715
rect 39285 13685 39315 13715
rect 39510 13910 39540 13940
rect 39365 13685 39395 13715
<< metal2 >>
rect 1175 15470 1215 15475
rect 1175 15440 1180 15470
rect 1210 15440 1215 15470
rect 3670 15470 3710 15475
rect 1175 15435 1215 15440
rect 2075 15435 2080 15465
rect 2110 15435 2115 15465
rect 1175 13945 1190 15435
rect 1205 15400 1245 15405
rect 1205 15370 1210 15400
rect 1240 15370 1245 15400
rect 1205 15365 1245 15370
rect 2045 15365 2050 15395
rect 2080 15365 2085 15395
rect 1175 13940 1205 13945
rect 1175 13905 1205 13910
rect 1220 13920 1235 15365
rect 1855 14210 1895 14215
rect 1855 14180 1860 14210
rect 1890 14180 1895 14210
rect 1855 14175 1895 14180
rect 1930 14175 1935 14205
rect 1965 14175 1970 14205
rect 1320 14140 1360 14145
rect 1320 14110 1325 14140
rect 1355 14110 1360 14140
rect 1320 14105 1360 14110
rect 1220 13905 1305 13920
rect 1290 13680 1305 13905
rect 1320 13715 1355 14105
rect 1860 13720 1895 14175
rect 1955 13720 1970 14175
rect 2055 13920 2070 15365
rect 2100 13945 2115 15435
rect 1855 13715 1895 13720
rect 1320 13685 1325 13715
rect 1355 13685 1360 13715
rect 1320 13680 1360 13685
rect 1855 13685 1860 13715
rect 1890 13685 1895 13715
rect 1855 13680 1895 13685
rect 1940 13715 1970 13720
rect 1940 13680 1970 13685
rect 1985 13905 2070 13920
rect 2085 13940 2115 13945
rect 2085 13905 2115 13910
rect 3670 15440 3675 15470
rect 3705 15440 3710 15470
rect 6165 15470 6205 15475
rect 3670 15435 3710 15440
rect 4570 15435 4575 15465
rect 4605 15435 4610 15465
rect 3670 13945 3685 15435
rect 3700 15400 3740 15405
rect 3700 15370 3705 15400
rect 3735 15370 3740 15400
rect 3700 15365 3740 15370
rect 4540 15365 4545 15395
rect 4575 15365 4580 15395
rect 3670 13940 3700 13945
rect 3670 13905 3700 13910
rect 3715 13920 3730 15365
rect 4350 14210 4390 14215
rect 4350 14180 4355 14210
rect 4385 14180 4390 14210
rect 4350 14175 4390 14180
rect 4425 14175 4430 14205
rect 4460 14175 4465 14205
rect 3815 14140 3855 14145
rect 3815 14110 3820 14140
rect 3850 14110 3855 14140
rect 3815 14105 3855 14110
rect 3715 13905 3800 13920
rect 1985 13680 2000 13905
rect 3785 13680 3800 13905
rect 3815 13715 3850 14105
rect 4355 13720 4390 14175
rect 4450 13720 4465 14175
rect 4550 13920 4565 15365
rect 4595 13945 4610 15435
rect 6165 15440 6170 15470
rect 6200 15440 6205 15470
rect 8660 15470 8700 15475
rect 6165 15435 6205 15440
rect 7065 15435 7070 15465
rect 7100 15435 7105 15465
rect 4350 13715 4390 13720
rect 3815 13685 3820 13715
rect 3850 13685 3855 13715
rect 3815 13680 3855 13685
rect 4350 13685 4355 13715
rect 4385 13685 4390 13715
rect 4350 13680 4390 13685
rect 4435 13715 4465 13720
rect 4435 13680 4465 13685
rect 4480 13905 4565 13920
rect 4580 13940 4610 13945
rect 4580 13905 4610 13910
rect 6075 15330 6115 15335
rect 6075 15300 6080 15330
rect 6110 15300 6115 15330
rect 6075 15295 6115 15300
rect 6075 13915 6090 15295
rect 6105 15260 6145 15265
rect 6105 15230 6110 15260
rect 6140 15230 6145 15260
rect 6105 15225 6145 15230
rect 6075 13910 6105 13915
rect 4480 13680 4495 13905
rect 6075 13875 6105 13880
rect 6120 13890 6135 15225
rect 6165 13945 6180 15435
rect 6195 15400 6235 15405
rect 6195 15370 6200 15400
rect 6230 15370 6235 15400
rect 6195 15365 6235 15370
rect 7035 15365 7040 15395
rect 7070 15365 7075 15395
rect 6165 13940 6195 13945
rect 6165 13905 6195 13910
rect 6210 13920 6225 15365
rect 6845 14210 6885 14215
rect 6845 14180 6850 14210
rect 6880 14180 6885 14210
rect 6845 14175 6885 14180
rect 6920 14175 6925 14205
rect 6955 14175 6960 14205
rect 6310 14140 6350 14145
rect 6310 14110 6315 14140
rect 6345 14110 6350 14140
rect 6310 14105 6350 14110
rect 6210 13905 6295 13920
rect 6120 13875 6235 13890
rect 6220 13680 6235 13875
rect 6280 13680 6295 13905
rect 6310 13715 6345 14105
rect 6850 13720 6885 14175
rect 6945 13720 6960 14175
rect 7045 13920 7060 15365
rect 7090 13945 7105 15435
rect 8660 15440 8665 15470
rect 8695 15440 8700 15470
rect 11155 15470 11195 15475
rect 8660 15435 8700 15440
rect 9560 15435 9565 15465
rect 9595 15435 9600 15465
rect 8570 15330 8610 15335
rect 7155 15295 7160 15325
rect 7190 15295 7195 15325
rect 7125 15225 7130 15255
rect 7160 15225 7165 15255
rect 6845 13715 6885 13720
rect 6310 13685 6315 13715
rect 6345 13685 6350 13715
rect 6310 13680 6350 13685
rect 6845 13685 6850 13715
rect 6880 13685 6885 13715
rect 6845 13680 6885 13685
rect 6930 13715 6960 13720
rect 6930 13680 6960 13685
rect 6975 13905 7060 13920
rect 7075 13940 7105 13945
rect 7075 13905 7105 13910
rect 6975 13680 6990 13905
rect 7135 13890 7150 15225
rect 7180 13915 7195 15295
rect 7035 13875 7150 13890
rect 7165 13910 7195 13915
rect 7165 13875 7195 13880
rect 8570 15300 8575 15330
rect 8605 15300 8610 15330
rect 8570 15295 8610 15300
rect 8570 13915 8585 15295
rect 8600 15260 8640 15265
rect 8600 15230 8605 15260
rect 8635 15230 8640 15260
rect 8600 15225 8640 15230
rect 8570 13910 8600 13915
rect 8570 13875 8600 13880
rect 8615 13890 8630 15225
rect 8660 13945 8675 15435
rect 8690 15400 8730 15405
rect 8690 15370 8695 15400
rect 8725 15370 8730 15400
rect 8690 15365 8730 15370
rect 9530 15365 9535 15395
rect 9565 15365 9570 15395
rect 8660 13940 8690 13945
rect 8660 13905 8690 13910
rect 8705 13920 8720 15365
rect 9340 14210 9380 14215
rect 9340 14180 9345 14210
rect 9375 14180 9380 14210
rect 9340 14175 9380 14180
rect 9415 14175 9420 14205
rect 9450 14175 9455 14205
rect 8805 14140 8845 14145
rect 8805 14110 8810 14140
rect 8840 14110 8845 14140
rect 8805 14105 8845 14110
rect 8705 13905 8790 13920
rect 8615 13875 8730 13890
rect 7035 13680 7050 13875
rect 8715 13680 8730 13875
rect 8775 13680 8790 13905
rect 8805 13715 8840 14105
rect 9345 13720 9380 14175
rect 9440 13720 9455 14175
rect 9540 13920 9555 15365
rect 9585 13945 9600 15435
rect 11155 15440 11160 15470
rect 11190 15440 11195 15470
rect 13650 15470 13690 15475
rect 11155 15435 11195 15440
rect 12055 15435 12060 15465
rect 12090 15435 12095 15465
rect 11065 15330 11105 15335
rect 9650 15295 9655 15325
rect 9685 15295 9690 15325
rect 9620 15225 9625 15255
rect 9655 15225 9660 15255
rect 9340 13715 9380 13720
rect 8805 13685 8810 13715
rect 8840 13685 8845 13715
rect 8805 13680 8845 13685
rect 9340 13685 9345 13715
rect 9375 13685 9380 13715
rect 9340 13680 9380 13685
rect 9425 13715 9455 13720
rect 9425 13680 9455 13685
rect 9470 13905 9555 13920
rect 9570 13940 9600 13945
rect 9570 13905 9600 13910
rect 9470 13680 9485 13905
rect 9630 13890 9645 15225
rect 9675 13915 9690 15295
rect 11065 15300 11070 15330
rect 11100 15300 11105 15330
rect 11065 15295 11105 15300
rect 9530 13875 9645 13890
rect 9660 13910 9690 13915
rect 9660 13875 9690 13880
rect 10885 15190 10925 15195
rect 10885 15160 10890 15190
rect 10920 15160 10925 15190
rect 10885 15155 10925 15160
rect 9530 13680 9545 13875
rect 10885 13855 10900 15155
rect 10915 15120 10955 15125
rect 10915 15090 10920 15120
rect 10950 15090 10955 15120
rect 10915 15085 10955 15090
rect 10885 13850 10915 13855
rect 10885 13815 10915 13820
rect 10930 13830 10945 15085
rect 10975 15050 11015 15055
rect 10975 15020 10980 15050
rect 11010 15020 11015 15050
rect 10975 15015 11015 15020
rect 10975 13885 10990 15015
rect 11005 14980 11045 14985
rect 11005 14950 11010 14980
rect 11040 14950 11045 14980
rect 11005 14945 11045 14950
rect 10975 13880 11005 13885
rect 10975 13845 11005 13850
rect 11020 13860 11035 14945
rect 11065 13915 11080 15295
rect 11095 15260 11135 15265
rect 11095 15230 11100 15260
rect 11130 15230 11135 15260
rect 11095 15225 11135 15230
rect 11065 13910 11095 13915
rect 11065 13875 11095 13880
rect 11110 13890 11125 15225
rect 11155 13945 11170 15435
rect 11185 15400 11225 15405
rect 11185 15370 11190 15400
rect 11220 15370 11225 15400
rect 11185 15365 11225 15370
rect 12025 15365 12030 15395
rect 12060 15365 12065 15395
rect 11155 13940 11185 13945
rect 11155 13905 11185 13910
rect 11200 13920 11215 15365
rect 11835 14210 11875 14215
rect 11835 14180 11840 14210
rect 11870 14180 11875 14210
rect 11835 14175 11875 14180
rect 11910 14175 11915 14205
rect 11945 14175 11950 14205
rect 11300 14140 11340 14145
rect 11300 14110 11305 14140
rect 11335 14110 11340 14140
rect 11300 14105 11340 14110
rect 11200 13905 11285 13920
rect 11110 13875 11225 13890
rect 11020 13845 11165 13860
rect 10930 13815 11105 13830
rect 11090 13680 11105 13815
rect 11150 13680 11165 13845
rect 11210 13680 11225 13875
rect 11270 13680 11285 13905
rect 11300 13715 11335 14105
rect 11840 13720 11875 14175
rect 11935 13720 11950 14175
rect 12035 13920 12050 15365
rect 12080 13945 12095 15435
rect 13650 15440 13655 15470
rect 13685 15440 13690 15470
rect 16145 15470 16185 15475
rect 13650 15435 13690 15440
rect 14550 15435 14555 15465
rect 14585 15435 14590 15465
rect 13560 15330 13600 15335
rect 12145 15295 12150 15325
rect 12180 15295 12185 15325
rect 12115 15225 12120 15255
rect 12150 15225 12155 15255
rect 11835 13715 11875 13720
rect 11300 13685 11305 13715
rect 11335 13685 11340 13715
rect 11300 13680 11340 13685
rect 11835 13685 11840 13715
rect 11870 13685 11875 13715
rect 11835 13680 11875 13685
rect 11920 13715 11950 13720
rect 11920 13680 11950 13685
rect 11965 13905 12050 13920
rect 12065 13940 12095 13945
rect 12065 13905 12095 13910
rect 11965 13680 11980 13905
rect 12125 13890 12140 15225
rect 12170 13915 12185 15295
rect 13560 15300 13565 15330
rect 13595 15300 13600 15330
rect 13560 15295 13600 15300
rect 13380 15190 13420 15195
rect 12325 15155 12330 15185
rect 12360 15155 12365 15185
rect 12295 15085 12300 15115
rect 12330 15085 12335 15115
rect 12235 15015 12240 15045
rect 12270 15015 12275 15045
rect 12205 14945 12210 14975
rect 12240 14945 12245 14975
rect 12025 13875 12140 13890
rect 12155 13910 12185 13915
rect 12155 13875 12185 13880
rect 12025 13680 12040 13875
rect 12215 13860 12230 14945
rect 12260 13885 12275 15015
rect 12085 13845 12230 13860
rect 12245 13880 12275 13885
rect 12245 13845 12275 13850
rect 12085 13680 12100 13845
rect 12305 13830 12320 15085
rect 12350 13855 12365 15155
rect 12145 13815 12320 13830
rect 12335 13850 12365 13855
rect 12335 13815 12365 13820
rect 13380 15160 13385 15190
rect 13415 15160 13420 15190
rect 13380 15155 13420 15160
rect 13380 13855 13395 15155
rect 13410 15120 13450 15125
rect 13410 15090 13415 15120
rect 13445 15090 13450 15120
rect 13410 15085 13450 15090
rect 13380 13850 13410 13855
rect 13380 13815 13410 13820
rect 13425 13830 13440 15085
rect 13470 15050 13510 15055
rect 13470 15020 13475 15050
rect 13505 15020 13510 15050
rect 13470 15015 13510 15020
rect 13470 13885 13485 15015
rect 13500 14980 13540 14985
rect 13500 14950 13505 14980
rect 13535 14950 13540 14980
rect 13500 14945 13540 14950
rect 13470 13880 13500 13885
rect 13470 13845 13500 13850
rect 13515 13860 13530 14945
rect 13560 13915 13575 15295
rect 13590 15260 13630 15265
rect 13590 15230 13595 15260
rect 13625 15230 13630 15260
rect 13590 15225 13630 15230
rect 13560 13910 13590 13915
rect 13560 13875 13590 13880
rect 13605 13890 13620 15225
rect 13650 13945 13665 15435
rect 13680 15400 13720 15405
rect 13680 15370 13685 15400
rect 13715 15370 13720 15400
rect 13680 15365 13720 15370
rect 14520 15365 14525 15395
rect 14555 15365 14560 15395
rect 13650 13940 13680 13945
rect 13650 13905 13680 13910
rect 13695 13920 13710 15365
rect 14330 14210 14370 14215
rect 14330 14180 14335 14210
rect 14365 14180 14370 14210
rect 14330 14175 14370 14180
rect 14405 14175 14410 14205
rect 14440 14175 14445 14205
rect 13795 14140 13835 14145
rect 13795 14110 13800 14140
rect 13830 14110 13835 14140
rect 13795 14105 13835 14110
rect 13695 13905 13780 13920
rect 13605 13875 13720 13890
rect 13515 13845 13660 13860
rect 13425 13815 13600 13830
rect 12145 13680 12160 13815
rect 13585 13680 13600 13815
rect 13645 13680 13660 13845
rect 13705 13680 13720 13875
rect 13765 13680 13780 13905
rect 13795 13715 13830 14105
rect 14335 13720 14370 14175
rect 14430 13720 14445 14175
rect 14530 13920 14545 15365
rect 14575 13945 14590 15435
rect 16145 15440 16150 15470
rect 16180 15440 16185 15470
rect 18640 15470 18680 15475
rect 16145 15435 16185 15440
rect 17045 15435 17050 15465
rect 17080 15435 17085 15465
rect 16055 15330 16095 15335
rect 14640 15295 14645 15325
rect 14675 15295 14680 15325
rect 14610 15225 14615 15255
rect 14645 15225 14650 15255
rect 14330 13715 14370 13720
rect 13795 13685 13800 13715
rect 13830 13685 13835 13715
rect 13795 13680 13835 13685
rect 14330 13685 14335 13715
rect 14365 13685 14370 13715
rect 14330 13680 14370 13685
rect 14415 13715 14445 13720
rect 14415 13680 14445 13685
rect 14460 13905 14545 13920
rect 14560 13940 14590 13945
rect 14560 13905 14590 13910
rect 14460 13680 14475 13905
rect 14620 13890 14635 15225
rect 14665 13915 14680 15295
rect 16055 15300 16060 15330
rect 16090 15300 16095 15330
rect 16055 15295 16095 15300
rect 15965 15190 16005 15195
rect 14820 15155 14825 15185
rect 14855 15155 14860 15185
rect 14790 15085 14795 15115
rect 14825 15085 14830 15115
rect 14730 15015 14735 15045
rect 14765 15015 14770 15045
rect 14700 14945 14705 14975
rect 14735 14945 14740 14975
rect 14520 13875 14635 13890
rect 14650 13910 14680 13915
rect 14650 13875 14680 13880
rect 14520 13680 14535 13875
rect 14710 13860 14725 14945
rect 14755 13885 14770 15015
rect 14580 13845 14725 13860
rect 14740 13880 14770 13885
rect 14740 13845 14770 13850
rect 14580 13680 14595 13845
rect 14800 13830 14815 15085
rect 14845 13855 14860 15155
rect 15965 15160 15970 15190
rect 16000 15160 16005 15190
rect 15965 15155 16005 15160
rect 15875 15050 15915 15055
rect 15875 15020 15880 15050
rect 15910 15020 15915 15050
rect 15875 15015 15915 15020
rect 14640 13815 14815 13830
rect 14830 13850 14860 13855
rect 14830 13815 14860 13820
rect 15695 14910 15735 14915
rect 15695 14880 15700 14910
rect 15730 14880 15735 14910
rect 15695 14875 15735 14880
rect 14640 13680 14655 13815
rect 15695 13795 15710 14875
rect 15725 14840 15765 14845
rect 15725 14810 15730 14840
rect 15760 14810 15765 14840
rect 15725 14805 15765 14810
rect 15695 13790 15725 13795
rect 15695 13755 15725 13760
rect 15740 13770 15755 14805
rect 15785 14770 15825 14775
rect 15785 14740 15790 14770
rect 15820 14740 15825 14770
rect 15785 14735 15825 14740
rect 15785 13825 15800 14735
rect 15815 14700 15855 14705
rect 15815 14670 15820 14700
rect 15850 14670 15855 14700
rect 15815 14665 15855 14670
rect 15785 13820 15815 13825
rect 15785 13785 15815 13790
rect 15830 13800 15845 14665
rect 15875 13855 15890 15015
rect 15905 14980 15945 14985
rect 15905 14950 15910 14980
rect 15940 14950 15945 14980
rect 15905 14945 15945 14950
rect 15875 13850 15905 13855
rect 15875 13815 15905 13820
rect 15920 13830 15935 14945
rect 15965 13885 15980 15155
rect 15995 15120 16035 15125
rect 15995 15090 16000 15120
rect 16030 15090 16035 15120
rect 15995 15085 16035 15090
rect 15965 13880 15995 13885
rect 15965 13845 15995 13850
rect 16010 13860 16025 15085
rect 16055 13915 16070 15295
rect 16085 15260 16125 15265
rect 16085 15230 16090 15260
rect 16120 15230 16125 15260
rect 16085 15225 16125 15230
rect 16055 13910 16085 13915
rect 16055 13875 16085 13880
rect 16100 13890 16115 15225
rect 16145 13945 16160 15435
rect 16175 15400 16215 15405
rect 16175 15370 16180 15400
rect 16210 15370 16215 15400
rect 16175 15365 16215 15370
rect 17015 15365 17020 15395
rect 17050 15365 17055 15395
rect 16145 13940 16175 13945
rect 16145 13905 16175 13910
rect 16190 13920 16205 15365
rect 16825 14210 16865 14215
rect 16825 14180 16830 14210
rect 16860 14180 16865 14210
rect 16825 14175 16865 14180
rect 16900 14175 16905 14205
rect 16935 14175 16940 14205
rect 16290 14140 16330 14145
rect 16290 14110 16295 14140
rect 16325 14110 16330 14140
rect 16290 14105 16330 14110
rect 16190 13905 16275 13920
rect 16100 13875 16215 13890
rect 16010 13845 16155 13860
rect 15920 13815 16095 13830
rect 15830 13785 16035 13800
rect 15740 13755 15975 13770
rect 15960 13680 15975 13755
rect 16020 13680 16035 13785
rect 16080 13680 16095 13815
rect 16140 13680 16155 13845
rect 16200 13680 16215 13875
rect 16260 13680 16275 13905
rect 16290 13715 16325 14105
rect 16830 13720 16865 14175
rect 16925 13720 16940 14175
rect 17025 13920 17040 15365
rect 17070 13945 17085 15435
rect 18640 15440 18645 15470
rect 18675 15440 18680 15470
rect 21135 15470 21175 15475
rect 18640 15435 18680 15440
rect 19540 15435 19545 15465
rect 19575 15435 19580 15465
rect 18550 15330 18590 15335
rect 17135 15295 17140 15325
rect 17170 15295 17175 15325
rect 17105 15225 17110 15255
rect 17140 15225 17145 15255
rect 16825 13715 16865 13720
rect 16290 13685 16295 13715
rect 16325 13685 16330 13715
rect 16290 13680 16330 13685
rect 16825 13685 16830 13715
rect 16860 13685 16865 13715
rect 16825 13680 16865 13685
rect 16910 13715 16940 13720
rect 16910 13680 16940 13685
rect 16955 13905 17040 13920
rect 17055 13940 17085 13945
rect 17055 13905 17085 13910
rect 16955 13680 16970 13905
rect 17115 13890 17130 15225
rect 17160 13915 17175 15295
rect 18550 15300 18555 15330
rect 18585 15300 18590 15330
rect 18550 15295 18590 15300
rect 18460 15190 18500 15195
rect 17225 15155 17230 15185
rect 17260 15155 17265 15185
rect 17195 15085 17200 15115
rect 17230 15085 17235 15115
rect 17015 13875 17130 13890
rect 17145 13910 17175 13915
rect 17145 13875 17175 13880
rect 17015 13680 17030 13875
rect 17205 13860 17220 15085
rect 17250 13885 17265 15155
rect 18460 15160 18465 15190
rect 18495 15160 18500 15190
rect 18460 15155 18500 15160
rect 18370 15050 18410 15055
rect 17315 15015 17320 15045
rect 17350 15015 17355 15045
rect 17285 14945 17290 14975
rect 17320 14945 17325 14975
rect 17075 13845 17220 13860
rect 17235 13880 17265 13885
rect 17235 13845 17265 13850
rect 17075 13680 17090 13845
rect 17295 13830 17310 14945
rect 17340 13855 17355 15015
rect 18370 15020 18375 15050
rect 18405 15020 18410 15050
rect 18370 15015 18410 15020
rect 18280 14910 18320 14915
rect 17495 14875 17500 14905
rect 17530 14875 17535 14905
rect 17465 14805 17470 14835
rect 17500 14805 17505 14835
rect 17405 14735 17410 14765
rect 17440 14735 17445 14765
rect 17375 14665 17380 14695
rect 17410 14665 17415 14695
rect 17135 13815 17310 13830
rect 17325 13850 17355 13855
rect 17325 13815 17355 13820
rect 17135 13680 17150 13815
rect 17385 13800 17400 14665
rect 17430 13825 17445 14735
rect 17195 13785 17400 13800
rect 17415 13820 17445 13825
rect 17415 13785 17445 13790
rect 17195 13680 17210 13785
rect 17475 13770 17490 14805
rect 17520 13795 17535 14875
rect 18280 14880 18285 14910
rect 18315 14880 18320 14910
rect 18280 14875 18320 14880
rect 18190 14630 18230 14635
rect 18190 14600 18195 14630
rect 18225 14600 18230 14630
rect 18190 14595 18230 14600
rect 17255 13755 17490 13770
rect 17505 13790 17535 13795
rect 17505 13755 17535 13760
rect 18100 14350 18140 14355
rect 18100 14320 18105 14350
rect 18135 14320 18140 14350
rect 18100 14315 18140 14320
rect 18100 13765 18115 14315
rect 18130 14280 18170 14285
rect 18130 14250 18135 14280
rect 18165 14250 18170 14280
rect 18130 14245 18170 14250
rect 18100 13760 18130 13765
rect 17255 13680 17270 13755
rect 18100 13725 18130 13730
rect 18145 13740 18160 14245
rect 18190 13795 18205 14595
rect 18220 14560 18260 14565
rect 18220 14530 18225 14560
rect 18255 14530 18260 14560
rect 18220 14525 18260 14530
rect 18190 13790 18220 13795
rect 18190 13755 18220 13760
rect 18235 13770 18250 14525
rect 18280 13825 18295 14875
rect 18310 14840 18350 14845
rect 18310 14810 18315 14840
rect 18345 14810 18350 14840
rect 18310 14805 18350 14810
rect 18280 13820 18310 13825
rect 18280 13785 18310 13790
rect 18325 13800 18340 14805
rect 18370 13855 18385 15015
rect 18400 14980 18440 14985
rect 18400 14950 18405 14980
rect 18435 14950 18440 14980
rect 18400 14945 18440 14950
rect 18370 13850 18400 13855
rect 18370 13815 18400 13820
rect 18415 13830 18430 14945
rect 18460 13885 18475 15155
rect 18490 15120 18530 15125
rect 18490 15090 18495 15120
rect 18525 15090 18530 15120
rect 18490 15085 18530 15090
rect 18460 13880 18490 13885
rect 18460 13845 18490 13850
rect 18505 13860 18520 15085
rect 18550 13915 18565 15295
rect 18580 15260 18620 15265
rect 18580 15230 18585 15260
rect 18615 15230 18620 15260
rect 18580 15225 18620 15230
rect 18550 13910 18580 13915
rect 18550 13875 18580 13880
rect 18595 13890 18610 15225
rect 18640 13945 18655 15435
rect 18670 15400 18710 15405
rect 18670 15370 18675 15400
rect 18705 15370 18710 15400
rect 18670 15365 18710 15370
rect 19510 15365 19515 15395
rect 19545 15365 19550 15395
rect 18640 13940 18670 13945
rect 18640 13905 18670 13910
rect 18685 13920 18700 15365
rect 19320 14210 19360 14215
rect 19320 14180 19325 14210
rect 19355 14180 19360 14210
rect 19320 14175 19360 14180
rect 19395 14175 19400 14205
rect 19430 14175 19435 14205
rect 18785 14140 18825 14145
rect 18785 14110 18790 14140
rect 18820 14110 18825 14140
rect 18785 14105 18825 14110
rect 18685 13905 18770 13920
rect 18595 13875 18710 13890
rect 18505 13845 18650 13860
rect 18415 13815 18590 13830
rect 18325 13785 18530 13800
rect 18235 13755 18470 13770
rect 18145 13725 18410 13740
rect 18395 13680 18410 13725
rect 18455 13680 18470 13755
rect 18515 13680 18530 13785
rect 18575 13680 18590 13815
rect 18635 13680 18650 13845
rect 18695 13680 18710 13875
rect 18755 13680 18770 13905
rect 18785 13715 18820 14105
rect 19325 13720 19360 14175
rect 19420 13720 19435 14175
rect 19520 13920 19535 15365
rect 19565 13945 19580 15435
rect 21135 15440 21140 15470
rect 21170 15440 21175 15470
rect 23630 15470 23670 15475
rect 21135 15435 21175 15440
rect 22035 15435 22040 15465
rect 22070 15435 22075 15465
rect 21045 15330 21085 15335
rect 19630 15295 19635 15325
rect 19665 15295 19670 15325
rect 19600 15225 19605 15255
rect 19635 15225 19640 15255
rect 19320 13715 19360 13720
rect 18785 13685 18790 13715
rect 18820 13685 18825 13715
rect 18785 13680 18825 13685
rect 19320 13685 19325 13715
rect 19355 13685 19360 13715
rect 19320 13680 19360 13685
rect 19405 13715 19435 13720
rect 19405 13680 19435 13685
rect 19450 13905 19535 13920
rect 19550 13940 19580 13945
rect 19550 13905 19580 13910
rect 19450 13680 19465 13905
rect 19610 13890 19625 15225
rect 19655 13915 19670 15295
rect 21045 15300 21050 15330
rect 21080 15300 21085 15330
rect 21045 15295 21085 15300
rect 20955 15190 20995 15195
rect 19720 15155 19725 15185
rect 19755 15155 19760 15185
rect 19690 15085 19695 15115
rect 19725 15085 19730 15115
rect 19510 13875 19625 13890
rect 19640 13910 19670 13915
rect 19640 13875 19670 13880
rect 19510 13680 19525 13875
rect 19700 13860 19715 15085
rect 19745 13885 19760 15155
rect 20955 15160 20960 15190
rect 20990 15160 20995 15190
rect 20955 15155 20995 15160
rect 20865 15050 20905 15055
rect 19810 15015 19815 15045
rect 19845 15015 19850 15045
rect 19780 14945 19785 14975
rect 19815 14945 19820 14975
rect 19570 13845 19715 13860
rect 19730 13880 19760 13885
rect 19730 13845 19760 13850
rect 19570 13680 19585 13845
rect 19790 13830 19805 14945
rect 19835 13855 19850 15015
rect 20865 15020 20870 15050
rect 20900 15020 20905 15050
rect 20865 15015 20905 15020
rect 20775 14910 20815 14915
rect 19900 14875 19905 14905
rect 19935 14875 19940 14905
rect 19870 14805 19875 14835
rect 19905 14805 19910 14835
rect 19630 13815 19805 13830
rect 19820 13850 19850 13855
rect 19820 13815 19850 13820
rect 19630 13680 19645 13815
rect 19880 13800 19895 14805
rect 19925 13825 19940 14875
rect 20775 14880 20780 14910
rect 20810 14880 20815 14910
rect 20775 14875 20815 14880
rect 20595 14630 20635 14635
rect 19990 14595 19995 14625
rect 20025 14595 20030 14625
rect 19960 14525 19965 14555
rect 19995 14525 20000 14555
rect 19690 13785 19895 13800
rect 19910 13820 19940 13825
rect 19910 13785 19940 13790
rect 19690 13680 19705 13785
rect 19970 13770 19985 14525
rect 20015 13795 20030 14595
rect 20595 14600 20600 14630
rect 20630 14600 20635 14630
rect 20595 14595 20635 14600
rect 20080 14315 20085 14345
rect 20115 14315 20120 14345
rect 20045 14245 20050 14275
rect 20080 14245 20085 14275
rect 19750 13755 19985 13770
rect 20000 13790 20030 13795
rect 20000 13755 20030 13760
rect 19750 13680 19765 13755
rect 20060 13740 20075 14245
rect 20105 13765 20120 14315
rect 19810 13725 20075 13740
rect 20090 13760 20120 13765
rect 20090 13725 20120 13730
rect 20595 13765 20610 14595
rect 20625 14560 20665 14565
rect 20625 14530 20630 14560
rect 20660 14530 20665 14560
rect 20625 14525 20665 14530
rect 20595 13760 20625 13765
rect 20595 13725 20625 13730
rect 20640 13740 20655 14525
rect 20670 14490 20710 14495
rect 20670 14460 20675 14490
rect 20705 14460 20710 14490
rect 20670 14455 20710 14460
rect 20685 13795 20700 14455
rect 20715 14420 20755 14425
rect 20715 14390 20720 14420
rect 20750 14390 20755 14420
rect 20715 14385 20755 14390
rect 20685 13790 20715 13795
rect 20685 13755 20715 13760
rect 20730 13770 20745 14385
rect 20775 13825 20790 14875
rect 20805 14840 20845 14845
rect 20805 14810 20810 14840
rect 20840 14810 20845 14840
rect 20805 14805 20845 14810
rect 20775 13820 20805 13825
rect 20775 13785 20805 13790
rect 20820 13800 20835 14805
rect 20865 13855 20880 15015
rect 20895 14980 20935 14985
rect 20895 14950 20900 14980
rect 20930 14950 20935 14980
rect 20895 14945 20935 14950
rect 20865 13850 20895 13855
rect 20865 13815 20895 13820
rect 20910 13830 20925 14945
rect 20955 13885 20970 15155
rect 20985 15120 21025 15125
rect 20985 15090 20990 15120
rect 21020 15090 21025 15120
rect 20985 15085 21025 15090
rect 20955 13880 20985 13885
rect 20955 13845 20985 13850
rect 21000 13860 21015 15085
rect 21045 13915 21060 15295
rect 21075 15260 21115 15265
rect 21075 15230 21080 15260
rect 21110 15230 21115 15260
rect 21075 15225 21115 15230
rect 21045 13910 21075 13915
rect 21045 13875 21075 13880
rect 21090 13890 21105 15225
rect 21135 13945 21150 15435
rect 21165 15400 21205 15405
rect 21165 15370 21170 15400
rect 21200 15370 21205 15400
rect 21165 15365 21205 15370
rect 22005 15365 22010 15395
rect 22040 15365 22045 15395
rect 21135 13940 21165 13945
rect 21135 13905 21165 13910
rect 21180 13920 21195 15365
rect 21815 14210 21855 14215
rect 21815 14180 21820 14210
rect 21850 14180 21855 14210
rect 21815 14175 21855 14180
rect 21890 14175 21895 14205
rect 21925 14175 21930 14205
rect 21280 14140 21320 14145
rect 21280 14110 21285 14140
rect 21315 14110 21320 14140
rect 21280 14105 21320 14110
rect 21180 13905 21265 13920
rect 21090 13875 21205 13890
rect 21000 13845 21145 13860
rect 20910 13815 21085 13830
rect 20820 13785 21025 13800
rect 20730 13755 20965 13770
rect 20640 13725 20905 13740
rect 19810 13680 19825 13725
rect 20890 13680 20905 13725
rect 20950 13680 20965 13755
rect 21010 13680 21025 13785
rect 21070 13680 21085 13815
rect 21130 13680 21145 13845
rect 21190 13680 21205 13875
rect 21250 13680 21265 13905
rect 21280 13715 21315 14105
rect 21820 13720 21855 14175
rect 21915 13720 21930 14175
rect 22015 13920 22030 15365
rect 22060 13945 22075 15435
rect 23630 15440 23635 15470
rect 23665 15440 23670 15470
rect 26125 15470 26165 15475
rect 23630 15435 23670 15440
rect 24530 15435 24535 15465
rect 24565 15435 24570 15465
rect 23540 15330 23580 15335
rect 22125 15295 22130 15325
rect 22160 15295 22165 15325
rect 22095 15225 22100 15255
rect 22130 15225 22135 15255
rect 21815 13715 21855 13720
rect 21280 13685 21285 13715
rect 21315 13685 21320 13715
rect 21280 13680 21320 13685
rect 21815 13685 21820 13715
rect 21850 13685 21855 13715
rect 21815 13680 21855 13685
rect 21900 13715 21930 13720
rect 21900 13680 21930 13685
rect 21945 13905 22030 13920
rect 22045 13940 22075 13945
rect 22045 13905 22075 13910
rect 21945 13680 21960 13905
rect 22105 13890 22120 15225
rect 22150 13915 22165 15295
rect 23540 15300 23545 15330
rect 23575 15300 23580 15330
rect 23540 15295 23580 15300
rect 23450 15190 23490 15195
rect 22215 15155 22220 15185
rect 22250 15155 22255 15185
rect 22185 15085 22190 15115
rect 22220 15085 22225 15115
rect 22005 13875 22120 13890
rect 22135 13910 22165 13915
rect 22135 13875 22165 13880
rect 22005 13680 22020 13875
rect 22195 13860 22210 15085
rect 22240 13885 22255 15155
rect 23450 15160 23455 15190
rect 23485 15160 23490 15190
rect 23450 15155 23490 15160
rect 23360 15050 23400 15055
rect 22305 15015 22310 15045
rect 22340 15015 22345 15045
rect 22275 14945 22280 14975
rect 22310 14945 22315 14975
rect 22065 13845 22210 13860
rect 22225 13880 22255 13885
rect 22225 13845 22255 13850
rect 22065 13680 22080 13845
rect 22285 13830 22300 14945
rect 22330 13855 22345 15015
rect 23360 15020 23365 15050
rect 23395 15020 23400 15050
rect 23360 15015 23400 15020
rect 23180 14910 23220 14915
rect 22395 14875 22400 14905
rect 22430 14875 22435 14905
rect 22365 14805 22370 14835
rect 22400 14805 22405 14835
rect 22125 13815 22300 13830
rect 22315 13850 22345 13855
rect 22315 13815 22345 13820
rect 22125 13680 22140 13815
rect 22375 13800 22390 14805
rect 22420 13825 22435 14875
rect 23180 14880 23185 14910
rect 23215 14880 23220 14910
rect 23180 14875 23220 14880
rect 22575 14595 22580 14625
rect 22610 14595 22615 14625
rect 22545 14525 22550 14555
rect 22580 14525 22585 14555
rect 22500 14455 22505 14485
rect 22535 14455 22540 14485
rect 22455 14385 22460 14415
rect 22490 14385 22495 14415
rect 22185 13785 22390 13800
rect 22405 13820 22435 13825
rect 22405 13785 22435 13790
rect 22185 13665 22200 13785
rect 22465 13770 22480 14385
rect 22510 13795 22525 14455
rect 22245 13755 22480 13770
rect 22495 13790 22525 13795
rect 22495 13755 22525 13760
rect 22245 13680 22260 13755
rect 22555 13740 22570 14525
rect 22600 13765 22615 14595
rect 22305 13725 22570 13740
rect 22585 13760 22615 13765
rect 23180 13795 23195 14875
rect 23210 14840 23250 14845
rect 23210 14810 23215 14840
rect 23245 14810 23250 14840
rect 23210 14805 23250 14810
rect 23180 13790 23210 13795
rect 23180 13755 23210 13760
rect 23225 13770 23240 14805
rect 23270 14770 23310 14775
rect 23270 14740 23275 14770
rect 23305 14740 23310 14770
rect 23270 14735 23310 14740
rect 23270 13825 23285 14735
rect 23300 14700 23340 14705
rect 23300 14670 23305 14700
rect 23335 14670 23340 14700
rect 23300 14665 23340 14670
rect 23270 13820 23300 13825
rect 23270 13785 23300 13790
rect 23315 13800 23330 14665
rect 23360 13855 23375 15015
rect 23390 14980 23430 14985
rect 23390 14950 23395 14980
rect 23425 14950 23430 14980
rect 23390 14945 23430 14950
rect 23360 13850 23390 13855
rect 23360 13815 23390 13820
rect 23405 13830 23420 14945
rect 23450 13885 23465 15155
rect 23480 15120 23520 15125
rect 23480 15090 23485 15120
rect 23515 15090 23520 15120
rect 23480 15085 23520 15090
rect 23450 13880 23480 13885
rect 23450 13845 23480 13850
rect 23495 13860 23510 15085
rect 23540 13915 23555 15295
rect 23570 15260 23610 15265
rect 23570 15230 23575 15260
rect 23605 15230 23610 15260
rect 23570 15225 23610 15230
rect 23540 13910 23570 13915
rect 23540 13875 23570 13880
rect 23585 13890 23600 15225
rect 23630 13945 23645 15435
rect 23660 15400 23700 15405
rect 23660 15370 23665 15400
rect 23695 15370 23700 15400
rect 23660 15365 23700 15370
rect 24500 15365 24505 15395
rect 24535 15365 24540 15395
rect 23630 13940 23660 13945
rect 23630 13905 23660 13910
rect 23675 13920 23690 15365
rect 24310 14210 24350 14215
rect 24310 14180 24315 14210
rect 24345 14180 24350 14210
rect 24310 14175 24350 14180
rect 24385 14175 24390 14205
rect 24420 14175 24425 14205
rect 23775 14140 23815 14145
rect 23775 14110 23780 14140
rect 23810 14110 23815 14140
rect 23775 14105 23815 14110
rect 23675 13905 23760 13920
rect 23585 13875 23700 13890
rect 23495 13845 23640 13860
rect 23405 13815 23580 13830
rect 23315 13785 23520 13800
rect 23225 13755 23460 13770
rect 22585 13725 22615 13730
rect 22305 13680 22320 13725
rect 23445 13680 23460 13755
rect 23505 13680 23520 13785
rect 23565 13680 23580 13815
rect 23625 13680 23640 13845
rect 23685 13680 23700 13875
rect 23745 13680 23760 13905
rect 23775 13715 23810 14105
rect 24315 13720 24350 14175
rect 24410 13720 24425 14175
rect 24510 13920 24525 15365
rect 24555 13945 24570 15435
rect 26125 15440 26130 15470
rect 26160 15440 26165 15470
rect 28620 15470 28660 15475
rect 26125 15435 26165 15440
rect 27025 15435 27030 15465
rect 27060 15435 27065 15465
rect 26035 15330 26075 15335
rect 24620 15295 24625 15325
rect 24655 15295 24660 15325
rect 24590 15225 24595 15255
rect 24625 15225 24630 15255
rect 24310 13715 24350 13720
rect 23775 13685 23780 13715
rect 23810 13685 23815 13715
rect 23775 13680 23815 13685
rect 24310 13685 24315 13715
rect 24345 13685 24350 13715
rect 24310 13680 24350 13685
rect 24395 13715 24425 13720
rect 24395 13680 24425 13685
rect 24440 13905 24525 13920
rect 24540 13940 24570 13945
rect 24540 13905 24570 13910
rect 24440 13680 24455 13905
rect 24600 13890 24615 15225
rect 24645 13915 24660 15295
rect 26035 15300 26040 15330
rect 26070 15300 26075 15330
rect 26035 15295 26075 15300
rect 25855 15190 25895 15195
rect 24710 15155 24715 15185
rect 24745 15155 24750 15185
rect 24680 15085 24685 15115
rect 24715 15085 24720 15115
rect 24500 13875 24615 13890
rect 24630 13910 24660 13915
rect 24630 13875 24660 13880
rect 24500 13680 24515 13875
rect 24690 13860 24705 15085
rect 24735 13885 24750 15155
rect 25855 15160 25860 15190
rect 25890 15160 25895 15190
rect 25855 15155 25895 15160
rect 24800 15015 24805 15045
rect 24835 15015 24840 15045
rect 24770 14945 24775 14975
rect 24805 14945 24810 14975
rect 24560 13845 24705 13860
rect 24720 13880 24750 13885
rect 24720 13845 24750 13850
rect 24560 13680 24575 13845
rect 24780 13830 24795 14945
rect 24825 13855 24840 15015
rect 24980 14875 24985 14905
rect 25015 14875 25020 14905
rect 24950 14805 24955 14835
rect 24985 14805 24990 14835
rect 24890 14735 24895 14765
rect 24925 14735 24930 14765
rect 24860 14665 24865 14695
rect 24895 14665 24900 14695
rect 24620 13815 24795 13830
rect 24810 13850 24840 13855
rect 24810 13815 24840 13820
rect 24620 13680 24635 13815
rect 24870 13800 24885 14665
rect 24915 13825 24930 14735
rect 24680 13785 24885 13800
rect 24900 13820 24930 13825
rect 24900 13785 24930 13790
rect 24680 13680 24695 13785
rect 24960 13770 24975 14805
rect 25005 13795 25020 14875
rect 25855 13855 25870 15155
rect 25885 15120 25925 15125
rect 25885 15090 25890 15120
rect 25920 15090 25925 15120
rect 25885 15085 25925 15090
rect 25855 13850 25885 13855
rect 25855 13815 25885 13820
rect 25900 13830 25915 15085
rect 25945 15050 25985 15055
rect 25945 15020 25950 15050
rect 25980 15020 25985 15050
rect 25945 15015 25985 15020
rect 25945 13885 25960 15015
rect 25975 14980 26015 14985
rect 25975 14950 25980 14980
rect 26010 14950 26015 14980
rect 25975 14945 26015 14950
rect 25945 13880 25975 13885
rect 25945 13845 25975 13850
rect 25990 13860 26005 14945
rect 26035 13915 26050 15295
rect 26065 15260 26105 15265
rect 26065 15230 26070 15260
rect 26100 15230 26105 15260
rect 26065 15225 26105 15230
rect 26035 13910 26065 13915
rect 26035 13875 26065 13880
rect 26080 13890 26095 15225
rect 26125 13945 26140 15435
rect 26155 15400 26195 15405
rect 26155 15370 26160 15400
rect 26190 15370 26195 15400
rect 26155 15365 26195 15370
rect 26995 15365 27000 15395
rect 27030 15365 27035 15395
rect 26125 13940 26155 13945
rect 26125 13905 26155 13910
rect 26170 13920 26185 15365
rect 26805 14210 26845 14215
rect 26805 14180 26810 14210
rect 26840 14180 26845 14210
rect 26805 14175 26845 14180
rect 26880 14175 26885 14205
rect 26915 14175 26920 14205
rect 26270 14140 26310 14145
rect 26270 14110 26275 14140
rect 26305 14110 26310 14140
rect 26270 14105 26310 14110
rect 26170 13905 26255 13920
rect 26080 13875 26195 13890
rect 25990 13845 26135 13860
rect 25900 13815 26075 13830
rect 24740 13755 24975 13770
rect 24990 13790 25020 13795
rect 24990 13755 25020 13760
rect 24740 13680 24755 13755
rect 26060 13680 26075 13815
rect 26120 13680 26135 13845
rect 26180 13680 26195 13875
rect 26240 13680 26255 13905
rect 26270 13715 26305 14105
rect 26810 13720 26845 14175
rect 26905 13720 26920 14175
rect 27005 13920 27020 15365
rect 27050 13945 27065 15435
rect 28620 15440 28625 15470
rect 28655 15440 28660 15470
rect 31115 15470 31155 15475
rect 28620 15435 28660 15440
rect 29520 15435 29525 15465
rect 29555 15435 29560 15465
rect 28530 15330 28570 15335
rect 27115 15295 27120 15325
rect 27150 15295 27155 15325
rect 27085 15225 27090 15255
rect 27120 15225 27125 15255
rect 26805 13715 26845 13720
rect 26270 13685 26275 13715
rect 26305 13685 26310 13715
rect 26270 13680 26310 13685
rect 26805 13685 26810 13715
rect 26840 13685 26845 13715
rect 26805 13680 26845 13685
rect 26890 13715 26920 13720
rect 26890 13680 26920 13685
rect 26935 13905 27020 13920
rect 27035 13940 27065 13945
rect 27035 13905 27065 13910
rect 26935 13680 26950 13905
rect 27095 13890 27110 15225
rect 27140 13915 27155 15295
rect 28530 15300 28535 15330
rect 28565 15300 28570 15330
rect 28530 15295 28570 15300
rect 28350 15190 28390 15195
rect 27295 15155 27300 15185
rect 27330 15155 27335 15185
rect 27265 15085 27270 15115
rect 27300 15085 27305 15115
rect 27205 15015 27210 15045
rect 27240 15015 27245 15045
rect 27175 14945 27180 14975
rect 27210 14945 27215 14975
rect 26995 13875 27110 13890
rect 27125 13910 27155 13915
rect 27125 13875 27155 13880
rect 26995 13680 27010 13875
rect 27185 13860 27200 14945
rect 27230 13885 27245 15015
rect 27055 13845 27200 13860
rect 27215 13880 27245 13885
rect 27215 13845 27245 13850
rect 27055 13680 27070 13845
rect 27275 13830 27290 15085
rect 27320 13855 27335 15155
rect 27115 13815 27290 13830
rect 27305 13850 27335 13855
rect 27305 13815 27335 13820
rect 28350 15160 28355 15190
rect 28385 15160 28390 15190
rect 28350 15155 28390 15160
rect 28350 13855 28365 15155
rect 28380 15120 28420 15125
rect 28380 15090 28385 15120
rect 28415 15090 28420 15120
rect 28380 15085 28420 15090
rect 28350 13850 28380 13855
rect 28350 13815 28380 13820
rect 28395 13830 28410 15085
rect 28440 15050 28480 15055
rect 28440 15020 28445 15050
rect 28475 15020 28480 15050
rect 28440 15015 28480 15020
rect 28440 13885 28455 15015
rect 28470 14980 28510 14985
rect 28470 14950 28475 14980
rect 28505 14950 28510 14980
rect 28470 14945 28510 14950
rect 28440 13880 28470 13885
rect 28440 13845 28470 13850
rect 28485 13860 28500 14945
rect 28530 13915 28545 15295
rect 28560 15260 28600 15265
rect 28560 15230 28565 15260
rect 28595 15230 28600 15260
rect 28560 15225 28600 15230
rect 28530 13910 28560 13915
rect 28530 13875 28560 13880
rect 28575 13890 28590 15225
rect 28620 13945 28635 15435
rect 28650 15400 28690 15405
rect 28650 15370 28655 15400
rect 28685 15370 28690 15400
rect 28650 15365 28690 15370
rect 29490 15365 29495 15395
rect 29525 15365 29530 15395
rect 28620 13940 28650 13945
rect 28620 13905 28650 13910
rect 28665 13920 28680 15365
rect 29300 14210 29340 14215
rect 29300 14180 29305 14210
rect 29335 14180 29340 14210
rect 29300 14175 29340 14180
rect 29375 14175 29380 14205
rect 29410 14175 29415 14205
rect 28765 14140 28805 14145
rect 28765 14110 28770 14140
rect 28800 14110 28805 14140
rect 28765 14105 28805 14110
rect 28665 13905 28750 13920
rect 28575 13875 28690 13890
rect 28485 13845 28630 13860
rect 28395 13815 28570 13830
rect 27115 13680 27130 13815
rect 28555 13680 28570 13815
rect 28615 13680 28630 13845
rect 28675 13680 28690 13875
rect 28735 13680 28750 13905
rect 28765 13715 28800 14105
rect 29305 13720 29340 14175
rect 29400 13720 29415 14175
rect 29500 13920 29515 15365
rect 29545 13945 29560 15435
rect 31115 15440 31120 15470
rect 31150 15440 31155 15470
rect 33610 15470 33650 15475
rect 31115 15435 31155 15440
rect 32015 15435 32020 15465
rect 32050 15435 32055 15465
rect 31025 15330 31065 15335
rect 29610 15295 29615 15325
rect 29645 15295 29650 15325
rect 29580 15225 29585 15255
rect 29615 15225 29620 15255
rect 29300 13715 29340 13720
rect 28765 13685 28770 13715
rect 28800 13685 28805 13715
rect 28765 13680 28805 13685
rect 29300 13685 29305 13715
rect 29335 13685 29340 13715
rect 29300 13680 29340 13685
rect 29385 13715 29415 13720
rect 29385 13680 29415 13685
rect 29430 13905 29515 13920
rect 29530 13940 29560 13945
rect 29530 13905 29560 13910
rect 29430 13680 29445 13905
rect 29590 13890 29605 15225
rect 29635 13915 29650 15295
rect 31025 15300 31030 15330
rect 31060 15300 31065 15330
rect 31025 15295 31065 15300
rect 29790 15155 29795 15185
rect 29825 15155 29830 15185
rect 29760 15085 29765 15115
rect 29795 15085 29800 15115
rect 29700 15015 29705 15045
rect 29735 15015 29740 15045
rect 29670 14945 29675 14975
rect 29705 14945 29710 14975
rect 29490 13875 29605 13890
rect 29620 13910 29650 13915
rect 29620 13875 29650 13880
rect 29490 13680 29505 13875
rect 29680 13860 29695 14945
rect 29725 13885 29740 15015
rect 29550 13845 29695 13860
rect 29710 13880 29740 13885
rect 29710 13845 29740 13850
rect 29550 13680 29565 13845
rect 29770 13830 29785 15085
rect 29815 13855 29830 15155
rect 31025 13915 31040 15295
rect 31055 15260 31095 15265
rect 31055 15230 31060 15260
rect 31090 15230 31095 15260
rect 31055 15225 31095 15230
rect 31025 13910 31055 13915
rect 31025 13875 31055 13880
rect 31070 13890 31085 15225
rect 31115 13945 31130 15435
rect 31145 15400 31185 15405
rect 31145 15370 31150 15400
rect 31180 15370 31185 15400
rect 31145 15365 31185 15370
rect 31985 15365 31990 15395
rect 32020 15365 32025 15395
rect 31115 13940 31145 13945
rect 31115 13905 31145 13910
rect 31160 13920 31175 15365
rect 31795 14210 31835 14215
rect 31795 14180 31800 14210
rect 31830 14180 31835 14210
rect 31795 14175 31835 14180
rect 31870 14175 31875 14205
rect 31905 14175 31910 14205
rect 31260 14140 31300 14145
rect 31260 14110 31265 14140
rect 31295 14110 31300 14140
rect 31260 14105 31300 14110
rect 31160 13905 31245 13920
rect 31070 13875 31185 13890
rect 29610 13815 29785 13830
rect 29800 13850 29830 13855
rect 29800 13815 29830 13820
rect 29610 13680 29625 13815
rect 31170 13680 31185 13875
rect 31230 13680 31245 13905
rect 31260 13715 31295 14105
rect 31800 13720 31835 14175
rect 31895 13720 31910 14175
rect 31995 13920 32010 15365
rect 32040 13945 32055 15435
rect 33610 15440 33615 15470
rect 33645 15440 33650 15470
rect 36105 15470 36145 15475
rect 33610 15435 33650 15440
rect 34510 15435 34515 15465
rect 34545 15435 34550 15465
rect 33520 15330 33560 15335
rect 32105 15295 32110 15325
rect 32140 15295 32145 15325
rect 32075 15225 32080 15255
rect 32110 15225 32115 15255
rect 31795 13715 31835 13720
rect 31260 13685 31265 13715
rect 31295 13685 31300 13715
rect 31260 13680 31300 13685
rect 31795 13685 31800 13715
rect 31830 13685 31835 13715
rect 31795 13680 31835 13685
rect 31880 13715 31910 13720
rect 31880 13680 31910 13685
rect 31925 13905 32010 13920
rect 32025 13940 32055 13945
rect 32025 13905 32055 13910
rect 31925 13680 31940 13905
rect 32085 13890 32100 15225
rect 32130 13915 32145 15295
rect 31985 13875 32100 13890
rect 32115 13910 32145 13915
rect 32115 13875 32145 13880
rect 33520 15300 33525 15330
rect 33555 15300 33560 15330
rect 33520 15295 33560 15300
rect 33520 13915 33535 15295
rect 33550 15260 33590 15265
rect 33550 15230 33555 15260
rect 33585 15230 33590 15260
rect 33550 15225 33590 15230
rect 33520 13910 33550 13915
rect 33520 13875 33550 13880
rect 33565 13890 33580 15225
rect 33610 13945 33625 15435
rect 33640 15400 33680 15405
rect 33640 15370 33645 15400
rect 33675 15370 33680 15400
rect 33640 15365 33680 15370
rect 34480 15365 34485 15395
rect 34515 15365 34520 15395
rect 33610 13940 33640 13945
rect 33610 13905 33640 13910
rect 33655 13920 33670 15365
rect 34290 14210 34330 14215
rect 34290 14180 34295 14210
rect 34325 14180 34330 14210
rect 34290 14175 34330 14180
rect 34365 14175 34370 14205
rect 34400 14175 34405 14205
rect 33755 14140 33795 14145
rect 33755 14110 33760 14140
rect 33790 14110 33795 14140
rect 33755 14105 33795 14110
rect 33655 13905 33740 13920
rect 33565 13875 33680 13890
rect 31985 13680 32000 13875
rect 33665 13680 33680 13875
rect 33725 13680 33740 13905
rect 33755 13715 33790 14105
rect 34295 13720 34330 14175
rect 34390 13720 34405 14175
rect 34490 13920 34505 15365
rect 34535 13945 34550 15435
rect 36105 15440 36110 15470
rect 36140 15440 36145 15470
rect 38600 15470 38640 15475
rect 36105 15435 36145 15440
rect 37005 15435 37010 15465
rect 37040 15435 37045 15465
rect 34600 15295 34605 15325
rect 34635 15295 34640 15325
rect 34570 15225 34575 15255
rect 34605 15225 34610 15255
rect 34290 13715 34330 13720
rect 33755 13685 33760 13715
rect 33790 13685 33795 13715
rect 33755 13680 33795 13685
rect 34290 13685 34295 13715
rect 34325 13685 34330 13715
rect 34290 13680 34330 13685
rect 34375 13715 34405 13720
rect 34375 13680 34405 13685
rect 34420 13905 34505 13920
rect 34520 13940 34550 13945
rect 34520 13905 34550 13910
rect 34420 13680 34435 13905
rect 34580 13890 34595 15225
rect 34625 13915 34640 15295
rect 34480 13875 34595 13890
rect 34610 13910 34640 13915
rect 36105 13945 36120 15435
rect 36135 15400 36175 15405
rect 36135 15370 36140 15400
rect 36170 15370 36175 15400
rect 36135 15365 36175 15370
rect 36975 15365 36980 15395
rect 37010 15365 37015 15395
rect 36105 13940 36135 13945
rect 36105 13905 36135 13910
rect 36150 13920 36165 15365
rect 36785 14210 36825 14215
rect 36785 14180 36790 14210
rect 36820 14180 36825 14210
rect 36785 14175 36825 14180
rect 36860 14175 36865 14205
rect 36895 14175 36900 14205
rect 36250 14140 36290 14145
rect 36250 14110 36255 14140
rect 36285 14110 36290 14140
rect 36250 14105 36290 14110
rect 36150 13905 36235 13920
rect 34610 13875 34640 13880
rect 34480 13680 34495 13875
rect 36220 13680 36235 13905
rect 36250 13715 36285 14105
rect 36790 13720 36825 14175
rect 36885 13720 36900 14175
rect 36985 13920 37000 15365
rect 37030 13945 37045 15435
rect 36785 13715 36825 13720
rect 36250 13685 36255 13715
rect 36285 13685 36290 13715
rect 36250 13680 36290 13685
rect 36785 13685 36790 13715
rect 36820 13685 36825 13715
rect 36785 13680 36825 13685
rect 36870 13715 36900 13720
rect 36870 13680 36900 13685
rect 36915 13905 37000 13920
rect 37015 13940 37045 13945
rect 37015 13905 37045 13910
rect 38600 15440 38605 15470
rect 38635 15440 38640 15470
rect 38600 15435 38640 15440
rect 39500 15435 39505 15465
rect 39535 15435 39540 15465
rect 38600 13945 38615 15435
rect 38630 15400 38670 15405
rect 38630 15370 38635 15400
rect 38665 15370 38670 15400
rect 38630 15365 38670 15370
rect 39470 15365 39475 15395
rect 39505 15365 39510 15395
rect 38600 13940 38630 13945
rect 38600 13905 38630 13910
rect 38645 13920 38660 15365
rect 39280 14210 39320 14215
rect 39280 14180 39285 14210
rect 39315 14180 39320 14210
rect 39280 14175 39320 14180
rect 39355 14175 39360 14205
rect 39390 14175 39395 14205
rect 38745 14140 38785 14145
rect 38745 14110 38750 14140
rect 38780 14110 38785 14140
rect 38745 14105 38785 14110
rect 38645 13905 38730 13920
rect 36915 13680 36930 13905
rect 38715 13680 38730 13905
rect 38745 13715 38780 14105
rect 39285 13720 39320 14175
rect 39380 13720 39395 14175
rect 39480 13920 39495 15365
rect 39525 13945 39540 15435
rect 39280 13715 39320 13720
rect 38745 13685 38750 13715
rect 38780 13685 38785 13715
rect 38745 13680 38785 13685
rect 39280 13685 39285 13715
rect 39315 13685 39320 13715
rect 39280 13680 39320 13685
rect 39365 13715 39395 13720
rect 39365 13680 39395 13685
rect 39410 13905 39495 13920
rect 39510 13940 39540 13945
rect 39510 13905 39540 13910
rect 39410 13680 39425 13905
<< via2 >>
rect 1180 15440 1210 15470
rect 1210 15370 1240 15400
rect 1860 14180 1890 14210
rect 1325 14110 1355 14140
rect 3675 15440 3705 15470
rect 3705 15370 3735 15400
rect 4355 14180 4385 14210
rect 3820 14110 3850 14140
rect 6170 15440 6200 15470
rect 6080 15300 6110 15330
rect 6110 15230 6140 15260
rect 6200 15370 6230 15400
rect 6850 14180 6880 14210
rect 6315 14110 6345 14140
rect 8665 15440 8695 15470
rect 8575 15300 8605 15330
rect 8605 15230 8635 15260
rect 8695 15370 8725 15400
rect 9345 14180 9375 14210
rect 8810 14110 8840 14140
rect 11160 15440 11190 15470
rect 11070 15300 11100 15330
rect 10890 15160 10920 15190
rect 10920 15090 10950 15120
rect 10980 15020 11010 15050
rect 11010 14950 11040 14980
rect 11100 15230 11130 15260
rect 11190 15370 11220 15400
rect 11840 14180 11870 14210
rect 11305 14110 11335 14140
rect 13655 15440 13685 15470
rect 13565 15300 13595 15330
rect 13385 15160 13415 15190
rect 13415 15090 13445 15120
rect 13475 15020 13505 15050
rect 13505 14950 13535 14980
rect 13595 15230 13625 15260
rect 13685 15370 13715 15400
rect 14335 14180 14365 14210
rect 13800 14110 13830 14140
rect 16150 15440 16180 15470
rect 16060 15300 16090 15330
rect 15970 15160 16000 15190
rect 15880 15020 15910 15050
rect 15700 14880 15730 14910
rect 15730 14810 15760 14840
rect 15790 14740 15820 14770
rect 15820 14670 15850 14700
rect 15910 14950 15940 14980
rect 16000 15090 16030 15120
rect 16090 15230 16120 15260
rect 16180 15370 16210 15400
rect 16830 14180 16860 14210
rect 16295 14110 16325 14140
rect 18645 15440 18675 15470
rect 18555 15300 18585 15330
rect 18465 15160 18495 15190
rect 18375 15020 18405 15050
rect 18285 14880 18315 14910
rect 18195 14600 18225 14630
rect 18105 14320 18135 14350
rect 18135 14250 18165 14280
rect 18225 14530 18255 14560
rect 18315 14810 18345 14840
rect 18405 14950 18435 14980
rect 18495 15090 18525 15120
rect 18585 15230 18615 15260
rect 18675 15370 18705 15400
rect 19325 14180 19355 14210
rect 18790 14110 18820 14140
rect 21140 15440 21170 15470
rect 21050 15300 21080 15330
rect 20960 15160 20990 15190
rect 20870 15020 20900 15050
rect 20780 14880 20810 14910
rect 20600 14600 20630 14630
rect 20630 14530 20660 14560
rect 20675 14460 20705 14490
rect 20720 14390 20750 14420
rect 20810 14810 20840 14840
rect 20900 14950 20930 14980
rect 20990 15090 21020 15120
rect 21080 15230 21110 15260
rect 21170 15370 21200 15400
rect 21820 14180 21850 14210
rect 21285 14110 21315 14140
rect 23635 15440 23665 15470
rect 23545 15300 23575 15330
rect 23455 15160 23485 15190
rect 23365 15020 23395 15050
rect 23185 14880 23215 14910
rect 23215 14810 23245 14840
rect 23275 14740 23305 14770
rect 23305 14670 23335 14700
rect 23395 14950 23425 14980
rect 23485 15090 23515 15120
rect 23575 15230 23605 15260
rect 23665 15370 23695 15400
rect 24315 14180 24345 14210
rect 23780 14110 23810 14140
rect 26130 15440 26160 15470
rect 26040 15300 26070 15330
rect 25860 15160 25890 15190
rect 25890 15090 25920 15120
rect 25950 15020 25980 15050
rect 25980 14950 26010 14980
rect 26070 15230 26100 15260
rect 26160 15370 26190 15400
rect 26810 14180 26840 14210
rect 26275 14110 26305 14140
rect 28625 15440 28655 15470
rect 28535 15300 28565 15330
rect 28355 15160 28385 15190
rect 28385 15090 28415 15120
rect 28445 15020 28475 15050
rect 28475 14950 28505 14980
rect 28565 15230 28595 15260
rect 28655 15370 28685 15400
rect 29305 14180 29335 14210
rect 28770 14110 28800 14140
rect 31120 15440 31150 15470
rect 31030 15300 31060 15330
rect 31060 15230 31090 15260
rect 31150 15370 31180 15400
rect 31800 14180 31830 14210
rect 31265 14110 31295 14140
rect 33615 15440 33645 15470
rect 33525 15300 33555 15330
rect 33555 15230 33585 15260
rect 33645 15370 33675 15400
rect 34295 14180 34325 14210
rect 33760 14110 33790 14140
rect 36110 15440 36140 15470
rect 36140 15370 36170 15400
rect 36790 14180 36820 14210
rect 36255 14110 36285 14140
rect 38605 15440 38635 15470
rect 38635 15370 38665 15400
rect 39285 14180 39315 14210
rect 38750 14110 38780 14140
<< metal3 >>
rect 1175 15470 1215 15475
rect -33 15465 36 15468
rect 1175 15465 1180 15470
rect -33 15440 1180 15465
rect 1210 15465 1215 15470
rect 3670 15470 3710 15475
rect 3670 15465 3675 15470
rect 1210 15440 3675 15465
rect 3705 15465 3710 15470
rect 6165 15470 6205 15475
rect 6165 15465 6170 15470
rect 3705 15440 6170 15465
rect 6200 15465 6205 15470
rect 8660 15470 8700 15475
rect 8660 15465 8665 15470
rect 6200 15440 8665 15465
rect 8695 15465 8700 15470
rect 11155 15470 11195 15475
rect 11155 15465 11160 15470
rect 8695 15440 11160 15465
rect 11190 15465 11195 15470
rect 13650 15470 13690 15475
rect 13650 15465 13655 15470
rect 11190 15440 13655 15465
rect 13685 15465 13690 15470
rect 16145 15470 16185 15475
rect 16145 15465 16150 15470
rect 13685 15440 16150 15465
rect 16180 15465 16185 15470
rect 18640 15470 18680 15475
rect 18640 15465 18645 15470
rect 16180 15440 18645 15465
rect 18675 15465 18680 15470
rect 21135 15470 21175 15475
rect 21135 15465 21140 15470
rect 18675 15440 21140 15465
rect 21170 15465 21175 15470
rect 23630 15470 23670 15475
rect 23630 15465 23635 15470
rect 21170 15440 23635 15465
rect 23665 15465 23670 15470
rect 26125 15470 26165 15475
rect 26125 15465 26130 15470
rect 23665 15440 26130 15465
rect 26160 15465 26165 15470
rect 28620 15470 28660 15475
rect 28620 15465 28625 15470
rect 26160 15440 28625 15465
rect 28655 15465 28660 15470
rect 31115 15470 31155 15475
rect 31115 15465 31120 15470
rect 28655 15440 31120 15465
rect 31150 15465 31155 15470
rect 33610 15470 33650 15475
rect 33610 15465 33615 15470
rect 31150 15440 33615 15465
rect 33645 15465 33650 15470
rect 36105 15470 36145 15475
rect 36105 15465 36110 15470
rect 33645 15440 36110 15465
rect 36140 15465 36145 15470
rect 38600 15470 38640 15475
rect 38600 15465 38605 15470
rect 36140 15440 38605 15465
rect 38635 15465 38640 15470
rect 38635 15440 39850 15465
rect -33 15435 39850 15440
rect 1205 15400 1245 15405
rect 1205 15395 1210 15400
rect -31 15370 1210 15395
rect 1240 15395 1245 15400
rect 3700 15400 3740 15405
rect 3700 15395 3705 15400
rect 1240 15370 3705 15395
rect 3735 15395 3740 15400
rect 6195 15400 6235 15405
rect 6195 15395 6200 15400
rect 3735 15370 6200 15395
rect 6230 15395 6235 15400
rect 8690 15400 8730 15405
rect 8690 15395 8695 15400
rect 6230 15370 8695 15395
rect 8725 15395 8730 15400
rect 11185 15400 11225 15405
rect 11185 15395 11190 15400
rect 8725 15370 11190 15395
rect 11220 15395 11225 15400
rect 13680 15400 13720 15405
rect 13680 15395 13685 15400
rect 11220 15370 13685 15395
rect 13715 15395 13720 15400
rect 16175 15400 16215 15405
rect 16175 15395 16180 15400
rect 13715 15370 16180 15395
rect 16210 15395 16215 15400
rect 18670 15400 18710 15405
rect 18670 15395 18675 15400
rect 16210 15370 18675 15395
rect 18705 15395 18710 15400
rect 21165 15400 21205 15405
rect 21165 15395 21170 15400
rect 18705 15370 21170 15395
rect 21200 15395 21205 15400
rect 23660 15400 23700 15405
rect 23660 15395 23665 15400
rect 21200 15370 23665 15395
rect 23695 15395 23700 15400
rect 26155 15400 26195 15405
rect 26155 15395 26160 15400
rect 23695 15370 26160 15395
rect 26190 15395 26195 15400
rect 28650 15400 28690 15405
rect 28650 15395 28655 15400
rect 26190 15370 28655 15395
rect 28685 15395 28690 15400
rect 31145 15400 31185 15405
rect 31145 15395 31150 15400
rect 28685 15370 31150 15395
rect 31180 15395 31185 15400
rect 33640 15400 33680 15405
rect 33640 15395 33645 15400
rect 31180 15370 33645 15395
rect 33675 15395 33680 15400
rect 36135 15400 36175 15405
rect 36135 15395 36140 15400
rect 33675 15370 36140 15395
rect 36170 15395 36175 15400
rect 38630 15400 38670 15405
rect 38630 15395 38635 15400
rect 36170 15370 38635 15395
rect 38665 15395 38670 15400
rect 38665 15370 39850 15395
rect -31 15365 39850 15370
rect -31 15362 38 15365
rect 6075 15330 6115 15335
rect 6075 15325 6080 15330
rect -30 15300 6080 15325
rect 6110 15325 6115 15330
rect 8570 15330 8610 15335
rect 8570 15325 8575 15330
rect 6110 15300 8575 15325
rect 8605 15325 8610 15330
rect 11065 15330 11105 15335
rect 11065 15325 11070 15330
rect 8605 15300 11070 15325
rect 11100 15325 11105 15330
rect 13560 15330 13600 15335
rect 13560 15325 13565 15330
rect 11100 15300 13565 15325
rect 13595 15325 13600 15330
rect 16055 15330 16095 15335
rect 16055 15325 16060 15330
rect 13595 15300 16060 15325
rect 16090 15325 16095 15330
rect 18550 15330 18590 15335
rect 18550 15325 18555 15330
rect 16090 15300 18555 15325
rect 18585 15325 18590 15330
rect 21045 15330 21085 15335
rect 21045 15325 21050 15330
rect 18585 15300 21050 15325
rect 21080 15325 21085 15330
rect 23540 15330 23580 15335
rect 23540 15325 23545 15330
rect 21080 15300 23545 15325
rect 23575 15325 23580 15330
rect 26035 15330 26075 15335
rect 26035 15325 26040 15330
rect 23575 15300 26040 15325
rect 26070 15325 26075 15330
rect 28530 15330 28570 15335
rect 28530 15325 28535 15330
rect 26070 15300 28535 15325
rect 28565 15325 28570 15330
rect 31025 15330 31065 15335
rect 31025 15325 31030 15330
rect 28565 15300 31030 15325
rect 31060 15325 31065 15330
rect 33520 15330 33560 15335
rect 33520 15325 33525 15330
rect 31060 15300 33525 15325
rect 33555 15325 33560 15330
rect 33555 15300 39850 15325
rect -30 15295 39850 15300
rect -29 15291 40 15295
rect 6105 15260 6145 15265
rect -31 15255 38 15256
rect 6105 15255 6110 15260
rect -31 15230 6110 15255
rect 6140 15255 6145 15260
rect 8600 15260 8640 15265
rect 8600 15255 8605 15260
rect 6140 15230 8605 15255
rect 8635 15255 8640 15260
rect 11095 15260 11135 15265
rect 11095 15255 11100 15260
rect 8635 15230 11100 15255
rect 11130 15255 11135 15260
rect 13590 15260 13630 15265
rect 13590 15255 13595 15260
rect 11130 15230 13595 15255
rect 13625 15255 13630 15260
rect 16085 15260 16125 15265
rect 16085 15255 16090 15260
rect 13625 15230 16090 15255
rect 16120 15255 16125 15260
rect 18580 15260 18620 15265
rect 18580 15255 18585 15260
rect 16120 15230 18585 15255
rect 18615 15255 18620 15260
rect 21075 15260 21115 15265
rect 21075 15255 21080 15260
rect 18615 15230 21080 15255
rect 21110 15255 21115 15260
rect 23570 15260 23610 15265
rect 23570 15255 23575 15260
rect 21110 15230 23575 15255
rect 23605 15255 23610 15260
rect 26065 15260 26105 15265
rect 26065 15255 26070 15260
rect 23605 15230 26070 15255
rect 26100 15255 26105 15260
rect 28560 15260 28600 15265
rect 28560 15255 28565 15260
rect 26100 15230 28565 15255
rect 28595 15255 28600 15260
rect 31055 15260 31095 15265
rect 31055 15255 31060 15260
rect 28595 15230 31060 15255
rect 31090 15255 31095 15260
rect 33550 15260 33590 15265
rect 33550 15255 33555 15260
rect 31090 15230 33555 15255
rect 33585 15255 33590 15260
rect 33585 15230 39850 15255
rect -31 15225 39850 15230
rect -31 15223 38 15225
rect 10885 15190 10925 15195
rect 10885 15185 10890 15190
rect -32 15160 10890 15185
rect 10920 15185 10925 15190
rect 13380 15190 13420 15195
rect 13380 15185 13385 15190
rect 10920 15160 13385 15185
rect 13415 15185 13420 15190
rect 15965 15190 16005 15195
rect 15965 15185 15970 15190
rect 13415 15160 15970 15185
rect 16000 15185 16005 15190
rect 18460 15190 18500 15195
rect 18460 15185 18465 15190
rect 16000 15160 18465 15185
rect 18495 15185 18500 15190
rect 20955 15190 20995 15195
rect 20955 15185 20960 15190
rect 18495 15160 20960 15185
rect 20990 15185 20995 15190
rect 23450 15190 23490 15195
rect 23450 15185 23455 15190
rect 20990 15160 23455 15185
rect 23485 15185 23490 15190
rect 25855 15190 25895 15195
rect 25855 15185 25860 15190
rect 23485 15160 25860 15185
rect 25890 15185 25895 15190
rect 28350 15190 28390 15195
rect 28350 15185 28355 15190
rect 25890 15160 28355 15185
rect 28385 15185 28390 15190
rect 28385 15160 39850 15185
rect -32 15155 39850 15160
rect -32 15152 37 15155
rect 10915 15120 10955 15125
rect 10915 15115 10920 15120
rect -32 15090 10920 15115
rect 10950 15115 10955 15120
rect 13410 15120 13450 15125
rect 13410 15115 13415 15120
rect 10950 15090 13415 15115
rect 13445 15115 13450 15120
rect 15995 15120 16035 15125
rect 15995 15115 16000 15120
rect 13445 15090 16000 15115
rect 16030 15115 16035 15120
rect 18490 15120 18530 15125
rect 18490 15115 18495 15120
rect 16030 15090 18495 15115
rect 18525 15115 18530 15120
rect 20985 15120 21025 15125
rect 20985 15115 20990 15120
rect 18525 15090 20990 15115
rect 21020 15115 21025 15120
rect 23480 15120 23520 15125
rect 23480 15115 23485 15120
rect 21020 15090 23485 15115
rect 23515 15115 23520 15120
rect 25885 15120 25925 15125
rect 25885 15115 25890 15120
rect 23515 15090 25890 15115
rect 25920 15115 25925 15120
rect 28380 15120 28420 15125
rect 28380 15115 28385 15120
rect 25920 15090 28385 15115
rect 28415 15115 28420 15120
rect 28415 15090 39850 15115
rect -32 15085 39850 15090
rect -32 15082 37 15085
rect 10975 15050 11015 15055
rect -35 15045 34 15046
rect 10975 15045 10980 15050
rect -35 15020 10980 15045
rect 11010 15045 11015 15050
rect 13470 15050 13510 15055
rect 13470 15045 13475 15050
rect 11010 15020 13475 15045
rect 13505 15045 13510 15050
rect 15875 15050 15915 15055
rect 15875 15045 15880 15050
rect 13505 15020 15880 15045
rect 15910 15045 15915 15050
rect 18370 15050 18410 15055
rect 18370 15045 18375 15050
rect 15910 15020 18375 15045
rect 18405 15045 18410 15050
rect 20865 15050 20905 15055
rect 20865 15045 20870 15050
rect 18405 15020 20870 15045
rect 20900 15045 20905 15050
rect 23360 15050 23400 15055
rect 23360 15045 23365 15050
rect 20900 15020 23365 15045
rect 23395 15045 23400 15050
rect 25945 15050 25985 15055
rect 25945 15045 25950 15050
rect 23395 15020 25950 15045
rect 25980 15045 25985 15050
rect 28440 15050 28480 15055
rect 28440 15045 28445 15050
rect 25980 15020 28445 15045
rect 28475 15045 28480 15050
rect 28475 15020 39850 15045
rect -35 15015 39850 15020
rect -35 15013 34 15015
rect 11005 14980 11045 14985
rect -31 14975 38 14979
rect 11005 14975 11010 14980
rect -31 14950 11010 14975
rect 11040 14975 11045 14980
rect 13500 14980 13540 14985
rect 13500 14975 13505 14980
rect 11040 14950 13505 14975
rect 13535 14975 13540 14980
rect 15905 14980 15945 14985
rect 15905 14975 15910 14980
rect 13535 14950 15910 14975
rect 15940 14975 15945 14980
rect 18400 14980 18440 14985
rect 18400 14975 18405 14980
rect 15940 14950 18405 14975
rect 18435 14975 18440 14980
rect 20895 14980 20935 14985
rect 20895 14975 20900 14980
rect 18435 14950 20900 14975
rect 20930 14975 20935 14980
rect 23390 14980 23430 14985
rect 23390 14975 23395 14980
rect 20930 14950 23395 14975
rect 23425 14975 23430 14980
rect 25975 14980 26015 14985
rect 25975 14975 25980 14980
rect 23425 14950 25980 14975
rect 26010 14975 26015 14980
rect 28470 14980 28510 14985
rect 28470 14975 28475 14980
rect 26010 14950 28475 14975
rect 28505 14975 28510 14980
rect 28505 14950 39850 14975
rect -31 14946 39850 14950
rect -30 14945 39850 14946
rect 15695 14910 15735 14915
rect 15695 14905 15700 14910
rect -30 14904 15700 14905
rect -32 14880 15700 14904
rect 15730 14905 15735 14910
rect 18280 14910 18320 14915
rect 18280 14905 18285 14910
rect 15730 14880 18285 14905
rect 18315 14905 18320 14910
rect 20775 14910 20815 14915
rect 20775 14905 20780 14910
rect 18315 14880 20780 14905
rect 20810 14905 20815 14910
rect 23180 14910 23220 14915
rect 23180 14905 23185 14910
rect 20810 14880 23185 14905
rect 23215 14905 23220 14910
rect 23215 14880 39850 14905
rect -32 14875 39850 14880
rect -32 14871 37 14875
rect 15725 14840 15765 14845
rect 15725 14835 15730 14840
rect -31 14810 15730 14835
rect 15760 14835 15765 14840
rect 18310 14840 18350 14845
rect 18310 14835 18315 14840
rect 15760 14810 18315 14835
rect 18345 14835 18350 14840
rect 20805 14840 20845 14845
rect 20805 14835 20810 14840
rect 18345 14810 20810 14835
rect 20840 14835 20845 14840
rect 23210 14840 23250 14845
rect 23210 14835 23215 14840
rect 20840 14810 23215 14835
rect 23245 14835 23250 14840
rect 23245 14810 39850 14835
rect -31 14805 39850 14810
rect -31 14802 38 14805
rect 15785 14770 15825 14775
rect -32 14765 37 14768
rect 15785 14765 15790 14770
rect -32 14740 15790 14765
rect 15820 14765 15825 14770
rect 23270 14770 23310 14775
rect 23270 14765 23275 14770
rect 15820 14740 23275 14765
rect 23305 14765 23310 14770
rect 23305 14740 39850 14765
rect -32 14735 39850 14740
rect 15815 14700 15855 14705
rect 15815 14695 15820 14700
rect -30 14670 15820 14695
rect 15850 14695 15855 14700
rect 23300 14700 23340 14705
rect 23300 14695 23305 14700
rect 15850 14670 23305 14695
rect 23335 14695 23340 14700
rect 23335 14670 39850 14695
rect -30 14665 39850 14670
rect -29 14662 40 14665
rect 18190 14630 18230 14635
rect -33 14625 36 14626
rect 18190 14625 18195 14630
rect -33 14600 18195 14625
rect 18225 14625 18230 14630
rect 20595 14630 20635 14635
rect 20595 14625 20600 14630
rect 18225 14600 20600 14625
rect 20630 14625 20635 14630
rect 20630 14600 39850 14625
rect -33 14595 39850 14600
rect -33 14593 36 14595
rect 18220 14560 18260 14565
rect -31 14555 38 14557
rect 18220 14555 18225 14560
rect -31 14530 18225 14555
rect 18255 14555 18260 14560
rect 20625 14560 20665 14565
rect 20625 14555 20630 14560
rect 18255 14530 20630 14555
rect 20660 14555 20665 14560
rect 20660 14530 39850 14555
rect -31 14525 39850 14530
rect -31 14524 38 14525
rect 20670 14490 20710 14495
rect 20670 14485 20675 14490
rect -30 14460 20675 14485
rect 20705 14485 20710 14490
rect 20705 14460 39850 14485
rect -30 14455 39850 14460
rect -29 14450 40 14455
rect 20715 14420 20755 14425
rect -29 14415 40 14417
rect 20715 14415 20720 14420
rect -30 14390 20720 14415
rect 20750 14415 20755 14420
rect 20750 14390 39850 14415
rect -30 14385 39850 14390
rect -29 14384 40 14385
rect 18100 14350 18140 14355
rect 18100 14345 18105 14350
rect -30 14320 18105 14345
rect 18135 14345 18140 14350
rect 18135 14320 39850 14345
rect -30 14315 39850 14320
rect -29 14312 40 14315
rect 18130 14280 18170 14285
rect -29 14275 40 14276
rect 18130 14275 18135 14280
rect -30 14250 18135 14275
rect 18165 14275 18170 14280
rect 18165 14250 39850 14275
rect -30 14245 39850 14250
rect -29 14244 40 14245
rect 1855 14210 1895 14215
rect -30 14205 39 14207
rect 1855 14205 1860 14210
rect -30 14180 1860 14205
rect 1890 14205 1895 14210
rect 4350 14210 4390 14215
rect 4350 14205 4355 14210
rect 1890 14180 4355 14205
rect 4385 14205 4390 14210
rect 6845 14210 6885 14215
rect 6845 14205 6850 14210
rect 4385 14180 6850 14205
rect 6880 14205 6885 14210
rect 9340 14210 9380 14215
rect 9340 14205 9345 14210
rect 6880 14180 9345 14205
rect 9375 14205 9380 14210
rect 11835 14210 11875 14215
rect 11835 14205 11840 14210
rect 9375 14180 11840 14205
rect 11870 14205 11875 14210
rect 14330 14210 14370 14215
rect 14330 14205 14335 14210
rect 11870 14180 14335 14205
rect 14365 14205 14370 14210
rect 16825 14210 16865 14215
rect 16825 14205 16830 14210
rect 14365 14180 16830 14205
rect 16860 14205 16865 14210
rect 19320 14210 19360 14215
rect 19320 14205 19325 14210
rect 16860 14180 19325 14205
rect 19355 14205 19360 14210
rect 21815 14210 21855 14215
rect 21815 14205 21820 14210
rect 19355 14180 21820 14205
rect 21850 14205 21855 14210
rect 24310 14210 24350 14215
rect 24310 14205 24315 14210
rect 21850 14180 24315 14205
rect 24345 14205 24350 14210
rect 26805 14210 26845 14215
rect 26805 14205 26810 14210
rect 24345 14180 26810 14205
rect 26840 14205 26845 14210
rect 29300 14210 29340 14215
rect 29300 14205 29305 14210
rect 26840 14180 29305 14205
rect 29335 14205 29340 14210
rect 31795 14210 31835 14215
rect 31795 14205 31800 14210
rect 29335 14180 31800 14205
rect 31830 14205 31835 14210
rect 34290 14210 34330 14215
rect 34290 14205 34295 14210
rect 31830 14180 34295 14205
rect 34325 14205 34330 14210
rect 36785 14210 36825 14215
rect 36785 14205 36790 14210
rect 34325 14180 36790 14205
rect 36820 14205 36825 14210
rect 39280 14210 39320 14215
rect 39280 14205 39285 14210
rect 36820 14180 39285 14205
rect 39315 14205 39320 14210
rect 39315 14180 39850 14205
rect -30 14175 39850 14180
rect 1320 14140 1360 14145
rect 1320 14135 1325 14140
rect -30 14134 1325 14135
rect -31 14110 1325 14134
rect 1355 14135 1360 14140
rect 3815 14140 3855 14145
rect 3815 14135 3820 14140
rect 1355 14110 3820 14135
rect 3850 14135 3855 14140
rect 6310 14140 6350 14145
rect 6310 14135 6315 14140
rect 3850 14110 6315 14135
rect 6345 14135 6350 14140
rect 8805 14140 8845 14145
rect 8805 14135 8810 14140
rect 6345 14110 8810 14135
rect 8840 14135 8845 14140
rect 11300 14140 11340 14145
rect 11300 14135 11305 14140
rect 8840 14110 11305 14135
rect 11335 14135 11340 14140
rect 13795 14140 13835 14145
rect 13795 14135 13800 14140
rect 11335 14110 13800 14135
rect 13830 14135 13835 14140
rect 16290 14140 16330 14145
rect 16290 14135 16295 14140
rect 13830 14110 16295 14135
rect 16325 14135 16330 14140
rect 18785 14140 18825 14145
rect 18785 14135 18790 14140
rect 16325 14110 18790 14135
rect 18820 14135 18825 14140
rect 21280 14140 21320 14145
rect 21280 14135 21285 14140
rect 18820 14110 21285 14135
rect 21315 14135 21320 14140
rect 23775 14140 23815 14145
rect 23775 14135 23780 14140
rect 21315 14110 23780 14135
rect 23810 14135 23815 14140
rect 26270 14140 26310 14145
rect 26270 14135 26275 14140
rect 23810 14110 26275 14135
rect 26305 14135 26310 14140
rect 28765 14140 28805 14145
rect 28765 14135 28770 14140
rect 26305 14110 28770 14135
rect 28800 14135 28805 14140
rect 31260 14140 31300 14145
rect 31260 14135 31265 14140
rect 28800 14110 31265 14135
rect 31295 14135 31300 14140
rect 33755 14140 33795 14145
rect 33755 14135 33760 14140
rect 31295 14110 33760 14135
rect 33790 14135 33795 14140
rect 36250 14140 36290 14145
rect 36250 14135 36255 14140
rect 33790 14110 36255 14135
rect 36285 14135 36290 14140
rect 38745 14140 38785 14145
rect 38745 14135 38750 14140
rect 36285 14110 38750 14135
rect 38780 14135 38785 14140
rect 38780 14110 39850 14135
rect -31 14105 39850 14110
rect -31 14103 40 14105
rect -29 14102 40 14103
<< metal4 >>
rect 40 -30 70 0
rect 2535 -30 2565 0
rect 5030 -30 5060 0
rect 7525 -30 7555 0
rect 10020 -30 10050 0
rect 12515 -30 12545 0
rect 15010 -30 15040 0
rect 17505 -30 17535 0
rect 20000 -30 20030 0
rect 22495 -30 22525 0
rect 24990 -30 25020 0
rect 27485 -30 27515 0
rect 29980 -30 30010 0
rect 32475 -30 32505 0
rect 34970 -30 35000 0
rect 37465 -30 37495 0
rect 0 -60 39785 -30
use end  end_0
timestamp 1729689530
transform 0 1 0 -1 0 13680
box 0 0 13680 2360
use end  end_1
timestamp 1729689530
transform 0 1 2495 -1 0 13680
box 0 0 13680 2360
use end  end_2
timestamp 1729689530
transform 0 1 34930 -1 0 13680
box 0 0 13680 2360
use end  end_3
timestamp 1729689530
transform 0 1 37425 -1 0 13680
box 0 0 13680 2360
use mid_2  mid_2_0
timestamp 1729709358
transform 1 0 17465 0 1 6840
box 0 -6840 4900 6840
use mid_2to4_  mid_2to4__0
timestamp 1729683266
transform 0 1 14970 -1 0 13680
box 0 0 13680 2360
use mid_2to4_  mid_2to4__1
timestamp 1729683266
transform 0 1 22455 -1 0 13680
box 0 0 13680 2360
use mid_4to8  mid_4to8_0
timestamp 1729685583
transform 0 1 9980 -1 0 13680
box 0 0 13680 2360
use mid_4to8  mid_4to8_1
timestamp 1729685583
transform 0 1 12475 -1 0 13680
box 0 0 13680 2360
use mid_4to8  mid_4to8_2
timestamp 1729685583
transform 0 1 24950 -1 0 13680
box 0 0 13680 2360
use mid_4to8  mid_4to8_3
timestamp 1729685583
transform 0 1 27445 -1 0 13680
box 0 0 13680 2360
use mid_6to8  mid_6to8_0
timestamp 1729688460
transform 0 1 4990 -1 0 13680
box 0 0 13680 2360
use mid_6to8  mid_6to8_1
timestamp 1729688460
transform 0 1 7485 -1 0 13680
box 0 0 13680 2360
use mid_6to8  mid_6to8_2
timestamp 1729688460
transform 0 1 29940 -1 0 13680
box 0 0 13680 2360
use mid_6to8  mid_6to8_3
timestamp 1729688460
transform 0 1 32435 -1 0 13680
box 0 0 13680 2360
<< labels >>
flabel metal3 -31 14103 39 14134 0 FreeSans 80 0 0 0 Sub
flabel metal3 -30 14175 39 14207 0 FreeSans 80 0 0 0 Vdd
port 4 nsew
flabel metal3 -29 14244 40 14276 0 FreeSans 80 0 0 0 smpl
port 12 nsew
flabel space 66 14244 119 14260 0 FreeSans 80 0 0 0 smpl_out_n
port 14 nsew
flabel metal3 -29 14312 40 14344 0 FreeSans 80 0 0 0 smpl_n_d12
port 16 nsew
flabel metal3 -29 14384 40 14417 0 FreeSans 80 0 0 0 phi10
port 18 nsew
flabel metal3 -29 14450 40 14483 0 FreeSans 80 0 0 0 phi20
port 20 nsew
flabel metal3 -31 14524 38 14557 0 FreeSans 80 0 0 0 phi11
port 22 nsew
flabel metal3 -33 14593 36 14626 0 FreeSans 80 0 0 0 phi21
port 24 nsew
flabel metal3 -29 14662 40 14695 0 FreeSans 80 0 0 0 phi12
port 26 nsew
flabel metal3 -32 14735 37 14768 0 FreeSans 80 0 0 0 phi22
port 28 nsew
flabel metal3 -31 14802 38 14835 0 FreeSans 80 0 0 0 phi13
port 30 nsew
flabel metal3 -32 14871 37 14904 0 FreeSans 80 0 0 0 phi23
port 32 nsew
flabel metal3 -31 14946 38 14979 0 FreeSans 80 0 0 0 phi14
port 34 nsew
flabel metal3 -35 15013 34 15046 0 FreeSans 80 0 0 0 phi24
port 36 nsew
flabel metal3 -32 15082 37 15115 0 FreeSans 80 0 0 0 phi15
port 38 nsew
flabel metal3 -32 15152 37 15185 0 FreeSans 80 0 0 0 phi25
port 40 nsew
flabel metal3 -31 15223 38 15256 0 FreeSans 80 0 0 0 phi16
port 42 nsew
flabel metal3 -29 15291 40 15324 0 FreeSans 80 0 0 0 phi26
port 44 nsew
flabel metal3 -31 15362 38 15395 0 FreeSans 80 0 0 0 phi17
port 46 nsew
flabel metal3 -33 15435 36 15468 0 FreeSans 80 0 0 0 phi27
port 48 nsew
flabel metal1 67 14314 120 14330 0 FreeSans 80 0 0 0 smpl_n_d12_out_n
port 50 nsew
flabel metal1 65 14453 118 14469 0 FreeSans 80 0 0 0 phi2_n0
port 60 nsew
flabel metal1 62 14523 115 14539 0 FreeSans 80 0 0 0 phi1_n1
port 62 nsew
flabel metal1 63 14664 116 14680 0 FreeSans 80 0 0 0 phi1_n2
port 67 nsew
flabel metal1 58 14593 111 14609 0 FreeSans 80 0 0 0 phi2_n1
port 69 nsew
flabel metal1 61 14733 114 14749 0 FreeSans 80 0 0 0 phi2_n2
port 71 nsew
flabel metal1 58 14804 111 14820 0 FreeSans 80 0 0 0 phi1_n3
port 73 nsew
flabel metal1 58 14873 111 14889 0 FreeSans 80 0 0 0 phi2_n3
port 75 nsew
flabel metal1 55 14943 108 14959 0 FreeSans 80 0 0 0 phi1_n4
port 79 nsew
flabel metal1 58 15013 111 15029 0 FreeSans 80 0 0 0 phi2_n4
port 81 nsew
flabel metal1 59 15084 112 15100 0 FreeSans 80 0 0 0 phi1_n5
port 83 nsew
flabel metal1 59 15154 112 15170 0 FreeSans 80 0 0 0 phi2_n5
port 85 nsew
flabel metal1 61 15223 114 15239 0 FreeSans 80 0 0 0 phi1_n6
port 87 nsew
flabel metal1 63 15293 116 15309 0 FreeSans 80 0 0 0 phi2_n6
port 89 nsew
flabel metal1 65 15364 118 15380 0 FreeSans 80 0 0 0 phi1_n7
port 91 nsew
flabel metal1 64 15433 117 15449 0 FreeSans 80 0 0 0 phi2_n7
port 93 nsew
flabel metal1 68 14383 121 14400 0 FreeSans 80 0 0 0 phi1_n0
port 95 nsew
flabel metal1 66 14174 119 14190 0 FreeSans 80 0 0 0 vin
port 97 nsew
flabel metal1 68 14103 121 14119 0 FreeSans 80 0 0 0 gnd
port 99 nsew
flabel metal3 -29 14102 40 14134 0 FreeSans 80 0 0 0 sub
port 101 nsew
<< end >>
