magic
tech sky130A
timestamp 1729540174
<< pwell >>
rect 1465 4030 1500 4190
rect 1465 3180 1500 3340
rect 1465 2320 1500 2480
rect 1465 1465 1500 1625
rect 1465 605 1500 765
rect 1465 -240 1500 -80
<< metal1 >>
rect 1180 -960 1195 5875
rect 1210 -960 1225 5875
rect 1265 -960 1280 5875
rect 1295 -960 1310 5875
rect 1350 -960 1365 5875
rect 1380 -960 1395 5875
rect 1435 -960 1450 5875
rect 1465 5755 1500 5875
rect 2005 5755 2040 5875
rect 1465 4890 1500 5050
rect 2005 4870 2040 5030
rect 1465 4030 1500 4190
rect 2005 4030 2040 4190
rect 1465 3180 1500 3340
rect 2005 3180 2040 3340
rect 1465 2320 1500 2480
rect 2005 2325 2040 2485
rect 1465 1465 1500 1625
rect 2005 1465 2040 1625
rect 1465 605 1500 765
rect 2005 620 2040 780
rect 1465 -240 1500 -80
rect 2005 -235 2040 -75
rect 2055 -960 2070 5875
rect 2100 -960 2115 5875
rect 2130 -960 2145 5875
rect 2185 -960 2200 5875
rect 2215 -960 2230 5875
rect 2270 -960 2285 5875
rect 2300 -960 2315 5875
rect 2355 -960 2370 5875
rect 2385 -960 2400 5875
<< metal4 >>
rect 295 5710 325 5875
rect 295 4860 325 5070
rect 295 4005 325 4215
rect 295 3145 325 3360
rect 295 2295 325 2510
rect 295 1435 325 1650
rect 295 585 325 800
rect 295 -270 325 -55
use cap_model3  cap_model3_1 ~/dac_lay
timestamp 1729540174
transform 0 1 1940 1 0 3975
box 190 -1685 930 460
use cap_model3  cap_model3_2
timestamp 1729540174
transform 0 1 1940 1 0 3120
box 190 -1685 930 460
use cap_model3  cap_model3_3
timestamp 1729540174
transform 0 1 1940 1 0 2265
box 190 -1685 930 460
use cap_model3  cap_model3_4
timestamp 1729540174
transform 0 1 1940 1 0 1410
box 190 -1685 930 460
use cap_model3  cap_model3_5
timestamp 1729540174
transform 0 1 1940 1 0 555
box 190 -1685 930 460
use cap_model3  cap_model3_6
timestamp 1729540174
transform 0 1 1940 1 0 -300
box 190 -1685 930 460
use cap_model3  cap_model3_7
timestamp 1729540174
transform 0 1 1940 1 0 -1155
box 190 -1685 930 460
use cap_model3  cap_model3_8
timestamp 1729540174
transform 0 1 1940 1 0 4830
box 190 -1685 930 460
<< end >>
