magic
tech sky130A
timestamp 1729561501
<< end >>
