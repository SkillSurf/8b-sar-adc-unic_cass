magic
tech sky130A
timestamp 1729561427
<< end >>
