** sch_path: /foss/designs/sar_8bit.sch
**.subckt sar_8bit clk rst_n avss comp_out dvdd dvss vinp vinm vcm vrefp ibsnk_1u dout7,dout6,dout5,dout4,dout3,dout2,dout1,dout0
*+ data_rdy avdd vrefm
*.opin data_rdy
*.iopin avss
*.iopin avdd
*.ipin clk
*.ipin rst_n
*.opin dout7,dout6,dout5,dout4,dout3,dout2,dout1,dout0
*.iopin dvss
*.iopin dvdd
*.ipin vinp
*.ipin vinm
*.ipin vcm
*.ipin vrefp
*.ipin ibsnk_1u
*.opin comp_out
*.ipin vrefm
x1 avdd comp_out ibsnk_1u comp_p comp_m avss latch adc_comp
XM2 dvss cap_1 dvss dvss sky130_fd_pr__nfet_01v8 L=5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM3 dvss cap_2 dvss dvss sky130_fd_pr__nfet_01v8 L=5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
x3 phi1x7 phi1x6 phi1x5 phi1x4 phi1x3 phi1x2 phi1x1 phi1x0 sphi1 avss vinp phi1x_n7 phi1x_n6 phi1x_n5 phi1x_n4 phi1x_n3 phi1x_n2
+ phi1x_n1 phi1x_n0 sphi1_n avss sample vrefp phi2x7 phi2x6 phi2x5 phi2x4 phi2x3 phi2x2 phi2x1 phi2x0 sphi2 avdd sample_n vcm sphi2_n
+ phi2x_n7 phi2x_n6 phi2x_n5 phi2x_n4 phi2x_n3 phi2x_n2 phi2x_n1 phi2x_n0 comp_p capdac_p
x4 vinm sphi1 phi27 phi26 phi25 phi24 phi23 phi22 phi21 phi20 avss sample phi2_n7 phi2_n6 phi2_n5 phi2_n4 phi2_n3 phi2_n2 phi2_n1
+ phi2_n0 sphi1_n sample_n avss vrefm phi17 phi16 phi15 phi14 phi13 phi12 phi11 phi10 sphi2 avdd vcm sphi2_n phi1_n7 phi1_n6 phi1_n5
+ phi1_n4 phi1_n3 phi1_n2 phi1_n1 phi1_n0 comp_m capdac_m
x2 dvdd clk rst_n dvss comp_out cap_1 cap_2 data_rdy sample sample_n phi17 phi16 phi15 phi14 phi13 phi12 phi11 phi10 phi27 phi26
+ phi25 phi24 phi23 phi22 phi21 phi20 phi1_n7 phi1_n6 phi1_n5 phi1_n4 phi1_n3 phi1_n2 phi1_n1 phi1_n0 phi2_n7 phi2_n6 phi2_n5 phi2_n4
+ phi2_n3 phi2_n2 phi2_n1 phi2_n0 phi1x_n7 phi1x_n6 phi1x_n5 phi1x_n4 phi1x_n3 phi1x_n2 phi1x_n1 phi1x_n0 phi2x_n7 phi2x_n6 phi2x_n5
+ phi2x_n4 phi2x_n3 phi2x_n2 phi2x_n1 phi2x_n0 phi1x7 phi1x6 phi1x5 phi1x4 phi1x3 phi1x2 phi1x1 phi1x0 phi2x7 phi2x6 phi2x5 phi2x4 phi2x3
+ phi2x2 phi2x1 phi2x0 dout7 dout6 dout5 dout4 dout3 dout2 dout1 dout0 sphi1 sphi1_n sphi2_n sphi2 latch sar_digital
**.ends

* expanding   symbol:  adc_comp.sym # of pins=7
** sym_path: /foss/designs/adc_comp.sym
** sch_path: /foss/designs/adc_comp.sch
.subckt adc_comp vdd vo ibn_1u vp vm vss latch
*.iopin vss
*.iopin vdd
*.ipin vp
*.ipin vm
*.ipin latch
*.ipin ibn_1u
*.opin vo
XM3 vom1 vp vx vss sky130_fd_pr__nfet_01v8_lvt L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8
XM4 vop1 vm vx vss sky130_fd_pr__nfet_01v8_lvt L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8
XM2 vop1 vbp vdd vdd sky130_fd_pr__pfet_01v8_lvt L=5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
XM1 vom1 vbp vdd vdd sky130_fd_pr__pfet_01v8_lvt L=5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
XM6 ibn_1u ibn_1u vss vss sky130_fd_pr__nfet_01v8 L=20 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM5 vx ibn_1u vss vss sky130_fd_pr__nfet_01v8 L=20 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=12 m=12
XM7 vbp ibn_1u vss vss sky130_fd_pr__nfet_01v8 L=20 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 vbp vbp vdd vdd sky130_fd_pr__pfet_01v8_lvt L=5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 vx vop1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM10 vx vom1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM11 vop2 vom2 vss vss sky130_fd_pr__nfet_01v8 L=2 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 vom2 vop2 vss vss sky130_fd_pr__nfet_01v8 L=2 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 net5 vom1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 net4 vop1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 vom2 latch_n vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18 vop2 latch_n vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM19 net1 vop2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM20 net1 vop2 vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM21 net2 net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM22 net2 net1 vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM23 net3 vom2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM24 net3 vom2 vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 net6 vop2 net4 vdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16 net7 vom2 net5 vdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM25 net6 latch vom2 vss sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM26 net7 latch vop2 vss sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x30 latch vss vss vdd vdd latch_n sky130_fd_sc_hd__inv_1
XM27 vss ibn_1u vss vss sky130_fd_pr__nfet_01v8 L=20 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM28 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM29 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=20 m=20
XM30 vdd vbp vdd vdd sky130_fd_pr__pfet_01v8_lvt L=5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
XM31 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
x7 net2 vss vss vdd vdd vo sky130_fd_sc_hd__inv_4
.ends


* expanding   symbol:  capdac_p.sym # of pins=17
** sym_path: /foss/designs/capdac_p.sym
** sch_path: /foss/designs/capdac_p.sch
.subckt capdac_p phi17 phi16 phi15 phi14 phi13 phi12 phi11 phi10 sphi1 sub vin phi1_n7 phi1_n6 phi1_n5 phi1_n4 phi1_n3 phi1_n2
+ phi1_n1 phi1_n0 sphi1_n GND sample vref phi27 phi26 phi25 phi24 phi23 phi22 phi21 phi20 sphi2 vdd sample_n vcm sphi2_n phi2_n7 phi2_n6
+ phi2_n5 phi2_n4 phi2_n3 phi2_n2 phi2_n1 phi2_n0 com_x
*.ipin phi17,phi16,phi15,phi14,phi13,phi12,phi11,phi10
*.ipin phi1_n7,phi1_n6,phi1_n5,phi1_n4,phi1_n3,phi1_n2,phi1_n1,phi1_n0
*.iopin vdd
*.iopin GND
*.iopin sub
*.ipin phi27,phi26,phi25,phi24,phi23,phi22,phi21,phi20
*.ipin phi2_n7,phi2_n6,phi2_n5,phi2_n4,phi2_n3,phi2_n2,phi2_n1,phi2_n0
*.opin com_x
*.ipin sphi1
*.ipin sphi1_n
*.ipin sphi2
*.ipin sphi2_n
*.ipin vcm
*.ipin vref
*.ipin vin
*.ipin sample_n
*.ipin sample
x2 net1 sub GND vdd sphi1 sphi2 sphi2_n sphi1_n com_x cap_switch_block
x1 net1 sub GND vdd phi10 phi20 phi2_n0 phi1_n0 com_x cap_switch_block
x12 net1 sub GND vdd phi11 phi21 phi2_n1 phi1_n1 com_x cap_switch_block
x11 net1 sub GND vdd phi11 phi21 phi2_n1 phi1_n1 com_x cap_switch_block
x54 net1 sub GND vdd phi12 phi22 phi2_n2 phi1_n2 com_x cap_switch_block
x53 net1 sub GND vdd phi12 phi22 phi2_n2 phi1_n2 com_x cap_switch_block
x52 net1 sub GND vdd phi12 phi22 phi2_n2 phi1_n2 com_x cap_switch_block
x51 net1 sub GND vdd phi12 phi22 phi2_n2 phi1_n2 com_x cap_switch_block
x68 net1 sub GND vdd phi13 phi23 phi2_n3 phi1_n3 com_x cap_switch_block
x67 net1 sub GND vdd phi13 phi23 phi2_n3 phi1_n3 com_x cap_switch_block
x66 net1 sub GND vdd phi13 phi23 phi2_n3 phi1_n3 com_x cap_switch_block
x65 net1 sub GND vdd phi13 phi23 phi2_n3 phi1_n3 com_x cap_switch_block
x64 net1 sub GND vdd phi13 phi23 phi2_n3 phi1_n3 com_x cap_switch_block
x63 net1 sub GND vdd phi13 phi23 phi2_n3 phi1_n3 com_x cap_switch_block
x62 net1 sub GND vdd phi13 phi23 phi2_n3 phi1_n3 com_x cap_switch_block
x61 net1 sub GND vdd phi13 phi23 phi2_n3 phi1_n3 com_x cap_switch_block
x716 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x715 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x714 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x713 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x712 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x711 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x710 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x79 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x78 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x77 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x76 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x75 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x74 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x73 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x72 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x71 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x832 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x831 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x830 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x829 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x828 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x827 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x826 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x825 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x824 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x823 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x822 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x821 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x820 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x819 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x818 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x817 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x816 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x815 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x814 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x813 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x812 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x811 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x810 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x89 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x88 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x87 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x86 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x85 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x84 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x83 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x82 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x81 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x964 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x963 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x962 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x961 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x960 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x959 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x958 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x957 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x956 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x955 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x954 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x953 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x952 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x951 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x950 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x949 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x948 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x947 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x946 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x945 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x944 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x943 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x942 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x941 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x940 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x939 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x938 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x937 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x936 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x935 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x934 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x933 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x932 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x931 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x930 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x929 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x928 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x927 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x926 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x925 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x924 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x923 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x922 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x921 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x920 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x919 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x918 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x917 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x916 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x915 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x914 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x913 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x912 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x911 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x910 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x99 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x98 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x97 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x96 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x95 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x94 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x93 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x92 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x91 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x10128 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10127 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10126 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10125 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10124 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10123 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10122 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10121 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10120 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10119 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10118 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10117 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10116 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10115 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10114 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10113 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10112 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10111 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10110 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10109 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10108 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10107 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10106 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10105 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10104 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10103 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10102 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10101 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10100 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1099 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1098 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1097 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1096 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1095 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1094 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1093 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1092 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1091 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1090 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1089 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1088 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1087 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1086 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1085 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1084 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1083 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1082 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1081 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1080 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1079 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1078 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1077 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1076 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1075 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1074 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1073 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1072 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1071 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1070 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1069 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1068 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1067 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1066 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1065 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1064 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1063 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1062 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1061 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1060 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1059 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1058 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1057 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1056 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1055 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1054 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1053 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1052 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1051 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1050 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1049 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1048 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1047 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1046 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1045 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1044 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1043 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1042 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1041 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1040 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1039 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1038 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1037 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1036 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1035 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1034 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1033 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1032 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1031 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1030 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1029 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1028 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1027 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1026 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1025 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1024 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1023 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1022 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1021 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1020 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1019 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1018 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1017 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1016 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1015 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1014 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1013 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1012 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1011 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1010 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x109 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x108 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x107 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x106 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x105 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x104 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x103 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x102 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x101 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x5[10] sphi2 sub net1 vref vdd sphi2_n tg_final
x5[9] sphi2 sub net1 vref vdd sphi2_n tg_final
x5[8] sphi2 sub net1 vref vdd sphi2_n tg_final
x5[7] sphi2 sub net1 vref vdd sphi2_n tg_final
x5[6] sphi2 sub net1 vref vdd sphi2_n tg_final
x5[5] sphi2 sub net1 vref vdd sphi2_n tg_final
x5[4] sphi2 sub net1 vref vdd sphi2_n tg_final
x5[3] sphi2 sub net1 vref vdd sphi2_n tg_final
x5[2] sphi2 sub net1 vref vdd sphi2_n tg_final
x5[1] sphi2 sub net1 vref vdd sphi2_n tg_final
x6[10] sphi1 sub net1 vin vdd sphi1_n tg_final
x6[9] sphi1 sub net1 vin vdd sphi1_n tg_final
x6[8] sphi1 sub net1 vin vdd sphi1_n tg_final
x6[7] sphi1 sub net1 vin vdd sphi1_n tg_final
x6[6] sphi1 sub net1 vin vdd sphi1_n tg_final
x6[5] sphi1 sub net1 vin vdd sphi1_n tg_final
x6[4] sphi1 sub net1 vin vdd sphi1_n tg_final
x6[3] sphi1 sub net1 vin vdd sphi1_n tg_final
x6[2] sphi1 sub net1 vin vdd sphi1_n tg_final
x6[1] sphi1 sub net1 vin vdd sphi1_n tg_final
x3[10] sample sub com_x vcm vdd sample_n tg_final
x3[9] sample sub com_x vcm vdd sample_n tg_final
x3[8] sample sub com_x vcm vdd sample_n tg_final
x3[7] sample sub com_x vcm vdd sample_n tg_final
x3[6] sample sub com_x vcm vdd sample_n tg_final
x3[5] sample sub com_x vcm vdd sample_n tg_final
x3[4] sample sub com_x vcm vdd sample_n tg_final
x3[3] sample sub com_x vcm vdd sample_n tg_final
x3[2] sample sub com_x vcm vdd sample_n tg_final
x3[1] sample sub com_x vcm vdd sample_n tg_final
x268 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x267 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x266 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x265 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x264 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x263 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x262 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x261 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x260 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x259 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x258 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x257 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x256 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x255 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x254 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x253 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x252 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x251 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x250 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x249 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x248 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x247 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x246 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x245 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x244 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x243 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x242 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x241 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x240 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x239 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x238 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x237 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x236 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x235 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x234 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x233 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x232 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x231 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x230 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x229 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x228 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x227 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x226 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x225 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x224 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x223 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x222 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x221 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x220 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x219 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x218 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x217 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x216 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x215 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x214 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x213 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x212 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x211 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x210 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x29 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x28 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x27 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x26 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x25 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x24 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x23 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x22 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x21 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
.ends


* expanding   symbol:  capdac_m.sym # of pins=17
** sym_path: /foss/designs/capdac_m.sym
** sch_path: /foss/designs/capdac_m.sch
.subckt capdac_m vin sphi1 phi17 phi16 phi15 phi14 phi13 phi12 phi11 phi10 sub sample phi1_n7 phi1_n6 phi1_n5 phi1_n4 phi1_n3
+ phi1_n2 phi1_n1 phi1_n0 sphi1_n sample_n GND vref phi27 phi26 phi25 phi24 phi23 phi22 phi21 phi20 sphi2 vdd vcm sphi2_n phi2_n7 phi2_n6
+ phi2_n5 phi2_n4 phi2_n3 phi2_n2 phi2_n1 phi2_n0 com_x
*.ipin phi17,phi16,phi15,phi14,phi13,phi12,phi11,phi10
*.ipin phi1_n7,phi1_n6,phi1_n5,phi1_n4,phi1_n3,phi1_n2,phi1_n1,phi1_n0
*.iopin vdd
*.iopin GND
*.iopin sub
*.ipin phi27,phi26,phi25,phi24,phi23,phi22,phi21,phi20
*.ipin phi2_n7,phi2_n6,phi2_n5,phi2_n4,phi2_n3,phi2_n2,phi2_n1,phi2_n0
*.opin com_x
*.ipin sphi1
*.ipin sphi1_n
*.ipin sphi2
*.ipin sphi2_n
*.ipin vcm
*.ipin vref
*.ipin sample
*.ipin sample_n
*.ipin vin
x2 net1 sub net1 vdd sphi1 sphi2 sphi2_n sphi1_n com_x cap_switch_block
x1 net1 sub GND vdd phi10 phi20 phi2_n0 phi1_n0 com_x cap_switch_block
x12 net1 sub GND vdd phi11 phi21 phi2_n1 phi1_n1 com_x cap_switch_block
x11 net1 sub GND vdd phi11 phi21 phi2_n1 phi1_n1 com_x cap_switch_block
x54 net1 sub GND vdd phi12 phi22 phi2_n2 phi1_n2 com_x cap_switch_block
x53 net1 sub GND vdd phi12 phi22 phi2_n2 phi1_n2 com_x cap_switch_block
x52 net1 sub GND vdd phi12 phi22 phi2_n2 phi1_n2 com_x cap_switch_block
x51 net1 sub GND vdd phi12 phi22 phi2_n2 phi1_n2 com_x cap_switch_block
x68 net1 sub GND vdd phi13 phi23 phi2_n3 phi1_n3 com_x cap_switch_block
x67 net1 sub GND vdd phi13 phi23 phi2_n3 phi1_n3 com_x cap_switch_block
x66 net1 sub GND vdd phi13 phi23 phi2_n3 phi1_n3 com_x cap_switch_block
x65 net1 sub GND vdd phi13 phi23 phi2_n3 phi1_n3 com_x cap_switch_block
x64 net1 sub GND vdd phi13 phi23 phi2_n3 phi1_n3 com_x cap_switch_block
x63 net1 sub GND vdd phi13 phi23 phi2_n3 phi1_n3 com_x cap_switch_block
x62 net1 sub GND vdd phi13 phi23 phi2_n3 phi1_n3 com_x cap_switch_block
x61 net1 sub GND vdd phi13 phi23 phi2_n3 phi1_n3 com_x cap_switch_block
x716 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x715 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x714 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x713 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x712 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x711 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x710 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x79 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x78 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x77 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x76 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x75 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x74 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x73 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x72 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x71 net1 sub GND vdd phi14 phi24 phi2_n4 phi1_n4 com_x cap_switch_block
x832 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x831 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x830 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x829 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x828 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x827 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x826 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x825 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x824 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x823 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x822 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x821 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x820 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x819 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x818 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x817 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x816 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x815 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x814 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x813 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x812 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x811 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x810 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x89 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x88 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x87 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x86 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x85 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x84 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x83 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x82 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x81 net1 sub GND vdd phi15 phi25 phi2_n5 phi1_n5 com_x cap_switch_block
x964 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x963 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x962 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x961 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x960 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x959 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x958 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x957 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x956 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x955 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x954 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x953 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x952 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x951 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x950 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x949 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x948 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x947 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x946 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x945 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x944 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x943 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x942 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x941 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x940 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x939 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x938 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x937 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x936 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x935 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x934 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x933 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x932 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x931 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x930 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x929 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x928 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x927 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x926 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x925 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x924 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x923 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x922 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x921 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x920 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x919 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x918 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x917 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x916 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x915 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x914 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x913 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x912 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x911 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x910 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x99 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x98 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x97 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x96 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x95 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x94 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x93 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x92 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x91 net1 sub GND vdd phi16 phi26 phi2_n6 phi1_n6 com_x cap_switch_block
x10128 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10127 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10126 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10125 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10124 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10123 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10122 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10121 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10120 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10119 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10118 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10117 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10116 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10115 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10114 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10113 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10112 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10111 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10110 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10109 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10108 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10107 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10106 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10105 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10104 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10103 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10102 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10101 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x10100 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1099 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1098 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1097 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1096 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1095 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1094 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1093 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1092 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1091 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1090 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1089 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1088 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1087 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1086 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1085 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1084 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1083 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1082 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1081 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1080 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1079 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1078 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1077 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1076 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1075 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1074 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1073 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1072 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1071 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1070 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1069 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1068 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1067 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1066 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1065 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1064 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1063 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1062 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1061 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1060 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1059 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1058 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1057 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1056 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1055 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1054 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1053 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1052 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1051 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1050 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1049 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1048 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1047 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1046 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1045 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1044 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1043 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1042 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1041 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1040 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1039 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1038 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1037 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1036 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1035 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1034 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1033 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1032 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1031 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1030 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1029 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1028 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1027 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1026 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1025 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1024 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1023 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1022 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1021 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1020 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1019 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1018 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1017 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1016 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1015 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1014 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1013 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1012 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1011 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x1010 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x109 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x108 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x107 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x106 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x105 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x104 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x103 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x102 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x101 net1 sub GND vdd phi17 phi27 phi2_n7 phi1_n7 com_x cap_switch_block
x410 sphi2 sub net1 vref vdd sphi2_n tg_final
x49 sphi2 sub net1 vref vdd sphi2_n tg_final
x48 sphi2 sub net1 vref vdd sphi2_n tg_final
x47 sphi2 sub net1 vref vdd sphi2_n tg_final
x46 sphi2 sub net1 vref vdd sphi2_n tg_final
x45 sphi2 sub net1 vref vdd sphi2_n tg_final
x44 sphi2 sub net1 vref vdd sphi2_n tg_final
x43 sphi2 sub net1 vref vdd sphi2_n tg_final
x42 sphi2 sub net1 vref vdd sphi2_n tg_final
x41 sphi2 sub net1 vref vdd sphi2_n tg_final
x210 sphi1 sub net1 vin vdd sphi1_n tg_final
x29 sphi1 sub net1 vin vdd sphi1_n tg_final
x28 sphi1 sub net1 vin vdd sphi1_n tg_final
x27 sphi1 sub net1 vin vdd sphi1_n tg_final
x26 sphi1 sub net1 vin vdd sphi1_n tg_final
x25 sphi1 sub net1 vin vdd sphi1_n tg_final
x24 sphi1 sub net1 vin vdd sphi1_n tg_final
x23 sphi1 sub net1 vin vdd sphi1_n tg_final
x22 sphi1 sub net1 vin vdd sphi1_n tg_final
x21 sphi1 sub net1 vin vdd sphi1_n tg_final
x310 sample sub com_x vcm vdd sample_n tg_final
x39 sample sub com_x vcm vdd sample_n tg_final
x38 sample sub com_x vcm vdd sample_n tg_final
x37 sample sub com_x vcm vdd sample_n tg_final
x36 sample sub com_x vcm vdd sample_n tg_final
x35 sample sub com_x vcm vdd sample_n tg_final
x34 sample sub com_x vcm vdd sample_n tg_final
x33 sample sub com_x vcm vdd sample_n tg_final
x32 sample sub com_x vcm vdd sample_n tg_final
x31 sample sub com_x vcm vdd sample_n tg_final
x1168 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1167 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1166 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1165 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1164 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1163 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1162 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1161 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1160 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1159 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1158 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1157 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1156 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1155 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1154 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1153 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1152 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1151 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1150 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1149 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1148 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1147 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1146 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1145 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1144 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1143 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1142 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1141 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1140 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1139 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1138 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1137 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1136 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1135 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1134 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1133 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1132 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1131 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1130 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1129 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1128 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1127 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1126 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1125 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1124 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1123 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1122 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1121 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1120 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1119 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1118 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1117 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1116 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1115 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1114 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1113 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1112 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1111 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x1110 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x119 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x118 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x117 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x116 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x115 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x114 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x113 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x112 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
x111 GND sub GND vdd vdd vdd GND GND GND cap_switch_block
.ends


* expanding   symbol:  sar_digital.sym # of pins=24
** sym_path: /foss/designs/sar_digital.sym
** sch_path: /foss/designs/sar_digital.sch
.subckt sar_digital vdd clk rst_n vss comp_out cap_1 cap_2 data_rdy sample sample_n phi17 phi16 phi15 phi14 phi13 phi12 phi11
+ phi10 phi27 phi26 phi25 phi24 phi23 phi22 phi21 phi20 phi1_n7 phi1_n6 phi1_n5 phi1_n4 phi1_n3 phi1_n2 phi1_n1 phi1_n0 phi2_n7 phi2_n6
+ phi2_n5 phi2_n4 phi2_n3 phi2_n2 phi2_n1 phi2_n0 phi1x_n7 phi1x_n6 phi1x_n5 phi1x_n4 phi1x_n3 phi1x_n2 phi1x_n1 phi1x_n0 phi2x_n7 phi2x_n6
+ phi2x_n5 phi2x_n4 phi2x_n3 phi2x_n2 phi2x_n1 phi2x_n0 phi1x7 phi1x6 phi1x5 phi1x4 phi1x3 phi1x2 phi1x1 phi1x0 phi2x7 phi2x6 phi2x5 phi2x4
+ phi2x3 phi2x2 phi2x1 phi2x0 dout7 dout6 dout5 dout4 dout3 dout2 dout1 dout0 sphi1 sphi1_n sphi2_n sphi2 latch
*.opin data_rdy
*.iopin vss
*.iopin vdd
*.ipin clk
*.ipin rst_n
*.ipin comp_out
*.opin sample
*.opin sample_n
*.iopin cap_1
*.iopin cap_2
*.opin phi17,phi16,phi15,phi14,phi13,phi12,phi11,phi10
*.opin phi1_n7,phi1_n6,phi1_n5,phi1_n4,phi1_n3,phi1_n2,phi1_n1,phi1_n0
*.opin phi1x_n7,phi1x_n6,phi1x_n5,phi1x_n4,phi1x_n3,phi1x_n2,phi1x_n1,phi1x_n0
*.opin phi1x7,phi1x6,phi1x5,phi1x4,phi1x3,phi1x2,phi1x1,phi1x0
*.opin sphi1
*.opin sphi1_n
*.opin sphi2_n
*.opin sphi2
*.opin phi27,phi26,phi25,phi24,phi23,phi22,phi21,phi20
*.opin phi2_n7,phi2_n6,phi2_n5,phi2_n4,phi2_n3,phi2_n2,phi2_n1,phi2_n0
*.opin phi2x_n7,phi2x_n6,phi2x_n5,phi2x_n4,phi2x_n3,phi2x_n2,phi2x_n1,phi2x_n0
*.opin phi2x7,phi2x6,phi2x5,phi2x4,phi2x3,phi2x2,phi2x1,phi2x0
*.opin latch
*.opin dout7,dout6,dout5,dout4,dout3,dout2,dout1,dout0
x2 clk data_rdy sample rst_n sample_n comp_out vss vdd data7 data6 data5 data4 data3 data2 data1 data0 data_n7 data_n6 data_n5
+ data_n4 data_n3 data_n2 data_n1 data_n0 sar_controller
x2[7] data7 vss vss vdd vdd net1[7] sky130_fd_sc_hd__inv_2
x2[6] data6 vss vss vdd vdd net1[6] sky130_fd_sc_hd__inv_2
x2[5] data5 vss vss vdd vdd net1[5] sky130_fd_sc_hd__inv_2
x2[4] data4 vss vss vdd vdd net1[4] sky130_fd_sc_hd__inv_2
x2[3] data3 vss vss vdd vdd net1[3] sky130_fd_sc_hd__inv_2
x2[2] data2 vss vss vdd vdd net1[2] sky130_fd_sc_hd__inv_2
x2[1] data1 vss vss vdd vdd net1[1] sky130_fd_sc_hd__inv_2
x2[0] data0 vss vss vdd vdd net1[0] sky130_fd_sc_hd__inv_2
x6[7] data7 d7 vss vss vdd vdd net2[7] sky130_fd_sc_hd__nor2_1
x6[6] data6 d6 vss vss vdd vdd net2[6] sky130_fd_sc_hd__nor2_1
x6[5] data5 d5 vss vss vdd vdd net2[5] sky130_fd_sc_hd__nor2_1
x6[4] data4 d4 vss vss vdd vdd net2[4] sky130_fd_sc_hd__nor2_1
x6[3] data3 d3 vss vss vdd vdd net2[3] sky130_fd_sc_hd__nor2_1
x6[2] data2 d2 vss vss vdd vdd net2[2] sky130_fd_sc_hd__nor2_1
x6[1] data1 d1 vss vss vdd vdd net2[1] sky130_fd_sc_hd__nor2_1
x6[0] data0 d0 vss vss vdd vdd net2[0] sky130_fd_sc_hd__nor2_1
x16[7] dn7 net1[7] vss vss vdd vdd net5[7] sky130_fd_sc_hd__nor2_1
x16[6] dn6 net1[6] vss vss vdd vdd net5[6] sky130_fd_sc_hd__nor2_1
x16[5] dn5 net1[5] vss vss vdd vdd net5[5] sky130_fd_sc_hd__nor2_1
x16[4] dn4 net1[4] vss vss vdd vdd net5[4] sky130_fd_sc_hd__nor2_1
x16[3] dn3 net1[3] vss vss vdd vdd net5[3] sky130_fd_sc_hd__nor2_1
x16[2] dn2 net1[2] vss vss vdd vdd net5[2] sky130_fd_sc_hd__nor2_1
x16[1] dn1 net1[1] vss vss vdd vdd net5[1] sky130_fd_sc_hd__nor2_1
x16[0] dn0 net1[0] vss vss vdd vdd net5[0] sky130_fd_sc_hd__nor2_1
x17[7] net2[7] vss vss vdd vdd net3[7] sky130_fd_sc_hd__buf_1
x17[6] net2[6] vss vss vdd vdd net3[6] sky130_fd_sc_hd__buf_1
x17[5] net2[5] vss vss vdd vdd net3[5] sky130_fd_sc_hd__buf_1
x17[4] net2[4] vss vss vdd vdd net3[4] sky130_fd_sc_hd__buf_1
x17[3] net2[3] vss vss vdd vdd net3[3] sky130_fd_sc_hd__buf_1
x17[2] net2[2] vss vss vdd vdd net3[2] sky130_fd_sc_hd__buf_1
x17[1] net2[1] vss vss vdd vdd net3[1] sky130_fd_sc_hd__buf_1
x17[0] net2[0] vss vss vdd vdd net3[0] sky130_fd_sc_hd__buf_1
x35[7] net3[7] vss vss vdd vdd net4[7] sky130_fd_sc_hd__buf_2
x35[6] net3[6] vss vss vdd vdd net4[6] sky130_fd_sc_hd__buf_2
x35[5] net3[5] vss vss vdd vdd net4[5] sky130_fd_sc_hd__buf_2
x35[4] net3[4] vss vss vdd vdd net4[4] sky130_fd_sc_hd__buf_2
x35[3] net3[3] vss vss vdd vdd net4[3] sky130_fd_sc_hd__buf_2
x35[2] net3[2] vss vss vdd vdd net4[2] sky130_fd_sc_hd__buf_2
x35[1] net3[1] vss vss vdd vdd net4[1] sky130_fd_sc_hd__buf_2
x35[0] net3[0] vss vss vdd vdd net4[0] sky130_fd_sc_hd__buf_2
x36[7] net4[7] vss vss vdd vdd dn7 sky130_fd_sc_hd__buf_1
x36[6] net4[6] vss vss vdd vdd dn6 sky130_fd_sc_hd__buf_1
x36[5] net4[5] vss vss vdd vdd dn5 sky130_fd_sc_hd__buf_1
x36[4] net4[4] vss vss vdd vdd dn4 sky130_fd_sc_hd__buf_1
x36[3] net4[3] vss vss vdd vdd dn3 sky130_fd_sc_hd__buf_1
x36[2] net4[2] vss vss vdd vdd dn2 sky130_fd_sc_hd__buf_1
x36[1] net4[1] vss vss vdd vdd dn1 sky130_fd_sc_hd__buf_1
x36[0] net4[0] vss vss vdd vdd dn0 sky130_fd_sc_hd__buf_1
x37[7] net5[7] vss vss vdd vdd net6[7] sky130_fd_sc_hd__buf_1
x37[6] net5[6] vss vss vdd vdd net6[6] sky130_fd_sc_hd__buf_1
x37[5] net5[5] vss vss vdd vdd net6[5] sky130_fd_sc_hd__buf_1
x37[4] net5[4] vss vss vdd vdd net6[4] sky130_fd_sc_hd__buf_1
x37[3] net5[3] vss vss vdd vdd net6[3] sky130_fd_sc_hd__buf_1
x37[2] net5[2] vss vss vdd vdd net6[2] sky130_fd_sc_hd__buf_1
x37[1] net5[1] vss vss vdd vdd net6[1] sky130_fd_sc_hd__buf_1
x37[0] net5[0] vss vss vdd vdd net6[0] sky130_fd_sc_hd__buf_1
x38[7] net6[7] vss vss vdd vdd net7[7] sky130_fd_sc_hd__buf_2
x38[6] net6[6] vss vss vdd vdd net7[6] sky130_fd_sc_hd__buf_2
x38[5] net6[5] vss vss vdd vdd net7[5] sky130_fd_sc_hd__buf_2
x38[4] net6[4] vss vss vdd vdd net7[4] sky130_fd_sc_hd__buf_2
x38[3] net6[3] vss vss vdd vdd net7[3] sky130_fd_sc_hd__buf_2
x38[2] net6[2] vss vss vdd vdd net7[2] sky130_fd_sc_hd__buf_2
x38[1] net6[1] vss vss vdd vdd net7[1] sky130_fd_sc_hd__buf_2
x38[0] net6[0] vss vss vdd vdd net7[0] sky130_fd_sc_hd__buf_2
x39[7] net7[7] vss vss vdd vdd d7 sky130_fd_sc_hd__buf_1
x39[6] net7[6] vss vss vdd vdd d6 sky130_fd_sc_hd__buf_1
x39[5] net7[5] vss vss vdd vdd d5 sky130_fd_sc_hd__buf_1
x39[4] net7[4] vss vss vdd vdd d4 sky130_fd_sc_hd__buf_1
x39[3] net7[3] vss vss vdd vdd d3 sky130_fd_sc_hd__buf_1
x39[2] net7[2] vss vss vdd vdd d2 sky130_fd_sc_hd__buf_1
x39[1] net7[1] vss vss vdd vdd d1 sky130_fd_sc_hd__buf_1
x39[0] net7[0] vss vss vdd vdd d0 sky130_fd_sc_hd__buf_1
x5[7] d7 sphi1 vss vss vdd vdd net8 sky130_fd_sc_hd__or2_2
x1[6] sample_n dn6 vss vss vdd vdd net30[6] sky130_fd_sc_hd__and2_2
x1[5] sample_n dn5 vss vss vdd vdd net30[5] sky130_fd_sc_hd__and2_2
x1[4] sample_n dn4 vss vss vdd vdd net30[4] sky130_fd_sc_hd__and2_2
x1[3] sample_n dn3 vss vss vdd vdd net30[3] sky130_fd_sc_hd__and2_2
x1[2] sample_n dn2 vss vss vdd vdd net30[2] sky130_fd_sc_hd__and2_2
x1[1] sample_n dn1 vss vss vdd vdd net30[1] sky130_fd_sc_hd__and2_2
x1[0] sample_n dn0 vss vss vdd vdd net30[0] sky130_fd_sc_hd__and2_2
x42 clk vss vss vdd vdd cap_1 sky130_fd_sc_hd__buf_1
x43 cap_1 vss vss vdd vdd cap_2 sky130_fd_sc_hd__buf_1
x44 net9 vss vss vdd vdd latch sky130_fd_sc_hd__inv_2
x45 cap_2 vss vss vdd vdd net9 sky130_fd_sc_hd__buf_1
x46 sample vss vss vdd vdd net10 sky130_fd_sc_hd__inv_2
x47 sample net12 vss vss vdd vdd net13 sky130_fd_sc_hd__nor2_1
x48 net11 net10 vss vss vdd vdd net17 sky130_fd_sc_hd__nor2_1
x49 net13 vss vss vdd vdd net14 sky130_fd_sc_hd__buf_1
x50 net14 vss vss vdd vdd net15 sky130_fd_sc_hd__buf_6
x51 net15 vss vss vdd vdd net16 sky130_fd_sc_hd__buf_1
x52 net17 vss vss vdd vdd net18 sky130_fd_sc_hd__buf_1
x53 net18 vss vss vdd vdd net19 sky130_fd_sc_hd__buf_6
x54 net19 vss vss vdd vdd net20 sky130_fd_sc_hd__buf_1
x55 net16 vss vss vdd vdd net24 sky130_fd_sc_hd__buf_6
x56 net20 vss vss vdd vdd net22 sky130_fd_sc_hd__buf_6
x41[6] d6 sample vss vss vdd vdd net21[6] sky130_fd_sc_hd__or2_2
x41[5] d5 sample vss vss vdd vdd net21[5] sky130_fd_sc_hd__or2_2
x41[4] d4 sample vss vss vdd vdd net21[4] sky130_fd_sc_hd__or2_2
x41[3] d3 sample vss vss vdd vdd net21[3] sky130_fd_sc_hd__or2_2
x41[2] d2 sample vss vss vdd vdd net21[2] sky130_fd_sc_hd__or2_2
x41[1] d1 sample vss vss vdd vdd net21[1] sky130_fd_sc_hd__or2_2
x41[0] d0 sample vss vss vdd vdd net21[0] sky130_fd_sc_hd__or2_2
x57 sphi2 dn7 vss vss vdd vdd net31 sky130_fd_sc_hd__and2_2
x58 net22 vss vss vdd vdd net23 sky130_fd_sc_hd__buf_1
x59 net23 vss vss vdd vdd net26 sky130_fd_sc_hd__buf_6
x60 net24 vss vss vdd vdd net25 sky130_fd_sc_hd__buf_1
x61 net25 vss vss vdd vdd net28 sky130_fd_sc_hd__buf_6
x62 net26 vss vss vdd vdd net27 sky130_fd_sc_hd__buf_1
x63 net27 vss vss vdd vdd net12 sky130_fd_sc_hd__buf_4
x64 net28 vss vss vdd vdd net29 sky130_fd_sc_hd__buf_1
x65 net29 vss vss vdd vdd net11 sky130_fd_sc_hd__buf_4
x43[7] d7 vss vss vdd vdd net32[7] sky130_fd_sc_hd__buf_1
x43[6] d6 vss vss vdd vdd net32[6] sky130_fd_sc_hd__buf_1
x43[5] d5 vss vss vdd vdd net32[5] sky130_fd_sc_hd__buf_1
x43[4] d4 vss vss vdd vdd net32[4] sky130_fd_sc_hd__buf_1
x43[3] d3 vss vss vdd vdd net32[3] sky130_fd_sc_hd__buf_1
x43[2] d2 vss vss vdd vdd net32[2] sky130_fd_sc_hd__buf_1
x43[1] d1 vss vss vdd vdd net32[1] sky130_fd_sc_hd__buf_1
x43[0] d0 vss vss vdd vdd net32[0] sky130_fd_sc_hd__buf_1
x44[7] net32[7] vss vss vdd vdd net33[7] sky130_fd_sc_hd__buf_2
x44[6] net32[6] vss vss vdd vdd net33[6] sky130_fd_sc_hd__buf_2
x44[5] net32[5] vss vss vdd vdd net33[5] sky130_fd_sc_hd__buf_2
x44[4] net32[4] vss vss vdd vdd net33[4] sky130_fd_sc_hd__buf_2
x44[3] net32[3] vss vss vdd vdd net33[3] sky130_fd_sc_hd__buf_2
x44[2] net32[2] vss vss vdd vdd net33[2] sky130_fd_sc_hd__buf_2
x44[1] net32[1] vss vss vdd vdd net33[1] sky130_fd_sc_hd__buf_2
x44[0] net32[0] vss vss vdd vdd net33[0] sky130_fd_sc_hd__buf_2
x45[7] net33[7] vss vss vdd vdd net34[7] sky130_fd_sc_hd__buf_4
x45[6] net33[6] vss vss vdd vdd net34[6] sky130_fd_sc_hd__buf_4
x45[5] net33[5] vss vss vdd vdd net34[5] sky130_fd_sc_hd__buf_4
x45[4] net33[4] vss vss vdd vdd net34[4] sky130_fd_sc_hd__buf_4
x45[3] net33[3] vss vss vdd vdd net34[3] sky130_fd_sc_hd__buf_4
x45[2] net33[2] vss vss vdd vdd net34[2] sky130_fd_sc_hd__buf_4
x45[1] net33[1] vss vss vdd vdd net34[1] sky130_fd_sc_hd__buf_4
x45[0] net33[0] vss vss vdd vdd net34[0] sky130_fd_sc_hd__buf_4
x46[7] net34[7] vss vss vdd vdd phi17 sky130_fd_sc_hd__buf_8
x46[6] net34[6] vss vss vdd vdd phi16 sky130_fd_sc_hd__buf_8
x46[5] net34[5] vss vss vdd vdd phi15 sky130_fd_sc_hd__buf_8
x46[4] net34[4] vss vss vdd vdd phi14 sky130_fd_sc_hd__buf_8
x46[3] net34[3] vss vss vdd vdd phi13 sky130_fd_sc_hd__buf_8
x46[2] net34[2] vss vss vdd vdd phi12 sky130_fd_sc_hd__buf_8
x46[1] net34[1] vss vss vdd vdd phi11 sky130_fd_sc_hd__buf_8
x46[0] net34[0] vss vss vdd vdd phi10 sky130_fd_sc_hd__buf_8
x47[7] dn7 vss vss vdd vdd net35[7] sky130_fd_sc_hd__buf_1
x47[6] dn6 vss vss vdd vdd net35[6] sky130_fd_sc_hd__buf_1
x47[5] dn5 vss vss vdd vdd net35[5] sky130_fd_sc_hd__buf_1
x47[4] dn4 vss vss vdd vdd net35[4] sky130_fd_sc_hd__buf_1
x47[3] dn3 vss vss vdd vdd net35[3] sky130_fd_sc_hd__buf_1
x47[2] dn2 vss vss vdd vdd net35[2] sky130_fd_sc_hd__buf_1
x47[1] dn1 vss vss vdd vdd net35[1] sky130_fd_sc_hd__buf_1
x47[0] dn0 vss vss vdd vdd net35[0] sky130_fd_sc_hd__buf_1
x48[7] net35[7] vss vss vdd vdd net36[7] sky130_fd_sc_hd__buf_2
x48[6] net35[6] vss vss vdd vdd net36[6] sky130_fd_sc_hd__buf_2
x48[5] net35[5] vss vss vdd vdd net36[5] sky130_fd_sc_hd__buf_2
x48[4] net35[4] vss vss vdd vdd net36[4] sky130_fd_sc_hd__buf_2
x48[3] net35[3] vss vss vdd vdd net36[3] sky130_fd_sc_hd__buf_2
x48[2] net35[2] vss vss vdd vdd net36[2] sky130_fd_sc_hd__buf_2
x48[1] net35[1] vss vss vdd vdd net36[1] sky130_fd_sc_hd__buf_2
x48[0] net35[0] vss vss vdd vdd net36[0] sky130_fd_sc_hd__buf_2
x49[7] net36[7] vss vss vdd vdd net37[7] sky130_fd_sc_hd__buf_4
x49[6] net36[6] vss vss vdd vdd net37[6] sky130_fd_sc_hd__buf_4
x49[5] net36[5] vss vss vdd vdd net37[5] sky130_fd_sc_hd__buf_4
x49[4] net36[4] vss vss vdd vdd net37[4] sky130_fd_sc_hd__buf_4
x49[3] net36[3] vss vss vdd vdd net37[3] sky130_fd_sc_hd__buf_4
x49[2] net36[2] vss vss vdd vdd net37[2] sky130_fd_sc_hd__buf_4
x49[1] net36[1] vss vss vdd vdd net37[1] sky130_fd_sc_hd__buf_4
x49[0] net36[0] vss vss vdd vdd net37[0] sky130_fd_sc_hd__buf_4
x50[7] net37[7] vss vss vdd vdd phi27 sky130_fd_sc_hd__buf_8
x50[6] net37[6] vss vss vdd vdd phi26 sky130_fd_sc_hd__buf_8
x50[5] net37[5] vss vss vdd vdd phi25 sky130_fd_sc_hd__buf_8
x50[4] net37[4] vss vss vdd vdd phi24 sky130_fd_sc_hd__buf_8
x50[3] net37[3] vss vss vdd vdd phi23 sky130_fd_sc_hd__buf_8
x50[2] net37[2] vss vss vdd vdd phi22 sky130_fd_sc_hd__buf_8
x50[1] net37[1] vss vss vdd vdd phi21 sky130_fd_sc_hd__buf_8
x50[0] net37[0] vss vss vdd vdd phi20 sky130_fd_sc_hd__buf_8
x51[7] phi27 vss vss vdd vdd phi2_n7 sky130_fd_sc_hd__inv_8
x51[6] phi26 vss vss vdd vdd phi2_n6 sky130_fd_sc_hd__inv_8
x51[5] phi25 vss vss vdd vdd phi2_n5 sky130_fd_sc_hd__inv_8
x51[4] phi24 vss vss vdd vdd phi2_n4 sky130_fd_sc_hd__inv_8
x51[3] phi23 vss vss vdd vdd phi2_n3 sky130_fd_sc_hd__inv_8
x51[2] phi22 vss vss vdd vdd phi2_n2 sky130_fd_sc_hd__inv_8
x51[1] phi21 vss vss vdd vdd phi2_n1 sky130_fd_sc_hd__inv_8
x51[0] phi20 vss vss vdd vdd phi2_n0 sky130_fd_sc_hd__inv_8
x52[7] phi17 vss vss vdd vdd phi1_n7 sky130_fd_sc_hd__inv_8
x52[6] phi16 vss vss vdd vdd phi1_n6 sky130_fd_sc_hd__inv_8
x52[5] phi15 vss vss vdd vdd phi1_n5 sky130_fd_sc_hd__inv_8
x52[4] phi14 vss vss vdd vdd phi1_n4 sky130_fd_sc_hd__inv_8
x52[3] phi13 vss vss vdd vdd phi1_n3 sky130_fd_sc_hd__inv_8
x52[2] phi12 vss vss vdd vdd phi1_n2 sky130_fd_sc_hd__inv_8
x52[1] phi11 vss vss vdd vdd phi1_n1 sky130_fd_sc_hd__inv_8
x52[0] phi10 vss vss vdd vdd phi1_n0 sky130_fd_sc_hd__inv_8
x66 net8 vss vss vdd vdd net38 sky130_fd_sc_hd__buf_1
x67 net38 vss vss vdd vdd net39 sky130_fd_sc_hd__buf_2
x71 net39 vss vss vdd vdd net40 sky130_fd_sc_hd__buf_4
x73 net40 vss vss vdd vdd phi1x7 sky130_fd_sc_hd__buf_8
x53[6] net21[6] vss vss vdd vdd net41[6] sky130_fd_sc_hd__buf_1
x53[5] net21[5] vss vss vdd vdd net41[5] sky130_fd_sc_hd__buf_1
x53[4] net21[4] vss vss vdd vdd net41[4] sky130_fd_sc_hd__buf_1
x53[3] net21[3] vss vss vdd vdd net41[3] sky130_fd_sc_hd__buf_1
x53[2] net21[2] vss vss vdd vdd net41[2] sky130_fd_sc_hd__buf_1
x53[1] net21[1] vss vss vdd vdd net41[1] sky130_fd_sc_hd__buf_1
x53[0] net21[0] vss vss vdd vdd net41[0] sky130_fd_sc_hd__buf_1
x54[6] net41[6] vss vss vdd vdd net42[6] sky130_fd_sc_hd__buf_2
x54[5] net41[5] vss vss vdd vdd net42[5] sky130_fd_sc_hd__buf_2
x54[4] net41[4] vss vss vdd vdd net42[4] sky130_fd_sc_hd__buf_2
x54[3] net41[3] vss vss vdd vdd net42[3] sky130_fd_sc_hd__buf_2
x54[2] net41[2] vss vss vdd vdd net42[2] sky130_fd_sc_hd__buf_2
x54[1] net41[1] vss vss vdd vdd net42[1] sky130_fd_sc_hd__buf_2
x54[0] net41[0] vss vss vdd vdd net42[0] sky130_fd_sc_hd__buf_2
x55[6] net42[6] vss vss vdd vdd net43[6] sky130_fd_sc_hd__buf_4
x55[5] net42[5] vss vss vdd vdd net43[5] sky130_fd_sc_hd__buf_4
x55[4] net42[4] vss vss vdd vdd net43[4] sky130_fd_sc_hd__buf_4
x55[3] net42[3] vss vss vdd vdd net43[3] sky130_fd_sc_hd__buf_4
x55[2] net42[2] vss vss vdd vdd net43[2] sky130_fd_sc_hd__buf_4
x55[1] net42[1] vss vss vdd vdd net43[1] sky130_fd_sc_hd__buf_4
x55[0] net42[0] vss vss vdd vdd net43[0] sky130_fd_sc_hd__buf_4
x56[6] net43[6] vss vss vdd vdd phi1x6 sky130_fd_sc_hd__buf_8
x56[5] net43[5] vss vss vdd vdd phi1x5 sky130_fd_sc_hd__buf_8
x56[4] net43[4] vss vss vdd vdd phi1x4 sky130_fd_sc_hd__buf_8
x56[3] net43[3] vss vss vdd vdd phi1x3 sky130_fd_sc_hd__buf_8
x56[2] net43[2] vss vss vdd vdd phi1x2 sky130_fd_sc_hd__buf_8
x56[1] net43[1] vss vss vdd vdd phi1x1 sky130_fd_sc_hd__buf_8
x56[0] net43[0] vss vss vdd vdd phi1x0 sky130_fd_sc_hd__buf_8
x57[6] net30[6] vss vss vdd vdd net44[6] sky130_fd_sc_hd__buf_1
x57[5] net30[5] vss vss vdd vdd net44[5] sky130_fd_sc_hd__buf_1
x57[4] net30[4] vss vss vdd vdd net44[4] sky130_fd_sc_hd__buf_1
x57[3] net30[3] vss vss vdd vdd net44[3] sky130_fd_sc_hd__buf_1
x57[2] net30[2] vss vss vdd vdd net44[2] sky130_fd_sc_hd__buf_1
x57[1] net30[1] vss vss vdd vdd net44[1] sky130_fd_sc_hd__buf_1
x57[0] net30[0] vss vss vdd vdd net44[0] sky130_fd_sc_hd__buf_1
x58[6] net44[6] vss vss vdd vdd net45[6] sky130_fd_sc_hd__buf_2
x58[5] net44[5] vss vss vdd vdd net45[5] sky130_fd_sc_hd__buf_2
x58[4] net44[4] vss vss vdd vdd net45[4] sky130_fd_sc_hd__buf_2
x58[3] net44[3] vss vss vdd vdd net45[3] sky130_fd_sc_hd__buf_2
x58[2] net44[2] vss vss vdd vdd net45[2] sky130_fd_sc_hd__buf_2
x58[1] net44[1] vss vss vdd vdd net45[1] sky130_fd_sc_hd__buf_2
x58[0] net44[0] vss vss vdd vdd net45[0] sky130_fd_sc_hd__buf_2
x59[6] net45[6] vss vss vdd vdd net46[6] sky130_fd_sc_hd__buf_4
x59[5] net45[5] vss vss vdd vdd net46[5] sky130_fd_sc_hd__buf_4
x59[4] net45[4] vss vss vdd vdd net46[4] sky130_fd_sc_hd__buf_4
x59[3] net45[3] vss vss vdd vdd net46[3] sky130_fd_sc_hd__buf_4
x59[2] net45[2] vss vss vdd vdd net46[2] sky130_fd_sc_hd__buf_4
x59[1] net45[1] vss vss vdd vdd net46[1] sky130_fd_sc_hd__buf_4
x59[0] net45[0] vss vss vdd vdd net46[0] sky130_fd_sc_hd__buf_4
x60[6] net46[6] vss vss vdd vdd phi2x6 sky130_fd_sc_hd__buf_8
x60[5] net46[5] vss vss vdd vdd phi2x5 sky130_fd_sc_hd__buf_8
x60[4] net46[4] vss vss vdd vdd phi2x4 sky130_fd_sc_hd__buf_8
x60[3] net46[3] vss vss vdd vdd phi2x3 sky130_fd_sc_hd__buf_8
x60[2] net46[2] vss vss vdd vdd phi2x2 sky130_fd_sc_hd__buf_8
x60[1] net46[1] vss vss vdd vdd phi2x1 sky130_fd_sc_hd__buf_8
x60[0] net46[0] vss vss vdd vdd phi2x0 sky130_fd_sc_hd__buf_8
x74 net31 vss vss vdd vdd net47 sky130_fd_sc_hd__buf_1
x75 net47 vss vss vdd vdd net48 sky130_fd_sc_hd__buf_2
x76 net48 vss vss vdd vdd net49 sky130_fd_sc_hd__buf_4
x78 net49 vss vss vdd vdd phi2x7 sky130_fd_sc_hd__buf_8
x79 phi2x7 vss vss vdd vdd phi2x_n7 sky130_fd_sc_hd__inv_8
x61[6] phi2x6 vss vss vdd vdd phi2x_n6 sky130_fd_sc_hd__inv_8
x61[5] phi2x5 vss vss vdd vdd phi2x_n5 sky130_fd_sc_hd__inv_8
x61[4] phi2x4 vss vss vdd vdd phi2x_n4 sky130_fd_sc_hd__inv_8
x61[3] phi2x3 vss vss vdd vdd phi2x_n3 sky130_fd_sc_hd__inv_8
x61[2] phi2x2 vss vss vdd vdd phi2x_n2 sky130_fd_sc_hd__inv_8
x61[1] phi2x1 vss vss vdd vdd phi2x_n1 sky130_fd_sc_hd__inv_8
x61[0] phi2x0 vss vss vdd vdd phi2x_n0 sky130_fd_sc_hd__inv_8
x80 phi1x7 vss vss vdd vdd phi1x_n7 sky130_fd_sc_hd__inv_8
x62[6] phi1x6 vss vss vdd vdd phi1x_n6 sky130_fd_sc_hd__inv_8
x62[5] phi1x5 vss vss vdd vdd phi1x_n5 sky130_fd_sc_hd__inv_8
x62[4] phi1x4 vss vss vdd vdd phi1x_n4 sky130_fd_sc_hd__inv_8
x62[3] phi1x3 vss vss vdd vdd phi1x_n3 sky130_fd_sc_hd__inv_8
x62[2] phi1x2 vss vss vdd vdd phi1x_n2 sky130_fd_sc_hd__inv_8
x62[1] phi1x1 vss vss vdd vdd phi1x_n1 sky130_fd_sc_hd__inv_8
x62[0] phi1x0 vss vss vdd vdd phi1x_n0 sky130_fd_sc_hd__inv_8
x81 net12 vss vss vdd vdd net50 sky130_fd_sc_hd__buf_1
x82 net50 vss vss vdd vdd net51 sky130_fd_sc_hd__buf_2
x83 net51 vss vss vdd vdd net52 sky130_fd_sc_hd__buf_4
x84 net52 vss vss vdd vdd sphi1 sky130_fd_sc_hd__buf_8
x85 net11 vss vss vdd vdd net53 sky130_fd_sc_hd__buf_1
x86 net53 vss vss vdd vdd net54 sky130_fd_sc_hd__buf_2
x87 net54 vss vss vdd vdd net55 sky130_fd_sc_hd__buf_4
x88 net55 vss vss vdd vdd sphi2 sky130_fd_sc_hd__buf_8
x89 sphi1 vss vss vdd vdd sphi1_n sky130_fd_sc_hd__inv_8
x90 sphi2 vss vss vdd vdd sphi2_n sky130_fd_sc_hd__inv_8
x3[7] data_n7 vss vss vdd vdd dout7 sky130_fd_sc_hd__inv_4
x3[6] data_n6 vss vss vdd vdd dout6 sky130_fd_sc_hd__inv_4
x3[5] data_n5 vss vss vdd vdd dout5 sky130_fd_sc_hd__inv_4
x3[4] data_n4 vss vss vdd vdd dout4 sky130_fd_sc_hd__inv_4
x3[3] data_n3 vss vss vdd vdd dout3 sky130_fd_sc_hd__inv_4
x3[2] data_n2 vss vss vdd vdd dout2 sky130_fd_sc_hd__inv_4
x3[1] data_n1 vss vss vdd vdd dout1 sky130_fd_sc_hd__inv_4
x3[0] data_n0 vss vss vdd vdd dout0 sky130_fd_sc_hd__inv_4
.ends


* expanding   symbol:  /foss/designs/test/design/cap_switch_block.sym # of pins=9
** sym_path: /foss/designs/test/design/cap_switch_block.sym
** sch_path: /foss/designs/test/design/cap_switch_block.sch
.subckt cap_switch_block Vin sub GND Vdd phi1 phi2 phi2_n phi1_n com_x
*.ipin Vin
*.opin com_x
*.ipin phi1
*.ipin phi1_n
*.iopin Vdd
*.iopin GND
*.iopin sub
*.ipin phi2
*.ipin phi2_n
XC9 com_x net1 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 MF=1 m=1
x1 phi1 sub net1 Vin Vdd phi1_n tg_final
x2 phi2 sub net1 GND Vdd phi2_n tg_final
.ends


* expanding   symbol:  /foss/designs/test/design/tg_final.sym # of pins=6
** sym_path: /foss/designs/test/design/tg_final.sym
** sch_path: /foss/designs/test/design/tg_final.sch
.subckt tg_final clk sub vout vin vdd clk_b
*.ipin clk
*.ipin vin
*.opin vout
*.ipin vdd
*.ipin sub
*.ipin clk_b
XM2 vout clk vin sub sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 vout clk_b vin vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/test/design/sar_controller.sym # of pins=10
** sym_path: /foss/designs/test/design/sar_controller.sym
** sch_path: /foss/designs/test/design/sar_controller.sch
.subckt sar_controller clk data_rdy smpl rst_n smpl_n comp_out vss vdd d7 d6 d5 d4 d3 d2 d1 d0 d_n7 d_n6 d_n5 d_n4 d_n3 d_n2 d_n1
+ d_n0
*.ipin rst_n
*.opin data_rdy
*.ipin clk
*.ipin comp_out
*.iopin vss
*.iopin vdd
*.opin d7,d6,d5,d4,d3,d2,d1,d0
*.opin d_n7,d_n6,d_n5,d_n4,d_n3,d_n2,d_n1,d_n0
*.opin smpl_n
*.opin smpl
x26 net2 net21 net22 net9 vss vss vdd vdd net1 net25 sky130_fd_sc_hd__dfbbp_1
x5 net19 net23 net20 vss vss vdd vdd cnv_7 net9 sky130_fd_sc_hd__dfrbp_1
* noconn #net33
x24 net19 net8 net20 vss vss vdd vdd net23 net24 sky130_fd_sc_hd__dfsbp_1
x6 net24 net20 vss vss vdd vdd net22 sky130_fd_sc_hd__and2_4
x1 net19 cnv_7 net20 vss vss vdd vdd cnv_6 net12 sky130_fd_sc_hd__dfrbp_1
x2 net19 cnv_6 net20 vss vss vdd vdd cnv_5 net13 sky130_fd_sc_hd__dfrbp_1
x3 net19 cnv_5 net20 vss vss vdd vdd cnv_4 net14 sky130_fd_sc_hd__dfrbp_1
x4 net19 cnv_4 net20 vss vss vdd vdd cnv_3 net15 sky130_fd_sc_hd__dfrbp_1
x7 net19 cnv_3 net20 vss vss vdd vdd cnv_2 net16 sky130_fd_sc_hd__dfrbp_1
x8 net19 cnv_2 net20 vss vss vdd vdd cnv_1 net17 sky130_fd_sc_hd__dfrbp_1
x9 net19 cnv_1 net20 vss vss vdd vdd cnv_0 net18 sky130_fd_sc_hd__dfrbp_1
x10 net19 cnv_0 net20 vss vss vdd vdd net8 net33 sky130_fd_sc_hd__dfrbp_1
x11 vss vss net22 vss vss vdd vdd net11 net34 sky130_fd_sc_hd__dfrbp_1
x12 net10 net21 net22 net12 vss vss vdd vdd net2 net26 sky130_fd_sc_hd__dfbbp_1
x13 net3 net21 net22 net13 vss vss vdd vdd net10 net27 sky130_fd_sc_hd__dfbbp_1
x14 net4 net21 net22 net14 vss vss vdd vdd net3 net28 sky130_fd_sc_hd__dfbbp_1
x15 net5 net21 net22 net15 vss vss vdd vdd net4 net29 sky130_fd_sc_hd__dfbbp_1
x16 net6 net21 net22 net16 vss vss vdd vdd net5 net30 sky130_fd_sc_hd__dfbbp_1
x17 net7 net21 net22 net17 vss vss vdd vdd net6 net31 sky130_fd_sc_hd__dfbbp_1
x18 net11 net21 net22 net18 vss vss vdd vdd net7 net32 sky130_fd_sc_hd__dfbbp_1
* noconn #net34
x19 net1 vss vss vdd vdd d7 sky130_fd_sc_hd__buf_2
x20 net25 vss vss vdd vdd d_n7 sky130_fd_sc_hd__buf_2
x21 net2 vss vss vdd vdd d6 sky130_fd_sc_hd__buf_2
x22 net26 vss vss vdd vdd d_n6 sky130_fd_sc_hd__buf_2
x23 net10 vss vss vdd vdd d5 sky130_fd_sc_hd__buf_2
x25 net27 vss vss vdd vdd d_n5 sky130_fd_sc_hd__buf_2
x27 net3 vss vss vdd vdd d4 sky130_fd_sc_hd__buf_2
x28 net28 vss vss vdd vdd d_n4 sky130_fd_sc_hd__buf_2
x29 net4 vss vss vdd vdd d3 sky130_fd_sc_hd__buf_2
x30 net29 vss vss vdd vdd d_n3 sky130_fd_sc_hd__buf_2
x31 net5 vss vss vdd vdd d2 sky130_fd_sc_hd__buf_2
x32 net30 vss vss vdd vdd d_n2 sky130_fd_sc_hd__buf_2
x33 net6 vss vss vdd vdd d1 sky130_fd_sc_hd__buf_2
x34 net31 vss vss vdd vdd d_n1 sky130_fd_sc_hd__buf_2
x35 net7 vss vss vdd vdd d0 sky130_fd_sc_hd__buf_2
x36 net32 vss vss vdd vdd d_n0 sky130_fd_sc_hd__buf_2
x37 net23 vss vss vdd vdd net35 sky130_fd_sc_hd__buf_2
x38 net24 vss vss vdd vdd net36 sky130_fd_sc_hd__buf_2
x39 net8 vss vss vdd vdd data_rdy sky130_fd_sc_hd__buf_2
x40 comp_out vss vss vdd vdd net21 sky130_fd_sc_hd__buf_4
x41 rst_n vss vss vdd vdd net20 sky130_fd_sc_hd__buf_4
x42 clk vss vss vdd vdd net19 sky130_fd_sc_hd__buf_4
x43 net35 vss vss vdd vdd net37 sky130_fd_sc_hd__buf_4
x44 net36 vss vss vdd vdd net38 sky130_fd_sc_hd__buf_4
x45 net37 vss vss vdd vdd smpl sky130_fd_sc_hd__buf_8
x46 net38 vss vss vdd vdd smpl_n sky130_fd_sc_hd__buf_8
.ends

.end
