magic
tech sky130A
magscale 1 2
timestamp 1730649634
<< error_s >>
rect 3730 27460 3840 27520
rect 8720 27460 8830 27520
rect 13710 27460 13820 27520
rect 18700 27460 18810 27520
rect 23690 27460 23800 27520
rect 28680 27460 28790 27520
rect 33670 27460 33780 27520
rect 38660 27460 38770 27520
rect 43650 27460 43760 27520
rect 48640 27460 48750 27520
rect 53630 27460 53740 27520
rect 58620 27460 58730 27520
rect 63610 27460 63720 27520
rect 68600 27460 68710 27520
rect 73590 27460 73700 27520
rect 78580 27460 78690 27520
rect 3780 27420 3840 27460
rect 8770 27420 8830 27460
rect 13760 27420 13820 27460
rect 18750 27420 18810 27460
rect 23740 27420 23800 27460
rect 28730 27420 28790 27460
rect 33720 27420 33780 27460
rect 38710 27420 38770 27460
rect 43700 27420 43760 27460
rect 48690 27420 48750 27460
rect 53680 27420 53740 27460
rect 58670 27420 58730 27460
rect 63660 27420 63720 27460
rect 68650 27420 68710 27460
rect 73640 27420 73700 27460
rect 78630 27420 78690 27460
<< nwell >>
rect 3210 27858 3778 28590
rect 8200 27858 8768 28590
rect 13190 27858 13758 28590
rect 18180 27858 18748 28590
rect 23170 27858 23738 28590
rect 28160 27858 28728 28590
rect 33150 27858 33718 28590
rect 38140 27858 38708 28590
rect 43130 27858 43698 28590
rect 48120 27858 48688 28590
rect 53110 27858 53678 28590
rect 58100 27858 58668 28590
rect 63090 27858 63658 28590
rect 68080 27858 68648 28590
rect 73070 27858 73638 28590
rect 78060 27858 78628 28590
rect 82780 27858 83348 28590
rect 82780 26148 83348 26880
rect 82780 24438 83348 25170
rect -1510 22728 -942 23460
rect 82780 22728 83348 23460
rect -1510 21018 -942 21750
rect 82780 21018 83348 21750
rect -1510 19308 -942 20040
rect 82780 19308 83348 20040
rect -1510 17598 -942 18330
rect 82780 17598 83348 18330
rect -1510 15888 -942 16620
rect 82780 15888 83348 16620
rect -1510 14178 -942 14910
rect 82780 14178 83348 14910
rect -1510 12468 -942 13200
rect 82780 12468 83348 13200
rect -1510 10758 -942 11490
rect 82780 10758 83348 11490
rect -1510 9048 -942 9780
rect 82780 9048 83348 9780
rect -1510 7338 -942 8070
rect 82780 7338 83348 8070
rect -1510 5628 -942 6360
rect 82780 5628 83348 6360
rect -1510 3918 -942 4650
rect 82780 3918 83348 4650
rect -1510 2208 -942 2940
rect 82780 2208 83348 2940
rect -1510 498 -942 1230
rect 82780 498 83348 1230
rect -1510 -1212 -942 -480
rect 3210 -1212 3778 -480
rect 8200 -1212 8768 -480
rect 13190 -1212 13758 -480
rect 18180 -1212 18748 -480
rect 23170 -1212 23738 -480
rect 28160 -1212 28728 -480
rect 33150 -1212 33718 -480
rect 38140 -1212 38708 -480
rect 43130 -1212 43698 -480
rect 48120 -1212 48688 -480
rect 53110 -1212 53678 -480
rect 58100 -1212 58668 -480
rect 63090 -1212 63658 -480
rect 68080 -1212 68648 -480
rect 73070 -1212 73638 -480
rect 78060 -1212 78628 -480
rect 82780 -1212 83348 -480
<< pwell >>
rect -6370 29900 -6300 29990
rect 2650 27858 3208 28590
rect 7640 27858 8198 28590
rect 12630 27858 13188 28590
rect 17620 27858 18178 28590
rect 22610 27858 23168 28590
rect 27600 27858 28158 28590
rect 32590 27858 33148 28590
rect 37580 27858 38138 28590
rect 42570 27858 43128 28590
rect 47560 27858 48118 28590
rect 52550 27858 53108 28590
rect 57540 27858 58098 28590
rect 62530 27858 63088 28590
rect 67520 27858 68078 28590
rect 72510 27858 73068 28590
rect 77500 27858 78058 28590
rect 82220 27858 82778 28590
rect 2640 27360 2710 27820
rect 7630 27360 7700 27820
rect 12620 27360 12690 27820
rect 17610 27360 17680 27820
rect 22600 27360 22670 27820
rect 27590 27360 27660 27820
rect 32580 27360 32650 27820
rect 37570 27360 37640 27820
rect 42560 27360 42630 27820
rect 47550 27360 47620 27820
rect 52540 27360 52610 27820
rect 57530 27360 57600 27820
rect 62520 27360 62590 27820
rect 67510 27360 67580 27820
rect 72500 27360 72570 27820
rect 77490 27360 77560 27820
rect 82210 27360 82280 27820
rect 82220 26148 82778 26880
rect 82210 25650 82280 26110
rect 82220 24438 82778 25170
rect 82210 23940 82280 24400
rect -2070 22728 -1512 23460
rect 82220 22728 82778 23460
rect -2080 22230 -2010 22690
rect 82210 22230 82280 22690
rect -2070 21018 -1512 21750
rect 82220 21018 82778 21750
rect -2080 20520 -2010 20980
rect 82210 20520 82280 20980
rect -2070 19308 -1512 20040
rect 82220 19308 82778 20040
rect -2080 18810 -2010 19270
rect 82210 18810 82280 19270
rect -2070 17598 -1512 18330
rect 82220 17598 82778 18330
rect -2080 17100 -2010 17560
rect 82210 17100 82280 17560
rect -2070 15888 -1512 16620
rect 82220 15888 82778 16620
rect -2080 15390 -2010 15850
rect 82210 15390 82280 15850
rect -2070 14178 -1512 14910
rect 82220 14178 82778 14910
rect -2080 13680 -2010 14140
rect 82210 13680 82280 14140
rect -2070 12468 -1512 13200
rect 82220 12468 82778 13200
rect -2080 11970 -2010 12430
rect 82210 11970 82280 12430
rect -2070 10758 -1512 11490
rect 82220 10758 82778 11490
rect -2080 10260 -2010 10720
rect 82210 10260 82280 10720
rect -2070 9048 -1512 9780
rect 82220 9048 82778 9780
rect -2080 8550 -2010 9010
rect 82210 8550 82280 9010
rect -2070 7338 -1512 8070
rect 82220 7338 82778 8070
rect -2080 6840 -2010 7300
rect 82210 6840 82280 7300
rect -2070 5628 -1512 6360
rect 82220 5628 82778 6360
rect -2080 5130 -2010 5590
rect 82210 5130 82280 5590
rect -2070 3918 -1512 4650
rect 82220 3918 82778 4650
rect -2080 3420 -2010 3880
rect 82210 3420 82280 3880
rect -2070 2208 -1512 2940
rect 82220 2208 82778 2940
rect -2080 1710 -2010 2170
rect 82210 1710 82280 2170
rect -2070 498 -1512 1230
rect 82220 498 82778 1230
rect -2080 150 -2010 460
rect 82210 150 82280 460
rect -2080 70 -2000 150
rect 2640 70 2720 150
rect 7630 70 7710 150
rect 12620 70 12700 150
rect 17610 70 17690 150
rect 22600 70 22680 150
rect 27590 70 27670 150
rect 32580 70 32660 150
rect 37570 70 37650 150
rect 42560 70 42640 150
rect 47550 70 47630 150
rect 52540 70 52620 150
rect 57530 70 57610 150
rect 62520 70 62600 150
rect 67510 70 67590 150
rect 72500 70 72580 150
rect 77490 70 77570 150
rect 82210 70 82290 150
rect -2080 0 -2010 70
rect 2640 0 2710 70
rect 7630 0 7700 70
rect 12620 0 12690 70
rect 17610 0 17680 70
rect 22600 0 22670 70
rect 27590 0 27660 70
rect 32580 0 32650 70
rect 37570 0 37640 70
rect 42560 0 42630 70
rect 47550 0 47620 70
rect 52540 0 52610 70
rect 57530 0 57600 70
rect 62520 0 62590 70
rect 67510 0 67580 70
rect 72500 0 72570 70
rect 77490 0 77560 70
rect 82210 0 82280 70
rect -2070 -1212 -1512 -480
rect 2650 -1212 3208 -480
rect 7640 -1212 8198 -480
rect 12630 -1212 13188 -480
rect 17620 -1212 18178 -480
rect 22610 -1212 23168 -480
rect 27600 -1212 28158 -480
rect 32590 -1212 33148 -480
rect 37580 -1212 38138 -480
rect 42570 -1212 43128 -480
rect 47560 -1212 48118 -480
rect 52550 -1212 53108 -480
rect 57540 -1212 58098 -480
rect 62530 -1212 63088 -480
rect 67520 -1212 68078 -480
rect 72510 -1212 73068 -480
rect 77500 -1212 78058 -480
rect 82220 -1212 82778 -480
rect -2080 -1710 -2010 -1250
rect 2640 -1710 2710 -1250
rect 7630 -1710 7700 -1250
rect 12620 -1710 12690 -1250
rect 17610 -1710 17680 -1250
rect 22600 -1710 22670 -1250
rect 27590 -1710 27660 -1250
rect 32580 -1710 32650 -1250
rect 37570 -1710 37640 -1250
rect 42560 -1710 42630 -1250
rect 47550 -1710 47620 -1250
rect 52540 -1710 52610 -1250
rect 57530 -1710 57600 -1250
rect 62520 -1710 62590 -1250
rect 67510 -1710 67580 -1250
rect 72500 -1710 72570 -1250
rect 77490 -1710 77560 -1250
rect 82210 -1710 82280 -1250
<< nmos >>
rect 2860 28364 3060 28394
rect 2860 28054 3060 28084
rect 7850 28364 8050 28394
rect 7850 28054 8050 28084
rect 12840 28364 13040 28394
rect 12840 28054 13040 28084
rect 17830 28364 18030 28394
rect 17830 28054 18030 28084
rect 22820 28364 23020 28394
rect 22820 28054 23020 28084
rect 27810 28364 28010 28394
rect 27810 28054 28010 28084
rect 32800 28364 33000 28394
rect 32800 28054 33000 28084
rect 37790 28364 37990 28394
rect 37790 28054 37990 28084
rect 42780 28364 42980 28394
rect 42780 28054 42980 28084
rect 47770 28364 47970 28394
rect 47770 28054 47970 28084
rect 52760 28364 52960 28394
rect 52760 28054 52960 28084
rect 57750 28364 57950 28394
rect 57750 28054 57950 28084
rect 62740 28364 62940 28394
rect 62740 28054 62940 28084
rect 67730 28364 67930 28394
rect 67730 28054 67930 28084
rect 72720 28364 72920 28394
rect 72720 28054 72920 28084
rect 77710 28364 77910 28394
rect 77710 28054 77910 28084
rect 82430 28364 82630 28394
rect 82430 28054 82630 28084
rect 82430 26654 82630 26684
rect 82430 26344 82630 26374
rect 82430 24944 82630 24974
rect 82430 24634 82630 24664
rect -1860 23234 -1660 23264
rect -1860 22924 -1660 22954
rect 82430 23234 82630 23264
rect 82430 22924 82630 22954
rect -1860 21524 -1660 21554
rect -1860 21214 -1660 21244
rect 82430 21524 82630 21554
rect 82430 21214 82630 21244
rect -1860 19814 -1660 19844
rect -1860 19504 -1660 19534
rect 82430 19814 82630 19844
rect 82430 19504 82630 19534
rect -1860 18104 -1660 18134
rect -1860 17794 -1660 17824
rect 82430 18104 82630 18134
rect 82430 17794 82630 17824
rect -1860 16394 -1660 16424
rect -1860 16084 -1660 16114
rect 82430 16394 82630 16424
rect 82430 16084 82630 16114
rect -1860 14684 -1660 14714
rect -1860 14374 -1660 14404
rect 82430 14684 82630 14714
rect 82430 14374 82630 14404
rect -1860 12974 -1660 13004
rect -1860 12664 -1660 12694
rect 82430 12974 82630 13004
rect 82430 12664 82630 12694
rect -1860 11264 -1660 11294
rect -1860 10954 -1660 10984
rect 82430 11264 82630 11294
rect 82430 10954 82630 10984
rect -1860 9554 -1660 9584
rect -1860 9244 -1660 9274
rect 82430 9554 82630 9584
rect 82430 9244 82630 9274
rect -1860 7844 -1660 7874
rect -1860 7534 -1660 7564
rect 82430 7844 82630 7874
rect 82430 7534 82630 7564
rect -1860 6134 -1660 6164
rect -1860 5824 -1660 5854
rect 82430 6134 82630 6164
rect 82430 5824 82630 5854
rect -1860 4424 -1660 4454
rect -1860 4114 -1660 4144
rect 82430 4424 82630 4454
rect 82430 4114 82630 4144
rect -1860 2714 -1660 2744
rect -1860 2404 -1660 2434
rect 82430 2714 82630 2744
rect 82430 2404 82630 2434
rect -1860 1004 -1660 1034
rect -1860 694 -1660 724
rect 82430 1004 82630 1034
rect 82430 694 82630 724
rect -1860 -706 -1660 -676
rect -1860 -1016 -1660 -986
rect 2860 -706 3060 -676
rect 2860 -1016 3060 -986
rect 7850 -706 8050 -676
rect 7850 -1016 8050 -986
rect 12840 -706 13040 -676
rect 12840 -1016 13040 -986
rect 17830 -706 18030 -676
rect 17830 -1016 18030 -986
rect 22820 -706 23020 -676
rect 22820 -1016 23020 -986
rect 27810 -706 28010 -676
rect 27810 -1016 28010 -986
rect 32800 -706 33000 -676
rect 32800 -1016 33000 -986
rect 37790 -706 37990 -676
rect 37790 -1016 37990 -986
rect 42780 -706 42980 -676
rect 42780 -1016 42980 -986
rect 47770 -706 47970 -676
rect 47770 -1016 47970 -986
rect 52760 -706 52960 -676
rect 52760 -1016 52960 -986
rect 57750 -706 57950 -676
rect 57750 -1016 57950 -986
rect 62740 -706 62940 -676
rect 62740 -1016 62940 -986
rect 67730 -706 67930 -676
rect 67730 -1016 67930 -986
rect 72720 -706 72920 -676
rect 72720 -1016 72920 -986
rect 77710 -706 77910 -676
rect 77710 -1016 77910 -986
rect 82430 -706 82630 -676
rect 82430 -1016 82630 -986
<< pmos >>
rect 3358 28364 3558 28394
rect 3358 28054 3558 28084
rect 8348 28364 8548 28394
rect 8348 28054 8548 28084
rect 13338 28364 13538 28394
rect 13338 28054 13538 28084
rect 18328 28364 18528 28394
rect 18328 28054 18528 28084
rect 23318 28364 23518 28394
rect 23318 28054 23518 28084
rect 28308 28364 28508 28394
rect 28308 28054 28508 28084
rect 33298 28364 33498 28394
rect 33298 28054 33498 28084
rect 38288 28364 38488 28394
rect 38288 28054 38488 28084
rect 43278 28364 43478 28394
rect 43278 28054 43478 28084
rect 48268 28364 48468 28394
rect 48268 28054 48468 28084
rect 53258 28364 53458 28394
rect 53258 28054 53458 28084
rect 58248 28364 58448 28394
rect 58248 28054 58448 28084
rect 63238 28364 63438 28394
rect 63238 28054 63438 28084
rect 68228 28364 68428 28394
rect 68228 28054 68428 28084
rect 73218 28364 73418 28394
rect 73218 28054 73418 28084
rect 78208 28364 78408 28394
rect 78208 28054 78408 28084
rect 82928 28364 83128 28394
rect 82928 28054 83128 28084
rect 82928 26654 83128 26684
rect 82928 26344 83128 26374
rect 82928 24944 83128 24974
rect 82928 24634 83128 24664
rect -1362 23234 -1162 23264
rect -1362 22924 -1162 22954
rect 82928 23234 83128 23264
rect 82928 22924 83128 22954
rect -1362 21524 -1162 21554
rect -1362 21214 -1162 21244
rect 82928 21524 83128 21554
rect 82928 21214 83128 21244
rect -1362 19814 -1162 19844
rect -1362 19504 -1162 19534
rect 82928 19814 83128 19844
rect 82928 19504 83128 19534
rect -1362 18104 -1162 18134
rect -1362 17794 -1162 17824
rect 82928 18104 83128 18134
rect 82928 17794 83128 17824
rect -1362 16394 -1162 16424
rect -1362 16084 -1162 16114
rect 82928 16394 83128 16424
rect 82928 16084 83128 16114
rect -1362 14684 -1162 14714
rect -1362 14374 -1162 14404
rect 82928 14684 83128 14714
rect 82928 14374 83128 14404
rect -1362 12974 -1162 13004
rect -1362 12664 -1162 12694
rect 82928 12974 83128 13004
rect 82928 12664 83128 12694
rect -1362 11264 -1162 11294
rect -1362 10954 -1162 10984
rect 82928 11264 83128 11294
rect 82928 10954 83128 10984
rect -1362 9554 -1162 9584
rect -1362 9244 -1162 9274
rect 82928 9554 83128 9584
rect 82928 9244 83128 9274
rect -1362 7844 -1162 7874
rect -1362 7534 -1162 7564
rect 82928 7844 83128 7874
rect 82928 7534 83128 7564
rect -1362 6134 -1162 6164
rect -1362 5824 -1162 5854
rect 82928 6134 83128 6164
rect 82928 5824 83128 5854
rect -1362 4424 -1162 4454
rect -1362 4114 -1162 4144
rect 82928 4424 83128 4454
rect 82928 4114 83128 4144
rect -1362 2714 -1162 2744
rect -1362 2404 -1162 2434
rect 82928 2714 83128 2744
rect 82928 2404 83128 2434
rect -1362 1004 -1162 1034
rect -1362 694 -1162 724
rect 82928 1004 83128 1034
rect 82928 694 83128 724
rect -1362 -706 -1162 -676
rect -1362 -1016 -1162 -986
rect 3358 -706 3558 -676
rect 3358 -1016 3558 -986
rect 8348 -706 8548 -676
rect 8348 -1016 8548 -986
rect 13338 -706 13538 -676
rect 13338 -1016 13538 -986
rect 18328 -706 18528 -676
rect 18328 -1016 18528 -986
rect 23318 -706 23518 -676
rect 23318 -1016 23518 -986
rect 28308 -706 28508 -676
rect 28308 -1016 28508 -986
rect 33298 -706 33498 -676
rect 33298 -1016 33498 -986
rect 38288 -706 38488 -676
rect 38288 -1016 38488 -986
rect 43278 -706 43478 -676
rect 43278 -1016 43478 -986
rect 48268 -706 48468 -676
rect 48268 -1016 48468 -986
rect 53258 -706 53458 -676
rect 53258 -1016 53458 -986
rect 58248 -706 58448 -676
rect 58248 -1016 58448 -986
rect 63238 -706 63438 -676
rect 63238 -1016 63438 -986
rect 68228 -706 68428 -676
rect 68228 -1016 68428 -986
rect 73218 -706 73418 -676
rect 73218 -1016 73418 -986
rect 78208 -706 78408 -676
rect 78208 -1016 78408 -986
rect 82928 -706 83128 -676
rect 82928 -1016 83128 -986
<< ndiff >>
rect 2860 28440 3060 28452
rect 2860 28406 2872 28440
rect 3048 28406 3060 28440
rect 2860 28394 3060 28406
rect 2860 28352 3060 28364
rect 2860 28318 2872 28352
rect 3048 28318 3060 28352
rect 2860 28306 3060 28318
rect 2860 28130 3060 28142
rect 2860 28096 2872 28130
rect 3048 28096 3060 28130
rect 2860 28084 3060 28096
rect 2860 28042 3060 28054
rect 2860 28008 2872 28042
rect 3048 28008 3060 28042
rect 2860 27996 3060 28008
rect 7850 28440 8050 28452
rect 7850 28406 7862 28440
rect 8038 28406 8050 28440
rect 7850 28394 8050 28406
rect 7850 28352 8050 28364
rect 7850 28318 7862 28352
rect 8038 28318 8050 28352
rect 7850 28306 8050 28318
rect 7850 28130 8050 28142
rect 7850 28096 7862 28130
rect 8038 28096 8050 28130
rect 7850 28084 8050 28096
rect 7850 28042 8050 28054
rect 7850 28008 7862 28042
rect 8038 28008 8050 28042
rect 7850 27996 8050 28008
rect 12840 28440 13040 28452
rect 12840 28406 12852 28440
rect 13028 28406 13040 28440
rect 12840 28394 13040 28406
rect 12840 28352 13040 28364
rect 12840 28318 12852 28352
rect 13028 28318 13040 28352
rect 12840 28306 13040 28318
rect 12840 28130 13040 28142
rect 12840 28096 12852 28130
rect 13028 28096 13040 28130
rect 12840 28084 13040 28096
rect 12840 28042 13040 28054
rect 12840 28008 12852 28042
rect 13028 28008 13040 28042
rect 12840 27996 13040 28008
rect 17830 28440 18030 28452
rect 17830 28406 17842 28440
rect 18018 28406 18030 28440
rect 17830 28394 18030 28406
rect 17830 28352 18030 28364
rect 17830 28318 17842 28352
rect 18018 28318 18030 28352
rect 17830 28306 18030 28318
rect 17830 28130 18030 28142
rect 17830 28096 17842 28130
rect 18018 28096 18030 28130
rect 17830 28084 18030 28096
rect 17830 28042 18030 28054
rect 17830 28008 17842 28042
rect 18018 28008 18030 28042
rect 17830 27996 18030 28008
rect 22820 28440 23020 28452
rect 22820 28406 22832 28440
rect 23008 28406 23020 28440
rect 22820 28394 23020 28406
rect 22820 28352 23020 28364
rect 22820 28318 22832 28352
rect 23008 28318 23020 28352
rect 22820 28306 23020 28318
rect 22820 28130 23020 28142
rect 22820 28096 22832 28130
rect 23008 28096 23020 28130
rect 22820 28084 23020 28096
rect 22820 28042 23020 28054
rect 22820 28008 22832 28042
rect 23008 28008 23020 28042
rect 22820 27996 23020 28008
rect 27810 28440 28010 28452
rect 27810 28406 27822 28440
rect 27998 28406 28010 28440
rect 27810 28394 28010 28406
rect 27810 28352 28010 28364
rect 27810 28318 27822 28352
rect 27998 28318 28010 28352
rect 27810 28306 28010 28318
rect 27810 28130 28010 28142
rect 27810 28096 27822 28130
rect 27998 28096 28010 28130
rect 27810 28084 28010 28096
rect 27810 28042 28010 28054
rect 27810 28008 27822 28042
rect 27998 28008 28010 28042
rect 27810 27996 28010 28008
rect 32800 28440 33000 28452
rect 32800 28406 32812 28440
rect 32988 28406 33000 28440
rect 32800 28394 33000 28406
rect 32800 28352 33000 28364
rect 32800 28318 32812 28352
rect 32988 28318 33000 28352
rect 32800 28306 33000 28318
rect 32800 28130 33000 28142
rect 32800 28096 32812 28130
rect 32988 28096 33000 28130
rect 32800 28084 33000 28096
rect 32800 28042 33000 28054
rect 32800 28008 32812 28042
rect 32988 28008 33000 28042
rect 32800 27996 33000 28008
rect 37790 28440 37990 28452
rect 37790 28406 37802 28440
rect 37978 28406 37990 28440
rect 37790 28394 37990 28406
rect 37790 28352 37990 28364
rect 37790 28318 37802 28352
rect 37978 28318 37990 28352
rect 37790 28306 37990 28318
rect 37790 28130 37990 28142
rect 37790 28096 37802 28130
rect 37978 28096 37990 28130
rect 37790 28084 37990 28096
rect 37790 28042 37990 28054
rect 37790 28008 37802 28042
rect 37978 28008 37990 28042
rect 37790 27996 37990 28008
rect 42780 28440 42980 28452
rect 42780 28406 42792 28440
rect 42968 28406 42980 28440
rect 42780 28394 42980 28406
rect 42780 28352 42980 28364
rect 42780 28318 42792 28352
rect 42968 28318 42980 28352
rect 42780 28306 42980 28318
rect 42780 28130 42980 28142
rect 42780 28096 42792 28130
rect 42968 28096 42980 28130
rect 42780 28084 42980 28096
rect 42780 28042 42980 28054
rect 42780 28008 42792 28042
rect 42968 28008 42980 28042
rect 42780 27996 42980 28008
rect 47770 28440 47970 28452
rect 47770 28406 47782 28440
rect 47958 28406 47970 28440
rect 47770 28394 47970 28406
rect 47770 28352 47970 28364
rect 47770 28318 47782 28352
rect 47958 28318 47970 28352
rect 47770 28306 47970 28318
rect 47770 28130 47970 28142
rect 47770 28096 47782 28130
rect 47958 28096 47970 28130
rect 47770 28084 47970 28096
rect 47770 28042 47970 28054
rect 47770 28008 47782 28042
rect 47958 28008 47970 28042
rect 47770 27996 47970 28008
rect 52760 28440 52960 28452
rect 52760 28406 52772 28440
rect 52948 28406 52960 28440
rect 52760 28394 52960 28406
rect 52760 28352 52960 28364
rect 52760 28318 52772 28352
rect 52948 28318 52960 28352
rect 52760 28306 52960 28318
rect 52760 28130 52960 28142
rect 52760 28096 52772 28130
rect 52948 28096 52960 28130
rect 52760 28084 52960 28096
rect 52760 28042 52960 28054
rect 52760 28008 52772 28042
rect 52948 28008 52960 28042
rect 52760 27996 52960 28008
rect 57750 28440 57950 28452
rect 57750 28406 57762 28440
rect 57938 28406 57950 28440
rect 57750 28394 57950 28406
rect 57750 28352 57950 28364
rect 57750 28318 57762 28352
rect 57938 28318 57950 28352
rect 57750 28306 57950 28318
rect 57750 28130 57950 28142
rect 57750 28096 57762 28130
rect 57938 28096 57950 28130
rect 57750 28084 57950 28096
rect 57750 28042 57950 28054
rect 57750 28008 57762 28042
rect 57938 28008 57950 28042
rect 57750 27996 57950 28008
rect 62740 28440 62940 28452
rect 62740 28406 62752 28440
rect 62928 28406 62940 28440
rect 62740 28394 62940 28406
rect 62740 28352 62940 28364
rect 62740 28318 62752 28352
rect 62928 28318 62940 28352
rect 62740 28306 62940 28318
rect 62740 28130 62940 28142
rect 62740 28096 62752 28130
rect 62928 28096 62940 28130
rect 62740 28084 62940 28096
rect 62740 28042 62940 28054
rect 62740 28008 62752 28042
rect 62928 28008 62940 28042
rect 62740 27996 62940 28008
rect 67730 28440 67930 28452
rect 67730 28406 67742 28440
rect 67918 28406 67930 28440
rect 67730 28394 67930 28406
rect 67730 28352 67930 28364
rect 67730 28318 67742 28352
rect 67918 28318 67930 28352
rect 67730 28306 67930 28318
rect 67730 28130 67930 28142
rect 67730 28096 67742 28130
rect 67918 28096 67930 28130
rect 67730 28084 67930 28096
rect 67730 28042 67930 28054
rect 67730 28008 67742 28042
rect 67918 28008 67930 28042
rect 67730 27996 67930 28008
rect 72720 28440 72920 28452
rect 72720 28406 72732 28440
rect 72908 28406 72920 28440
rect 72720 28394 72920 28406
rect 72720 28352 72920 28364
rect 72720 28318 72732 28352
rect 72908 28318 72920 28352
rect 72720 28306 72920 28318
rect 72720 28130 72920 28142
rect 72720 28096 72732 28130
rect 72908 28096 72920 28130
rect 72720 28084 72920 28096
rect 72720 28042 72920 28054
rect 72720 28008 72732 28042
rect 72908 28008 72920 28042
rect 72720 27996 72920 28008
rect 77710 28440 77910 28452
rect 77710 28406 77722 28440
rect 77898 28406 77910 28440
rect 77710 28394 77910 28406
rect 77710 28352 77910 28364
rect 77710 28318 77722 28352
rect 77898 28318 77910 28352
rect 77710 28306 77910 28318
rect 77710 28130 77910 28142
rect 77710 28096 77722 28130
rect 77898 28096 77910 28130
rect 77710 28084 77910 28096
rect 77710 28042 77910 28054
rect 77710 28008 77722 28042
rect 77898 28008 77910 28042
rect 77710 27996 77910 28008
rect 82430 28440 82630 28452
rect 82430 28406 82442 28440
rect 82618 28406 82630 28440
rect 82430 28394 82630 28406
rect 82430 28352 82630 28364
rect 82430 28318 82442 28352
rect 82618 28318 82630 28352
rect 82430 28306 82630 28318
rect 82430 28130 82630 28142
rect 82430 28096 82442 28130
rect 82618 28096 82630 28130
rect 82430 28084 82630 28096
rect 82430 28042 82630 28054
rect 82430 28008 82442 28042
rect 82618 28008 82630 28042
rect 82430 27996 82630 28008
rect 82430 26730 82630 26742
rect 82430 26696 82442 26730
rect 82618 26696 82630 26730
rect 82430 26684 82630 26696
rect 82430 26642 82630 26654
rect 82430 26608 82442 26642
rect 82618 26608 82630 26642
rect 82430 26596 82630 26608
rect 82430 26420 82630 26432
rect 82430 26386 82442 26420
rect 82618 26386 82630 26420
rect 82430 26374 82630 26386
rect 82430 26332 82630 26344
rect 82430 26298 82442 26332
rect 82618 26298 82630 26332
rect 82430 26286 82630 26298
rect 82430 25020 82630 25032
rect 82430 24986 82442 25020
rect 82618 24986 82630 25020
rect 82430 24974 82630 24986
rect 82430 24932 82630 24944
rect 82430 24898 82442 24932
rect 82618 24898 82630 24932
rect 82430 24886 82630 24898
rect 82430 24710 82630 24722
rect 82430 24676 82442 24710
rect 82618 24676 82630 24710
rect 82430 24664 82630 24676
rect 82430 24622 82630 24634
rect 82430 24588 82442 24622
rect 82618 24588 82630 24622
rect 82430 24576 82630 24588
rect -1860 23310 -1660 23322
rect -1860 23276 -1848 23310
rect -1672 23276 -1660 23310
rect -1860 23264 -1660 23276
rect -1860 23222 -1660 23234
rect -1860 23188 -1848 23222
rect -1672 23188 -1660 23222
rect -1860 23176 -1660 23188
rect -1860 23000 -1660 23012
rect -1860 22966 -1848 23000
rect -1672 22966 -1660 23000
rect -1860 22954 -1660 22966
rect -1860 22912 -1660 22924
rect -1860 22878 -1848 22912
rect -1672 22878 -1660 22912
rect -1860 22866 -1660 22878
rect 82430 23310 82630 23322
rect 82430 23276 82442 23310
rect 82618 23276 82630 23310
rect 82430 23264 82630 23276
rect 82430 23222 82630 23234
rect 82430 23188 82442 23222
rect 82618 23188 82630 23222
rect 82430 23176 82630 23188
rect 82430 23000 82630 23012
rect 82430 22966 82442 23000
rect 82618 22966 82630 23000
rect 82430 22954 82630 22966
rect 82430 22912 82630 22924
rect 82430 22878 82442 22912
rect 82618 22878 82630 22912
rect 82430 22866 82630 22878
rect -1860 21600 -1660 21612
rect -1860 21566 -1848 21600
rect -1672 21566 -1660 21600
rect -1860 21554 -1660 21566
rect -1860 21512 -1660 21524
rect -1860 21478 -1848 21512
rect -1672 21478 -1660 21512
rect -1860 21466 -1660 21478
rect -1860 21290 -1660 21302
rect -1860 21256 -1848 21290
rect -1672 21256 -1660 21290
rect -1860 21244 -1660 21256
rect -1860 21202 -1660 21214
rect -1860 21168 -1848 21202
rect -1672 21168 -1660 21202
rect -1860 21156 -1660 21168
rect 82430 21600 82630 21612
rect 82430 21566 82442 21600
rect 82618 21566 82630 21600
rect 82430 21554 82630 21566
rect 82430 21512 82630 21524
rect 82430 21478 82442 21512
rect 82618 21478 82630 21512
rect 82430 21466 82630 21478
rect 82430 21290 82630 21302
rect 82430 21256 82442 21290
rect 82618 21256 82630 21290
rect 82430 21244 82630 21256
rect 82430 21202 82630 21214
rect 82430 21168 82442 21202
rect 82618 21168 82630 21202
rect 82430 21156 82630 21168
rect -1860 19890 -1660 19902
rect -1860 19856 -1848 19890
rect -1672 19856 -1660 19890
rect -1860 19844 -1660 19856
rect -1860 19802 -1660 19814
rect -1860 19768 -1848 19802
rect -1672 19768 -1660 19802
rect -1860 19756 -1660 19768
rect -1860 19580 -1660 19592
rect -1860 19546 -1848 19580
rect -1672 19546 -1660 19580
rect -1860 19534 -1660 19546
rect -1860 19492 -1660 19504
rect -1860 19458 -1848 19492
rect -1672 19458 -1660 19492
rect -1860 19446 -1660 19458
rect 82430 19890 82630 19902
rect 82430 19856 82442 19890
rect 82618 19856 82630 19890
rect 82430 19844 82630 19856
rect 82430 19802 82630 19814
rect 82430 19768 82442 19802
rect 82618 19768 82630 19802
rect 82430 19756 82630 19768
rect 82430 19580 82630 19592
rect 82430 19546 82442 19580
rect 82618 19546 82630 19580
rect 82430 19534 82630 19546
rect 82430 19492 82630 19504
rect 82430 19458 82442 19492
rect 82618 19458 82630 19492
rect 82430 19446 82630 19458
rect -1860 18180 -1660 18192
rect -1860 18146 -1848 18180
rect -1672 18146 -1660 18180
rect -1860 18134 -1660 18146
rect -1860 18092 -1660 18104
rect -1860 18058 -1848 18092
rect -1672 18058 -1660 18092
rect -1860 18046 -1660 18058
rect -1860 17870 -1660 17882
rect -1860 17836 -1848 17870
rect -1672 17836 -1660 17870
rect -1860 17824 -1660 17836
rect -1860 17782 -1660 17794
rect -1860 17748 -1848 17782
rect -1672 17748 -1660 17782
rect -1860 17736 -1660 17748
rect 82430 18180 82630 18192
rect 82430 18146 82442 18180
rect 82618 18146 82630 18180
rect 82430 18134 82630 18146
rect 82430 18092 82630 18104
rect 82430 18058 82442 18092
rect 82618 18058 82630 18092
rect 82430 18046 82630 18058
rect 82430 17870 82630 17882
rect 82430 17836 82442 17870
rect 82618 17836 82630 17870
rect 82430 17824 82630 17836
rect 82430 17782 82630 17794
rect 82430 17748 82442 17782
rect 82618 17748 82630 17782
rect 82430 17736 82630 17748
rect -1860 16470 -1660 16482
rect -1860 16436 -1848 16470
rect -1672 16436 -1660 16470
rect -1860 16424 -1660 16436
rect -1860 16382 -1660 16394
rect -1860 16348 -1848 16382
rect -1672 16348 -1660 16382
rect -1860 16336 -1660 16348
rect -1860 16160 -1660 16172
rect -1860 16126 -1848 16160
rect -1672 16126 -1660 16160
rect -1860 16114 -1660 16126
rect -1860 16072 -1660 16084
rect -1860 16038 -1848 16072
rect -1672 16038 -1660 16072
rect -1860 16026 -1660 16038
rect 82430 16470 82630 16482
rect 82430 16436 82442 16470
rect 82618 16436 82630 16470
rect 82430 16424 82630 16436
rect 82430 16382 82630 16394
rect 82430 16348 82442 16382
rect 82618 16348 82630 16382
rect 82430 16336 82630 16348
rect 82430 16160 82630 16172
rect 82430 16126 82442 16160
rect 82618 16126 82630 16160
rect 82430 16114 82630 16126
rect 82430 16072 82630 16084
rect 82430 16038 82442 16072
rect 82618 16038 82630 16072
rect 82430 16026 82630 16038
rect -1860 14760 -1660 14772
rect -1860 14726 -1848 14760
rect -1672 14726 -1660 14760
rect -1860 14714 -1660 14726
rect -1860 14672 -1660 14684
rect -1860 14638 -1848 14672
rect -1672 14638 -1660 14672
rect -1860 14626 -1660 14638
rect -1860 14450 -1660 14462
rect -1860 14416 -1848 14450
rect -1672 14416 -1660 14450
rect -1860 14404 -1660 14416
rect -1860 14362 -1660 14374
rect -1860 14328 -1848 14362
rect -1672 14328 -1660 14362
rect -1860 14316 -1660 14328
rect 82430 14760 82630 14772
rect 82430 14726 82442 14760
rect 82618 14726 82630 14760
rect 82430 14714 82630 14726
rect 82430 14672 82630 14684
rect 82430 14638 82442 14672
rect 82618 14638 82630 14672
rect 82430 14626 82630 14638
rect 82430 14450 82630 14462
rect 82430 14416 82442 14450
rect 82618 14416 82630 14450
rect 82430 14404 82630 14416
rect 82430 14362 82630 14374
rect 82430 14328 82442 14362
rect 82618 14328 82630 14362
rect 82430 14316 82630 14328
rect -1860 13050 -1660 13062
rect -1860 13016 -1848 13050
rect -1672 13016 -1660 13050
rect -1860 13004 -1660 13016
rect -1860 12962 -1660 12974
rect -1860 12928 -1848 12962
rect -1672 12928 -1660 12962
rect -1860 12916 -1660 12928
rect -1860 12740 -1660 12752
rect -1860 12706 -1848 12740
rect -1672 12706 -1660 12740
rect -1860 12694 -1660 12706
rect -1860 12652 -1660 12664
rect -1860 12618 -1848 12652
rect -1672 12618 -1660 12652
rect -1860 12606 -1660 12618
rect 82430 13050 82630 13062
rect 82430 13016 82442 13050
rect 82618 13016 82630 13050
rect 82430 13004 82630 13016
rect 82430 12962 82630 12974
rect 82430 12928 82442 12962
rect 82618 12928 82630 12962
rect 82430 12916 82630 12928
rect 82430 12740 82630 12752
rect 82430 12706 82442 12740
rect 82618 12706 82630 12740
rect 82430 12694 82630 12706
rect 82430 12652 82630 12664
rect 82430 12618 82442 12652
rect 82618 12618 82630 12652
rect 82430 12606 82630 12618
rect -1860 11340 -1660 11352
rect -1860 11306 -1848 11340
rect -1672 11306 -1660 11340
rect -1860 11294 -1660 11306
rect -1860 11252 -1660 11264
rect -1860 11218 -1848 11252
rect -1672 11218 -1660 11252
rect -1860 11206 -1660 11218
rect -1860 11030 -1660 11042
rect -1860 10996 -1848 11030
rect -1672 10996 -1660 11030
rect -1860 10984 -1660 10996
rect -1860 10942 -1660 10954
rect -1860 10908 -1848 10942
rect -1672 10908 -1660 10942
rect -1860 10896 -1660 10908
rect 82430 11340 82630 11352
rect 82430 11306 82442 11340
rect 82618 11306 82630 11340
rect 82430 11294 82630 11306
rect 82430 11252 82630 11264
rect 82430 11218 82442 11252
rect 82618 11218 82630 11252
rect 82430 11206 82630 11218
rect 82430 11030 82630 11042
rect 82430 10996 82442 11030
rect 82618 10996 82630 11030
rect 82430 10984 82630 10996
rect 82430 10942 82630 10954
rect 82430 10908 82442 10942
rect 82618 10908 82630 10942
rect 82430 10896 82630 10908
rect -1860 9630 -1660 9642
rect -1860 9596 -1848 9630
rect -1672 9596 -1660 9630
rect -1860 9584 -1660 9596
rect -1860 9542 -1660 9554
rect -1860 9508 -1848 9542
rect -1672 9508 -1660 9542
rect -1860 9496 -1660 9508
rect -1860 9320 -1660 9332
rect -1860 9286 -1848 9320
rect -1672 9286 -1660 9320
rect -1860 9274 -1660 9286
rect -1860 9232 -1660 9244
rect -1860 9198 -1848 9232
rect -1672 9198 -1660 9232
rect -1860 9186 -1660 9198
rect 82430 9630 82630 9642
rect 82430 9596 82442 9630
rect 82618 9596 82630 9630
rect 82430 9584 82630 9596
rect 82430 9542 82630 9554
rect 82430 9508 82442 9542
rect 82618 9508 82630 9542
rect 82430 9496 82630 9508
rect 82430 9320 82630 9332
rect 82430 9286 82442 9320
rect 82618 9286 82630 9320
rect 82430 9274 82630 9286
rect 82430 9232 82630 9244
rect 82430 9198 82442 9232
rect 82618 9198 82630 9232
rect 82430 9186 82630 9198
rect -1860 7920 -1660 7932
rect -1860 7886 -1848 7920
rect -1672 7886 -1660 7920
rect -1860 7874 -1660 7886
rect -1860 7832 -1660 7844
rect -1860 7798 -1848 7832
rect -1672 7798 -1660 7832
rect -1860 7786 -1660 7798
rect -1860 7610 -1660 7622
rect -1860 7576 -1848 7610
rect -1672 7576 -1660 7610
rect -1860 7564 -1660 7576
rect -1860 7522 -1660 7534
rect -1860 7488 -1848 7522
rect -1672 7488 -1660 7522
rect -1860 7476 -1660 7488
rect 82430 7920 82630 7932
rect 82430 7886 82442 7920
rect 82618 7886 82630 7920
rect 82430 7874 82630 7886
rect 82430 7832 82630 7844
rect 82430 7798 82442 7832
rect 82618 7798 82630 7832
rect 82430 7786 82630 7798
rect 82430 7610 82630 7622
rect 82430 7576 82442 7610
rect 82618 7576 82630 7610
rect 82430 7564 82630 7576
rect 82430 7522 82630 7534
rect 82430 7488 82442 7522
rect 82618 7488 82630 7522
rect 82430 7476 82630 7488
rect -1860 6210 -1660 6222
rect -1860 6176 -1848 6210
rect -1672 6176 -1660 6210
rect -1860 6164 -1660 6176
rect -1860 6122 -1660 6134
rect -1860 6088 -1848 6122
rect -1672 6088 -1660 6122
rect -1860 6076 -1660 6088
rect -1860 5900 -1660 5912
rect -1860 5866 -1848 5900
rect -1672 5866 -1660 5900
rect -1860 5854 -1660 5866
rect -1860 5812 -1660 5824
rect -1860 5778 -1848 5812
rect -1672 5778 -1660 5812
rect -1860 5766 -1660 5778
rect 82430 6210 82630 6222
rect 82430 6176 82442 6210
rect 82618 6176 82630 6210
rect 82430 6164 82630 6176
rect 82430 6122 82630 6134
rect 82430 6088 82442 6122
rect 82618 6088 82630 6122
rect 82430 6076 82630 6088
rect 82430 5900 82630 5912
rect 82430 5866 82442 5900
rect 82618 5866 82630 5900
rect 82430 5854 82630 5866
rect 82430 5812 82630 5824
rect 82430 5778 82442 5812
rect 82618 5778 82630 5812
rect 82430 5766 82630 5778
rect -1860 4500 -1660 4512
rect -1860 4466 -1848 4500
rect -1672 4466 -1660 4500
rect -1860 4454 -1660 4466
rect -1860 4412 -1660 4424
rect -1860 4378 -1848 4412
rect -1672 4378 -1660 4412
rect -1860 4366 -1660 4378
rect -1860 4190 -1660 4202
rect -1860 4156 -1848 4190
rect -1672 4156 -1660 4190
rect -1860 4144 -1660 4156
rect -1860 4102 -1660 4114
rect -1860 4068 -1848 4102
rect -1672 4068 -1660 4102
rect -1860 4056 -1660 4068
rect 82430 4500 82630 4512
rect 82430 4466 82442 4500
rect 82618 4466 82630 4500
rect 82430 4454 82630 4466
rect 82430 4412 82630 4424
rect 82430 4378 82442 4412
rect 82618 4378 82630 4412
rect 82430 4366 82630 4378
rect 82430 4190 82630 4202
rect 82430 4156 82442 4190
rect 82618 4156 82630 4190
rect 82430 4144 82630 4156
rect 82430 4102 82630 4114
rect 82430 4068 82442 4102
rect 82618 4068 82630 4102
rect 82430 4056 82630 4068
rect -1860 2790 -1660 2802
rect -1860 2756 -1848 2790
rect -1672 2756 -1660 2790
rect -1860 2744 -1660 2756
rect -1860 2702 -1660 2714
rect -1860 2668 -1848 2702
rect -1672 2668 -1660 2702
rect -1860 2656 -1660 2668
rect -1860 2480 -1660 2492
rect -1860 2446 -1848 2480
rect -1672 2446 -1660 2480
rect -1860 2434 -1660 2446
rect -1860 2392 -1660 2404
rect -1860 2358 -1848 2392
rect -1672 2358 -1660 2392
rect -1860 2346 -1660 2358
rect 82430 2790 82630 2802
rect 82430 2756 82442 2790
rect 82618 2756 82630 2790
rect 82430 2744 82630 2756
rect 82430 2702 82630 2714
rect 82430 2668 82442 2702
rect 82618 2668 82630 2702
rect 82430 2656 82630 2668
rect 82430 2480 82630 2492
rect 82430 2446 82442 2480
rect 82618 2446 82630 2480
rect 82430 2434 82630 2446
rect 82430 2392 82630 2404
rect 82430 2358 82442 2392
rect 82618 2358 82630 2392
rect 82430 2346 82630 2358
rect -1860 1080 -1660 1092
rect -1860 1046 -1848 1080
rect -1672 1046 -1660 1080
rect -1860 1034 -1660 1046
rect -1860 992 -1660 1004
rect -1860 958 -1848 992
rect -1672 958 -1660 992
rect -1860 946 -1660 958
rect -1860 770 -1660 782
rect -1860 736 -1848 770
rect -1672 736 -1660 770
rect -1860 724 -1660 736
rect -1860 682 -1660 694
rect -1860 648 -1848 682
rect -1672 648 -1660 682
rect -1860 636 -1660 648
rect 82430 1080 82630 1092
rect 82430 1046 82442 1080
rect 82618 1046 82630 1080
rect 82430 1034 82630 1046
rect 82430 992 82630 1004
rect 82430 958 82442 992
rect 82618 958 82630 992
rect 82430 946 82630 958
rect 82430 770 82630 782
rect 82430 736 82442 770
rect 82618 736 82630 770
rect 82430 724 82630 736
rect 82430 682 82630 694
rect 82430 648 82442 682
rect 82618 648 82630 682
rect 82430 636 82630 648
rect -1860 -630 -1660 -618
rect -1860 -664 -1848 -630
rect -1672 -664 -1660 -630
rect -1860 -676 -1660 -664
rect -1860 -718 -1660 -706
rect -1860 -752 -1848 -718
rect -1672 -752 -1660 -718
rect -1860 -764 -1660 -752
rect -1860 -940 -1660 -928
rect -1860 -974 -1848 -940
rect -1672 -974 -1660 -940
rect -1860 -986 -1660 -974
rect -1860 -1028 -1660 -1016
rect -1860 -1062 -1848 -1028
rect -1672 -1062 -1660 -1028
rect -1860 -1074 -1660 -1062
rect 2860 -630 3060 -618
rect 2860 -664 2872 -630
rect 3048 -664 3060 -630
rect 2860 -676 3060 -664
rect 2860 -718 3060 -706
rect 2860 -752 2872 -718
rect 3048 -752 3060 -718
rect 2860 -764 3060 -752
rect 2860 -940 3060 -928
rect 2860 -974 2872 -940
rect 3048 -974 3060 -940
rect 2860 -986 3060 -974
rect 2860 -1028 3060 -1016
rect 2860 -1062 2872 -1028
rect 3048 -1062 3060 -1028
rect 2860 -1074 3060 -1062
rect 7850 -630 8050 -618
rect 7850 -664 7862 -630
rect 8038 -664 8050 -630
rect 7850 -676 8050 -664
rect 7850 -718 8050 -706
rect 7850 -752 7862 -718
rect 8038 -752 8050 -718
rect 7850 -764 8050 -752
rect 7850 -940 8050 -928
rect 7850 -974 7862 -940
rect 8038 -974 8050 -940
rect 7850 -986 8050 -974
rect 7850 -1028 8050 -1016
rect 7850 -1062 7862 -1028
rect 8038 -1062 8050 -1028
rect 7850 -1074 8050 -1062
rect 12840 -630 13040 -618
rect 12840 -664 12852 -630
rect 13028 -664 13040 -630
rect 12840 -676 13040 -664
rect 12840 -718 13040 -706
rect 12840 -752 12852 -718
rect 13028 -752 13040 -718
rect 12840 -764 13040 -752
rect 12840 -940 13040 -928
rect 12840 -974 12852 -940
rect 13028 -974 13040 -940
rect 12840 -986 13040 -974
rect 12840 -1028 13040 -1016
rect 12840 -1062 12852 -1028
rect 13028 -1062 13040 -1028
rect 12840 -1074 13040 -1062
rect 17830 -630 18030 -618
rect 17830 -664 17842 -630
rect 18018 -664 18030 -630
rect 17830 -676 18030 -664
rect 17830 -718 18030 -706
rect 17830 -752 17842 -718
rect 18018 -752 18030 -718
rect 17830 -764 18030 -752
rect 17830 -940 18030 -928
rect 17830 -974 17842 -940
rect 18018 -974 18030 -940
rect 17830 -986 18030 -974
rect 17830 -1028 18030 -1016
rect 17830 -1062 17842 -1028
rect 18018 -1062 18030 -1028
rect 17830 -1074 18030 -1062
rect 22820 -630 23020 -618
rect 22820 -664 22832 -630
rect 23008 -664 23020 -630
rect 22820 -676 23020 -664
rect 22820 -718 23020 -706
rect 22820 -752 22832 -718
rect 23008 -752 23020 -718
rect 22820 -764 23020 -752
rect 22820 -940 23020 -928
rect 22820 -974 22832 -940
rect 23008 -974 23020 -940
rect 22820 -986 23020 -974
rect 22820 -1028 23020 -1016
rect 22820 -1062 22832 -1028
rect 23008 -1062 23020 -1028
rect 22820 -1074 23020 -1062
rect 27810 -630 28010 -618
rect 27810 -664 27822 -630
rect 27998 -664 28010 -630
rect 27810 -676 28010 -664
rect 27810 -718 28010 -706
rect 27810 -752 27822 -718
rect 27998 -752 28010 -718
rect 27810 -764 28010 -752
rect 27810 -940 28010 -928
rect 27810 -974 27822 -940
rect 27998 -974 28010 -940
rect 27810 -986 28010 -974
rect 27810 -1028 28010 -1016
rect 27810 -1062 27822 -1028
rect 27998 -1062 28010 -1028
rect 27810 -1074 28010 -1062
rect 32800 -630 33000 -618
rect 32800 -664 32812 -630
rect 32988 -664 33000 -630
rect 32800 -676 33000 -664
rect 32800 -718 33000 -706
rect 32800 -752 32812 -718
rect 32988 -752 33000 -718
rect 32800 -764 33000 -752
rect 32800 -940 33000 -928
rect 32800 -974 32812 -940
rect 32988 -974 33000 -940
rect 32800 -986 33000 -974
rect 32800 -1028 33000 -1016
rect 32800 -1062 32812 -1028
rect 32988 -1062 33000 -1028
rect 32800 -1074 33000 -1062
rect 37790 -630 37990 -618
rect 37790 -664 37802 -630
rect 37978 -664 37990 -630
rect 37790 -676 37990 -664
rect 37790 -718 37990 -706
rect 37790 -752 37802 -718
rect 37978 -752 37990 -718
rect 37790 -764 37990 -752
rect 37790 -940 37990 -928
rect 37790 -974 37802 -940
rect 37978 -974 37990 -940
rect 37790 -986 37990 -974
rect 37790 -1028 37990 -1016
rect 37790 -1062 37802 -1028
rect 37978 -1062 37990 -1028
rect 37790 -1074 37990 -1062
rect 42780 -630 42980 -618
rect 42780 -664 42792 -630
rect 42968 -664 42980 -630
rect 42780 -676 42980 -664
rect 42780 -718 42980 -706
rect 42780 -752 42792 -718
rect 42968 -752 42980 -718
rect 42780 -764 42980 -752
rect 42780 -940 42980 -928
rect 42780 -974 42792 -940
rect 42968 -974 42980 -940
rect 42780 -986 42980 -974
rect 42780 -1028 42980 -1016
rect 42780 -1062 42792 -1028
rect 42968 -1062 42980 -1028
rect 42780 -1074 42980 -1062
rect 47770 -630 47970 -618
rect 47770 -664 47782 -630
rect 47958 -664 47970 -630
rect 47770 -676 47970 -664
rect 47770 -718 47970 -706
rect 47770 -752 47782 -718
rect 47958 -752 47970 -718
rect 47770 -764 47970 -752
rect 47770 -940 47970 -928
rect 47770 -974 47782 -940
rect 47958 -974 47970 -940
rect 47770 -986 47970 -974
rect 47770 -1028 47970 -1016
rect 47770 -1062 47782 -1028
rect 47958 -1062 47970 -1028
rect 47770 -1074 47970 -1062
rect 52760 -630 52960 -618
rect 52760 -664 52772 -630
rect 52948 -664 52960 -630
rect 52760 -676 52960 -664
rect 52760 -718 52960 -706
rect 52760 -752 52772 -718
rect 52948 -752 52960 -718
rect 52760 -764 52960 -752
rect 52760 -940 52960 -928
rect 52760 -974 52772 -940
rect 52948 -974 52960 -940
rect 52760 -986 52960 -974
rect 52760 -1028 52960 -1016
rect 52760 -1062 52772 -1028
rect 52948 -1062 52960 -1028
rect 52760 -1074 52960 -1062
rect 57750 -630 57950 -618
rect 57750 -664 57762 -630
rect 57938 -664 57950 -630
rect 57750 -676 57950 -664
rect 57750 -718 57950 -706
rect 57750 -752 57762 -718
rect 57938 -752 57950 -718
rect 57750 -764 57950 -752
rect 57750 -940 57950 -928
rect 57750 -974 57762 -940
rect 57938 -974 57950 -940
rect 57750 -986 57950 -974
rect 57750 -1028 57950 -1016
rect 57750 -1062 57762 -1028
rect 57938 -1062 57950 -1028
rect 57750 -1074 57950 -1062
rect 62740 -630 62940 -618
rect 62740 -664 62752 -630
rect 62928 -664 62940 -630
rect 62740 -676 62940 -664
rect 62740 -718 62940 -706
rect 62740 -752 62752 -718
rect 62928 -752 62940 -718
rect 62740 -764 62940 -752
rect 62740 -940 62940 -928
rect 62740 -974 62752 -940
rect 62928 -974 62940 -940
rect 62740 -986 62940 -974
rect 62740 -1028 62940 -1016
rect 62740 -1062 62752 -1028
rect 62928 -1062 62940 -1028
rect 62740 -1074 62940 -1062
rect 67730 -630 67930 -618
rect 67730 -664 67742 -630
rect 67918 -664 67930 -630
rect 67730 -676 67930 -664
rect 67730 -718 67930 -706
rect 67730 -752 67742 -718
rect 67918 -752 67930 -718
rect 67730 -764 67930 -752
rect 67730 -940 67930 -928
rect 67730 -974 67742 -940
rect 67918 -974 67930 -940
rect 67730 -986 67930 -974
rect 67730 -1028 67930 -1016
rect 67730 -1062 67742 -1028
rect 67918 -1062 67930 -1028
rect 67730 -1074 67930 -1062
rect 72720 -630 72920 -618
rect 72720 -664 72732 -630
rect 72908 -664 72920 -630
rect 72720 -676 72920 -664
rect 72720 -718 72920 -706
rect 72720 -752 72732 -718
rect 72908 -752 72920 -718
rect 72720 -764 72920 -752
rect 72720 -940 72920 -928
rect 72720 -974 72732 -940
rect 72908 -974 72920 -940
rect 72720 -986 72920 -974
rect 72720 -1028 72920 -1016
rect 72720 -1062 72732 -1028
rect 72908 -1062 72920 -1028
rect 72720 -1074 72920 -1062
rect 77710 -630 77910 -618
rect 77710 -664 77722 -630
rect 77898 -664 77910 -630
rect 77710 -676 77910 -664
rect 77710 -718 77910 -706
rect 77710 -752 77722 -718
rect 77898 -752 77910 -718
rect 77710 -764 77910 -752
rect 77710 -940 77910 -928
rect 77710 -974 77722 -940
rect 77898 -974 77910 -940
rect 77710 -986 77910 -974
rect 77710 -1028 77910 -1016
rect 77710 -1062 77722 -1028
rect 77898 -1062 77910 -1028
rect 77710 -1074 77910 -1062
rect 82430 -630 82630 -618
rect 82430 -664 82442 -630
rect 82618 -664 82630 -630
rect 82430 -676 82630 -664
rect 82430 -718 82630 -706
rect 82430 -752 82442 -718
rect 82618 -752 82630 -718
rect 82430 -764 82630 -752
rect 82430 -940 82630 -928
rect 82430 -974 82442 -940
rect 82618 -974 82630 -940
rect 82430 -986 82630 -974
rect 82430 -1028 82630 -1016
rect 82430 -1062 82442 -1028
rect 82618 -1062 82630 -1028
rect 82430 -1074 82630 -1062
<< pdiff >>
rect 3358 28440 3558 28452
rect 3358 28406 3370 28440
rect 3546 28406 3558 28440
rect 3358 28394 3558 28406
rect 3358 28352 3558 28364
rect 3358 28318 3370 28352
rect 3546 28318 3558 28352
rect 3358 28306 3558 28318
rect 3358 28130 3558 28142
rect 3358 28096 3370 28130
rect 3546 28096 3558 28130
rect 3358 28084 3558 28096
rect 3358 28042 3558 28054
rect 3358 28008 3370 28042
rect 3546 28008 3558 28042
rect 3358 27996 3558 28008
rect 8348 28440 8548 28452
rect 8348 28406 8360 28440
rect 8536 28406 8548 28440
rect 8348 28394 8548 28406
rect 8348 28352 8548 28364
rect 8348 28318 8360 28352
rect 8536 28318 8548 28352
rect 8348 28306 8548 28318
rect 8348 28130 8548 28142
rect 8348 28096 8360 28130
rect 8536 28096 8548 28130
rect 8348 28084 8548 28096
rect 8348 28042 8548 28054
rect 8348 28008 8360 28042
rect 8536 28008 8548 28042
rect 8348 27996 8548 28008
rect 13338 28440 13538 28452
rect 13338 28406 13350 28440
rect 13526 28406 13538 28440
rect 13338 28394 13538 28406
rect 13338 28352 13538 28364
rect 13338 28318 13350 28352
rect 13526 28318 13538 28352
rect 13338 28306 13538 28318
rect 13338 28130 13538 28142
rect 13338 28096 13350 28130
rect 13526 28096 13538 28130
rect 13338 28084 13538 28096
rect 13338 28042 13538 28054
rect 13338 28008 13350 28042
rect 13526 28008 13538 28042
rect 13338 27996 13538 28008
rect 18328 28440 18528 28452
rect 18328 28406 18340 28440
rect 18516 28406 18528 28440
rect 18328 28394 18528 28406
rect 18328 28352 18528 28364
rect 18328 28318 18340 28352
rect 18516 28318 18528 28352
rect 18328 28306 18528 28318
rect 18328 28130 18528 28142
rect 18328 28096 18340 28130
rect 18516 28096 18528 28130
rect 18328 28084 18528 28096
rect 18328 28042 18528 28054
rect 18328 28008 18340 28042
rect 18516 28008 18528 28042
rect 18328 27996 18528 28008
rect 23318 28440 23518 28452
rect 23318 28406 23330 28440
rect 23506 28406 23518 28440
rect 23318 28394 23518 28406
rect 23318 28352 23518 28364
rect 23318 28318 23330 28352
rect 23506 28318 23518 28352
rect 23318 28306 23518 28318
rect 23318 28130 23518 28142
rect 23318 28096 23330 28130
rect 23506 28096 23518 28130
rect 23318 28084 23518 28096
rect 23318 28042 23518 28054
rect 23318 28008 23330 28042
rect 23506 28008 23518 28042
rect 23318 27996 23518 28008
rect 28308 28440 28508 28452
rect 28308 28406 28320 28440
rect 28496 28406 28508 28440
rect 28308 28394 28508 28406
rect 28308 28352 28508 28364
rect 28308 28318 28320 28352
rect 28496 28318 28508 28352
rect 28308 28306 28508 28318
rect 28308 28130 28508 28142
rect 28308 28096 28320 28130
rect 28496 28096 28508 28130
rect 28308 28084 28508 28096
rect 28308 28042 28508 28054
rect 28308 28008 28320 28042
rect 28496 28008 28508 28042
rect 28308 27996 28508 28008
rect 33298 28440 33498 28452
rect 33298 28406 33310 28440
rect 33486 28406 33498 28440
rect 33298 28394 33498 28406
rect 33298 28352 33498 28364
rect 33298 28318 33310 28352
rect 33486 28318 33498 28352
rect 33298 28306 33498 28318
rect 33298 28130 33498 28142
rect 33298 28096 33310 28130
rect 33486 28096 33498 28130
rect 33298 28084 33498 28096
rect 33298 28042 33498 28054
rect 33298 28008 33310 28042
rect 33486 28008 33498 28042
rect 33298 27996 33498 28008
rect 38288 28440 38488 28452
rect 38288 28406 38300 28440
rect 38476 28406 38488 28440
rect 38288 28394 38488 28406
rect 38288 28352 38488 28364
rect 38288 28318 38300 28352
rect 38476 28318 38488 28352
rect 38288 28306 38488 28318
rect 38288 28130 38488 28142
rect 38288 28096 38300 28130
rect 38476 28096 38488 28130
rect 38288 28084 38488 28096
rect 38288 28042 38488 28054
rect 38288 28008 38300 28042
rect 38476 28008 38488 28042
rect 38288 27996 38488 28008
rect 43278 28440 43478 28452
rect 43278 28406 43290 28440
rect 43466 28406 43478 28440
rect 43278 28394 43478 28406
rect 43278 28352 43478 28364
rect 43278 28318 43290 28352
rect 43466 28318 43478 28352
rect 43278 28306 43478 28318
rect 43278 28130 43478 28142
rect 43278 28096 43290 28130
rect 43466 28096 43478 28130
rect 43278 28084 43478 28096
rect 43278 28042 43478 28054
rect 43278 28008 43290 28042
rect 43466 28008 43478 28042
rect 43278 27996 43478 28008
rect 48268 28440 48468 28452
rect 48268 28406 48280 28440
rect 48456 28406 48468 28440
rect 48268 28394 48468 28406
rect 48268 28352 48468 28364
rect 48268 28318 48280 28352
rect 48456 28318 48468 28352
rect 48268 28306 48468 28318
rect 48268 28130 48468 28142
rect 48268 28096 48280 28130
rect 48456 28096 48468 28130
rect 48268 28084 48468 28096
rect 48268 28042 48468 28054
rect 48268 28008 48280 28042
rect 48456 28008 48468 28042
rect 48268 27996 48468 28008
rect 53258 28440 53458 28452
rect 53258 28406 53270 28440
rect 53446 28406 53458 28440
rect 53258 28394 53458 28406
rect 53258 28352 53458 28364
rect 53258 28318 53270 28352
rect 53446 28318 53458 28352
rect 53258 28306 53458 28318
rect 53258 28130 53458 28142
rect 53258 28096 53270 28130
rect 53446 28096 53458 28130
rect 53258 28084 53458 28096
rect 53258 28042 53458 28054
rect 53258 28008 53270 28042
rect 53446 28008 53458 28042
rect 53258 27996 53458 28008
rect 58248 28440 58448 28452
rect 58248 28406 58260 28440
rect 58436 28406 58448 28440
rect 58248 28394 58448 28406
rect 58248 28352 58448 28364
rect 58248 28318 58260 28352
rect 58436 28318 58448 28352
rect 58248 28306 58448 28318
rect 58248 28130 58448 28142
rect 58248 28096 58260 28130
rect 58436 28096 58448 28130
rect 58248 28084 58448 28096
rect 58248 28042 58448 28054
rect 58248 28008 58260 28042
rect 58436 28008 58448 28042
rect 58248 27996 58448 28008
rect 63238 28440 63438 28452
rect 63238 28406 63250 28440
rect 63426 28406 63438 28440
rect 63238 28394 63438 28406
rect 63238 28352 63438 28364
rect 63238 28318 63250 28352
rect 63426 28318 63438 28352
rect 63238 28306 63438 28318
rect 63238 28130 63438 28142
rect 63238 28096 63250 28130
rect 63426 28096 63438 28130
rect 63238 28084 63438 28096
rect 63238 28042 63438 28054
rect 63238 28008 63250 28042
rect 63426 28008 63438 28042
rect 63238 27996 63438 28008
rect 68228 28440 68428 28452
rect 68228 28406 68240 28440
rect 68416 28406 68428 28440
rect 68228 28394 68428 28406
rect 68228 28352 68428 28364
rect 68228 28318 68240 28352
rect 68416 28318 68428 28352
rect 68228 28306 68428 28318
rect 68228 28130 68428 28142
rect 68228 28096 68240 28130
rect 68416 28096 68428 28130
rect 68228 28084 68428 28096
rect 68228 28042 68428 28054
rect 68228 28008 68240 28042
rect 68416 28008 68428 28042
rect 68228 27996 68428 28008
rect 73218 28440 73418 28452
rect 73218 28406 73230 28440
rect 73406 28406 73418 28440
rect 73218 28394 73418 28406
rect 73218 28352 73418 28364
rect 73218 28318 73230 28352
rect 73406 28318 73418 28352
rect 73218 28306 73418 28318
rect 73218 28130 73418 28142
rect 73218 28096 73230 28130
rect 73406 28096 73418 28130
rect 73218 28084 73418 28096
rect 73218 28042 73418 28054
rect 73218 28008 73230 28042
rect 73406 28008 73418 28042
rect 73218 27996 73418 28008
rect 78208 28440 78408 28452
rect 78208 28406 78220 28440
rect 78396 28406 78408 28440
rect 78208 28394 78408 28406
rect 78208 28352 78408 28364
rect 78208 28318 78220 28352
rect 78396 28318 78408 28352
rect 78208 28306 78408 28318
rect 78208 28130 78408 28142
rect 78208 28096 78220 28130
rect 78396 28096 78408 28130
rect 78208 28084 78408 28096
rect 78208 28042 78408 28054
rect 78208 28008 78220 28042
rect 78396 28008 78408 28042
rect 78208 27996 78408 28008
rect 82928 28440 83128 28452
rect 82928 28406 82940 28440
rect 83116 28406 83128 28440
rect 82928 28394 83128 28406
rect 82928 28352 83128 28364
rect 82928 28318 82940 28352
rect 83116 28318 83128 28352
rect 82928 28306 83128 28318
rect 82928 28130 83128 28142
rect 82928 28096 82940 28130
rect 83116 28096 83128 28130
rect 82928 28084 83128 28096
rect 82928 28042 83128 28054
rect 82928 28008 82940 28042
rect 83116 28008 83128 28042
rect 82928 27996 83128 28008
rect 82928 26730 83128 26742
rect 82928 26696 82940 26730
rect 83116 26696 83128 26730
rect 82928 26684 83128 26696
rect 82928 26642 83128 26654
rect 82928 26608 82940 26642
rect 83116 26608 83128 26642
rect 82928 26596 83128 26608
rect 82928 26420 83128 26432
rect 82928 26386 82940 26420
rect 83116 26386 83128 26420
rect 82928 26374 83128 26386
rect 82928 26332 83128 26344
rect 82928 26298 82940 26332
rect 83116 26298 83128 26332
rect 82928 26286 83128 26298
rect 82928 25020 83128 25032
rect 82928 24986 82940 25020
rect 83116 24986 83128 25020
rect 82928 24974 83128 24986
rect 82928 24932 83128 24944
rect 82928 24898 82940 24932
rect 83116 24898 83128 24932
rect 82928 24886 83128 24898
rect 82928 24710 83128 24722
rect 82928 24676 82940 24710
rect 83116 24676 83128 24710
rect 82928 24664 83128 24676
rect 82928 24622 83128 24634
rect 82928 24588 82940 24622
rect 83116 24588 83128 24622
rect 82928 24576 83128 24588
rect -1362 23310 -1162 23322
rect -1362 23276 -1350 23310
rect -1174 23276 -1162 23310
rect -1362 23264 -1162 23276
rect -1362 23222 -1162 23234
rect -1362 23188 -1350 23222
rect -1174 23188 -1162 23222
rect -1362 23176 -1162 23188
rect -1362 23000 -1162 23012
rect -1362 22966 -1350 23000
rect -1174 22966 -1162 23000
rect -1362 22954 -1162 22966
rect -1362 22912 -1162 22924
rect -1362 22878 -1350 22912
rect -1174 22878 -1162 22912
rect -1362 22866 -1162 22878
rect 82928 23310 83128 23322
rect 82928 23276 82940 23310
rect 83116 23276 83128 23310
rect 82928 23264 83128 23276
rect 82928 23222 83128 23234
rect 82928 23188 82940 23222
rect 83116 23188 83128 23222
rect 82928 23176 83128 23188
rect 82928 23000 83128 23012
rect 82928 22966 82940 23000
rect 83116 22966 83128 23000
rect 82928 22954 83128 22966
rect 82928 22912 83128 22924
rect 82928 22878 82940 22912
rect 83116 22878 83128 22912
rect 82928 22866 83128 22878
rect -1362 21600 -1162 21612
rect -1362 21566 -1350 21600
rect -1174 21566 -1162 21600
rect -1362 21554 -1162 21566
rect -1362 21512 -1162 21524
rect -1362 21478 -1350 21512
rect -1174 21478 -1162 21512
rect -1362 21466 -1162 21478
rect -1362 21290 -1162 21302
rect -1362 21256 -1350 21290
rect -1174 21256 -1162 21290
rect -1362 21244 -1162 21256
rect -1362 21202 -1162 21214
rect -1362 21168 -1350 21202
rect -1174 21168 -1162 21202
rect -1362 21156 -1162 21168
rect 82928 21600 83128 21612
rect 82928 21566 82940 21600
rect 83116 21566 83128 21600
rect 82928 21554 83128 21566
rect 82928 21512 83128 21524
rect 82928 21478 82940 21512
rect 83116 21478 83128 21512
rect 82928 21466 83128 21478
rect 82928 21290 83128 21302
rect 82928 21256 82940 21290
rect 83116 21256 83128 21290
rect 82928 21244 83128 21256
rect 82928 21202 83128 21214
rect 82928 21168 82940 21202
rect 83116 21168 83128 21202
rect 82928 21156 83128 21168
rect -1362 19890 -1162 19902
rect -1362 19856 -1350 19890
rect -1174 19856 -1162 19890
rect -1362 19844 -1162 19856
rect -1362 19802 -1162 19814
rect -1362 19768 -1350 19802
rect -1174 19768 -1162 19802
rect -1362 19756 -1162 19768
rect -1362 19580 -1162 19592
rect -1362 19546 -1350 19580
rect -1174 19546 -1162 19580
rect -1362 19534 -1162 19546
rect -1362 19492 -1162 19504
rect -1362 19458 -1350 19492
rect -1174 19458 -1162 19492
rect -1362 19446 -1162 19458
rect 82928 19890 83128 19902
rect 82928 19856 82940 19890
rect 83116 19856 83128 19890
rect 82928 19844 83128 19856
rect 82928 19802 83128 19814
rect 82928 19768 82940 19802
rect 83116 19768 83128 19802
rect 82928 19756 83128 19768
rect 82928 19580 83128 19592
rect 82928 19546 82940 19580
rect 83116 19546 83128 19580
rect 82928 19534 83128 19546
rect 82928 19492 83128 19504
rect 82928 19458 82940 19492
rect 83116 19458 83128 19492
rect 82928 19446 83128 19458
rect -1362 18180 -1162 18192
rect -1362 18146 -1350 18180
rect -1174 18146 -1162 18180
rect -1362 18134 -1162 18146
rect -1362 18092 -1162 18104
rect -1362 18058 -1350 18092
rect -1174 18058 -1162 18092
rect -1362 18046 -1162 18058
rect -1362 17870 -1162 17882
rect -1362 17836 -1350 17870
rect -1174 17836 -1162 17870
rect -1362 17824 -1162 17836
rect -1362 17782 -1162 17794
rect -1362 17748 -1350 17782
rect -1174 17748 -1162 17782
rect -1362 17736 -1162 17748
rect 82928 18180 83128 18192
rect 82928 18146 82940 18180
rect 83116 18146 83128 18180
rect 82928 18134 83128 18146
rect 82928 18092 83128 18104
rect 82928 18058 82940 18092
rect 83116 18058 83128 18092
rect 82928 18046 83128 18058
rect 82928 17870 83128 17882
rect 82928 17836 82940 17870
rect 83116 17836 83128 17870
rect 82928 17824 83128 17836
rect 82928 17782 83128 17794
rect 82928 17748 82940 17782
rect 83116 17748 83128 17782
rect 82928 17736 83128 17748
rect -1362 16470 -1162 16482
rect -1362 16436 -1350 16470
rect -1174 16436 -1162 16470
rect -1362 16424 -1162 16436
rect -1362 16382 -1162 16394
rect -1362 16348 -1350 16382
rect -1174 16348 -1162 16382
rect -1362 16336 -1162 16348
rect -1362 16160 -1162 16172
rect -1362 16126 -1350 16160
rect -1174 16126 -1162 16160
rect -1362 16114 -1162 16126
rect -1362 16072 -1162 16084
rect -1362 16038 -1350 16072
rect -1174 16038 -1162 16072
rect -1362 16026 -1162 16038
rect 82928 16470 83128 16482
rect 82928 16436 82940 16470
rect 83116 16436 83128 16470
rect 82928 16424 83128 16436
rect 82928 16382 83128 16394
rect 82928 16348 82940 16382
rect 83116 16348 83128 16382
rect 82928 16336 83128 16348
rect 82928 16160 83128 16172
rect 82928 16126 82940 16160
rect 83116 16126 83128 16160
rect 82928 16114 83128 16126
rect 82928 16072 83128 16084
rect 82928 16038 82940 16072
rect 83116 16038 83128 16072
rect 82928 16026 83128 16038
rect -1362 14760 -1162 14772
rect -1362 14726 -1350 14760
rect -1174 14726 -1162 14760
rect -1362 14714 -1162 14726
rect -1362 14672 -1162 14684
rect -1362 14638 -1350 14672
rect -1174 14638 -1162 14672
rect -1362 14626 -1162 14638
rect -1362 14450 -1162 14462
rect -1362 14416 -1350 14450
rect -1174 14416 -1162 14450
rect -1362 14404 -1162 14416
rect -1362 14362 -1162 14374
rect -1362 14328 -1350 14362
rect -1174 14328 -1162 14362
rect -1362 14316 -1162 14328
rect 82928 14760 83128 14772
rect 82928 14726 82940 14760
rect 83116 14726 83128 14760
rect 82928 14714 83128 14726
rect 82928 14672 83128 14684
rect 82928 14638 82940 14672
rect 83116 14638 83128 14672
rect 82928 14626 83128 14638
rect 82928 14450 83128 14462
rect 82928 14416 82940 14450
rect 83116 14416 83128 14450
rect 82928 14404 83128 14416
rect 82928 14362 83128 14374
rect 82928 14328 82940 14362
rect 83116 14328 83128 14362
rect 82928 14316 83128 14328
rect -1362 13050 -1162 13062
rect -1362 13016 -1350 13050
rect -1174 13016 -1162 13050
rect -1362 13004 -1162 13016
rect -1362 12962 -1162 12974
rect -1362 12928 -1350 12962
rect -1174 12928 -1162 12962
rect -1362 12916 -1162 12928
rect -1362 12740 -1162 12752
rect -1362 12706 -1350 12740
rect -1174 12706 -1162 12740
rect -1362 12694 -1162 12706
rect -1362 12652 -1162 12664
rect -1362 12618 -1350 12652
rect -1174 12618 -1162 12652
rect -1362 12606 -1162 12618
rect 82928 13050 83128 13062
rect 82928 13016 82940 13050
rect 83116 13016 83128 13050
rect 82928 13004 83128 13016
rect 82928 12962 83128 12974
rect 82928 12928 82940 12962
rect 83116 12928 83128 12962
rect 82928 12916 83128 12928
rect 82928 12740 83128 12752
rect 82928 12706 82940 12740
rect 83116 12706 83128 12740
rect 82928 12694 83128 12706
rect 82928 12652 83128 12664
rect 82928 12618 82940 12652
rect 83116 12618 83128 12652
rect 82928 12606 83128 12618
rect -1362 11340 -1162 11352
rect -1362 11306 -1350 11340
rect -1174 11306 -1162 11340
rect -1362 11294 -1162 11306
rect -1362 11252 -1162 11264
rect -1362 11218 -1350 11252
rect -1174 11218 -1162 11252
rect -1362 11206 -1162 11218
rect -1362 11030 -1162 11042
rect -1362 10996 -1350 11030
rect -1174 10996 -1162 11030
rect -1362 10984 -1162 10996
rect -1362 10942 -1162 10954
rect -1362 10908 -1350 10942
rect -1174 10908 -1162 10942
rect -1362 10896 -1162 10908
rect 82928 11340 83128 11352
rect 82928 11306 82940 11340
rect 83116 11306 83128 11340
rect 82928 11294 83128 11306
rect 82928 11252 83128 11264
rect 82928 11218 82940 11252
rect 83116 11218 83128 11252
rect 82928 11206 83128 11218
rect 82928 11030 83128 11042
rect 82928 10996 82940 11030
rect 83116 10996 83128 11030
rect 82928 10984 83128 10996
rect 82928 10942 83128 10954
rect 82928 10908 82940 10942
rect 83116 10908 83128 10942
rect 82928 10896 83128 10908
rect -1362 9630 -1162 9642
rect -1362 9596 -1350 9630
rect -1174 9596 -1162 9630
rect -1362 9584 -1162 9596
rect -1362 9542 -1162 9554
rect -1362 9508 -1350 9542
rect -1174 9508 -1162 9542
rect -1362 9496 -1162 9508
rect -1362 9320 -1162 9332
rect -1362 9286 -1350 9320
rect -1174 9286 -1162 9320
rect -1362 9274 -1162 9286
rect -1362 9232 -1162 9244
rect -1362 9198 -1350 9232
rect -1174 9198 -1162 9232
rect -1362 9186 -1162 9198
rect 82928 9630 83128 9642
rect 82928 9596 82940 9630
rect 83116 9596 83128 9630
rect 82928 9584 83128 9596
rect 82928 9542 83128 9554
rect 82928 9508 82940 9542
rect 83116 9508 83128 9542
rect 82928 9496 83128 9508
rect 82928 9320 83128 9332
rect 82928 9286 82940 9320
rect 83116 9286 83128 9320
rect 82928 9274 83128 9286
rect 82928 9232 83128 9244
rect 82928 9198 82940 9232
rect 83116 9198 83128 9232
rect 82928 9186 83128 9198
rect -1362 7920 -1162 7932
rect -1362 7886 -1350 7920
rect -1174 7886 -1162 7920
rect -1362 7874 -1162 7886
rect -1362 7832 -1162 7844
rect -1362 7798 -1350 7832
rect -1174 7798 -1162 7832
rect -1362 7786 -1162 7798
rect -1362 7610 -1162 7622
rect -1362 7576 -1350 7610
rect -1174 7576 -1162 7610
rect -1362 7564 -1162 7576
rect -1362 7522 -1162 7534
rect -1362 7488 -1350 7522
rect -1174 7488 -1162 7522
rect -1362 7476 -1162 7488
rect 82928 7920 83128 7932
rect 82928 7886 82940 7920
rect 83116 7886 83128 7920
rect 82928 7874 83128 7886
rect 82928 7832 83128 7844
rect 82928 7798 82940 7832
rect 83116 7798 83128 7832
rect 82928 7786 83128 7798
rect 82928 7610 83128 7622
rect 82928 7576 82940 7610
rect 83116 7576 83128 7610
rect 82928 7564 83128 7576
rect 82928 7522 83128 7534
rect 82928 7488 82940 7522
rect 83116 7488 83128 7522
rect 82928 7476 83128 7488
rect -1362 6210 -1162 6222
rect -1362 6176 -1350 6210
rect -1174 6176 -1162 6210
rect -1362 6164 -1162 6176
rect -1362 6122 -1162 6134
rect -1362 6088 -1350 6122
rect -1174 6088 -1162 6122
rect -1362 6076 -1162 6088
rect -1362 5900 -1162 5912
rect -1362 5866 -1350 5900
rect -1174 5866 -1162 5900
rect -1362 5854 -1162 5866
rect -1362 5812 -1162 5824
rect -1362 5778 -1350 5812
rect -1174 5778 -1162 5812
rect -1362 5766 -1162 5778
rect 82928 6210 83128 6222
rect 82928 6176 82940 6210
rect 83116 6176 83128 6210
rect 82928 6164 83128 6176
rect 82928 6122 83128 6134
rect 82928 6088 82940 6122
rect 83116 6088 83128 6122
rect 82928 6076 83128 6088
rect 82928 5900 83128 5912
rect 82928 5866 82940 5900
rect 83116 5866 83128 5900
rect 82928 5854 83128 5866
rect 82928 5812 83128 5824
rect 82928 5778 82940 5812
rect 83116 5778 83128 5812
rect 82928 5766 83128 5778
rect -1362 4500 -1162 4512
rect -1362 4466 -1350 4500
rect -1174 4466 -1162 4500
rect -1362 4454 -1162 4466
rect -1362 4412 -1162 4424
rect -1362 4378 -1350 4412
rect -1174 4378 -1162 4412
rect -1362 4366 -1162 4378
rect -1362 4190 -1162 4202
rect -1362 4156 -1350 4190
rect -1174 4156 -1162 4190
rect -1362 4144 -1162 4156
rect -1362 4102 -1162 4114
rect -1362 4068 -1350 4102
rect -1174 4068 -1162 4102
rect -1362 4056 -1162 4068
rect 82928 4500 83128 4512
rect 82928 4466 82940 4500
rect 83116 4466 83128 4500
rect 82928 4454 83128 4466
rect 82928 4412 83128 4424
rect 82928 4378 82940 4412
rect 83116 4378 83128 4412
rect 82928 4366 83128 4378
rect 82928 4190 83128 4202
rect 82928 4156 82940 4190
rect 83116 4156 83128 4190
rect 82928 4144 83128 4156
rect 82928 4102 83128 4114
rect 82928 4068 82940 4102
rect 83116 4068 83128 4102
rect 82928 4056 83128 4068
rect -1362 2790 -1162 2802
rect -1362 2756 -1350 2790
rect -1174 2756 -1162 2790
rect -1362 2744 -1162 2756
rect -1362 2702 -1162 2714
rect -1362 2668 -1350 2702
rect -1174 2668 -1162 2702
rect -1362 2656 -1162 2668
rect -1362 2480 -1162 2492
rect -1362 2446 -1350 2480
rect -1174 2446 -1162 2480
rect -1362 2434 -1162 2446
rect -1362 2392 -1162 2404
rect -1362 2358 -1350 2392
rect -1174 2358 -1162 2392
rect -1362 2346 -1162 2358
rect 82928 2790 83128 2802
rect 82928 2756 82940 2790
rect 83116 2756 83128 2790
rect 82928 2744 83128 2756
rect 82928 2702 83128 2714
rect 82928 2668 82940 2702
rect 83116 2668 83128 2702
rect 82928 2656 83128 2668
rect 82928 2480 83128 2492
rect 82928 2446 82940 2480
rect 83116 2446 83128 2480
rect 82928 2434 83128 2446
rect 82928 2392 83128 2404
rect 82928 2358 82940 2392
rect 83116 2358 83128 2392
rect 82928 2346 83128 2358
rect -1362 1080 -1162 1092
rect -1362 1046 -1350 1080
rect -1174 1046 -1162 1080
rect -1362 1034 -1162 1046
rect -1362 992 -1162 1004
rect -1362 958 -1350 992
rect -1174 958 -1162 992
rect -1362 946 -1162 958
rect -1362 770 -1162 782
rect -1362 736 -1350 770
rect -1174 736 -1162 770
rect -1362 724 -1162 736
rect -1362 682 -1162 694
rect -1362 648 -1350 682
rect -1174 648 -1162 682
rect -1362 636 -1162 648
rect 82928 1080 83128 1092
rect 82928 1046 82940 1080
rect 83116 1046 83128 1080
rect 82928 1034 83128 1046
rect 82928 992 83128 1004
rect 82928 958 82940 992
rect 83116 958 83128 992
rect 82928 946 83128 958
rect 82928 770 83128 782
rect 82928 736 82940 770
rect 83116 736 83128 770
rect 82928 724 83128 736
rect 82928 682 83128 694
rect 82928 648 82940 682
rect 83116 648 83128 682
rect 82928 636 83128 648
rect -1362 -630 -1162 -618
rect -1362 -664 -1350 -630
rect -1174 -664 -1162 -630
rect -1362 -676 -1162 -664
rect -1362 -718 -1162 -706
rect -1362 -752 -1350 -718
rect -1174 -752 -1162 -718
rect -1362 -764 -1162 -752
rect -1362 -940 -1162 -928
rect -1362 -974 -1350 -940
rect -1174 -974 -1162 -940
rect -1362 -986 -1162 -974
rect -1362 -1028 -1162 -1016
rect -1362 -1062 -1350 -1028
rect -1174 -1062 -1162 -1028
rect -1362 -1074 -1162 -1062
rect 3358 -630 3558 -618
rect 3358 -664 3370 -630
rect 3546 -664 3558 -630
rect 3358 -676 3558 -664
rect 3358 -718 3558 -706
rect 3358 -752 3370 -718
rect 3546 -752 3558 -718
rect 3358 -764 3558 -752
rect 3358 -940 3558 -928
rect 3358 -974 3370 -940
rect 3546 -974 3558 -940
rect 3358 -986 3558 -974
rect 3358 -1028 3558 -1016
rect 3358 -1062 3370 -1028
rect 3546 -1062 3558 -1028
rect 3358 -1074 3558 -1062
rect 8348 -630 8548 -618
rect 8348 -664 8360 -630
rect 8536 -664 8548 -630
rect 8348 -676 8548 -664
rect 8348 -718 8548 -706
rect 8348 -752 8360 -718
rect 8536 -752 8548 -718
rect 8348 -764 8548 -752
rect 8348 -940 8548 -928
rect 8348 -974 8360 -940
rect 8536 -974 8548 -940
rect 8348 -986 8548 -974
rect 8348 -1028 8548 -1016
rect 8348 -1062 8360 -1028
rect 8536 -1062 8548 -1028
rect 8348 -1074 8548 -1062
rect 13338 -630 13538 -618
rect 13338 -664 13350 -630
rect 13526 -664 13538 -630
rect 13338 -676 13538 -664
rect 13338 -718 13538 -706
rect 13338 -752 13350 -718
rect 13526 -752 13538 -718
rect 13338 -764 13538 -752
rect 13338 -940 13538 -928
rect 13338 -974 13350 -940
rect 13526 -974 13538 -940
rect 13338 -986 13538 -974
rect 13338 -1028 13538 -1016
rect 13338 -1062 13350 -1028
rect 13526 -1062 13538 -1028
rect 13338 -1074 13538 -1062
rect 18328 -630 18528 -618
rect 18328 -664 18340 -630
rect 18516 -664 18528 -630
rect 18328 -676 18528 -664
rect 18328 -718 18528 -706
rect 18328 -752 18340 -718
rect 18516 -752 18528 -718
rect 18328 -764 18528 -752
rect 18328 -940 18528 -928
rect 18328 -974 18340 -940
rect 18516 -974 18528 -940
rect 18328 -986 18528 -974
rect 18328 -1028 18528 -1016
rect 18328 -1062 18340 -1028
rect 18516 -1062 18528 -1028
rect 18328 -1074 18528 -1062
rect 23318 -630 23518 -618
rect 23318 -664 23330 -630
rect 23506 -664 23518 -630
rect 23318 -676 23518 -664
rect 23318 -718 23518 -706
rect 23318 -752 23330 -718
rect 23506 -752 23518 -718
rect 23318 -764 23518 -752
rect 23318 -940 23518 -928
rect 23318 -974 23330 -940
rect 23506 -974 23518 -940
rect 23318 -986 23518 -974
rect 23318 -1028 23518 -1016
rect 23318 -1062 23330 -1028
rect 23506 -1062 23518 -1028
rect 23318 -1074 23518 -1062
rect 28308 -630 28508 -618
rect 28308 -664 28320 -630
rect 28496 -664 28508 -630
rect 28308 -676 28508 -664
rect 28308 -718 28508 -706
rect 28308 -752 28320 -718
rect 28496 -752 28508 -718
rect 28308 -764 28508 -752
rect 28308 -940 28508 -928
rect 28308 -974 28320 -940
rect 28496 -974 28508 -940
rect 28308 -986 28508 -974
rect 28308 -1028 28508 -1016
rect 28308 -1062 28320 -1028
rect 28496 -1062 28508 -1028
rect 28308 -1074 28508 -1062
rect 33298 -630 33498 -618
rect 33298 -664 33310 -630
rect 33486 -664 33498 -630
rect 33298 -676 33498 -664
rect 33298 -718 33498 -706
rect 33298 -752 33310 -718
rect 33486 -752 33498 -718
rect 33298 -764 33498 -752
rect 33298 -940 33498 -928
rect 33298 -974 33310 -940
rect 33486 -974 33498 -940
rect 33298 -986 33498 -974
rect 33298 -1028 33498 -1016
rect 33298 -1062 33310 -1028
rect 33486 -1062 33498 -1028
rect 33298 -1074 33498 -1062
rect 38288 -630 38488 -618
rect 38288 -664 38300 -630
rect 38476 -664 38488 -630
rect 38288 -676 38488 -664
rect 38288 -718 38488 -706
rect 38288 -752 38300 -718
rect 38476 -752 38488 -718
rect 38288 -764 38488 -752
rect 38288 -940 38488 -928
rect 38288 -974 38300 -940
rect 38476 -974 38488 -940
rect 38288 -986 38488 -974
rect 38288 -1028 38488 -1016
rect 38288 -1062 38300 -1028
rect 38476 -1062 38488 -1028
rect 38288 -1074 38488 -1062
rect 43278 -630 43478 -618
rect 43278 -664 43290 -630
rect 43466 -664 43478 -630
rect 43278 -676 43478 -664
rect 43278 -718 43478 -706
rect 43278 -752 43290 -718
rect 43466 -752 43478 -718
rect 43278 -764 43478 -752
rect 43278 -940 43478 -928
rect 43278 -974 43290 -940
rect 43466 -974 43478 -940
rect 43278 -986 43478 -974
rect 43278 -1028 43478 -1016
rect 43278 -1062 43290 -1028
rect 43466 -1062 43478 -1028
rect 43278 -1074 43478 -1062
rect 48268 -630 48468 -618
rect 48268 -664 48280 -630
rect 48456 -664 48468 -630
rect 48268 -676 48468 -664
rect 48268 -718 48468 -706
rect 48268 -752 48280 -718
rect 48456 -752 48468 -718
rect 48268 -764 48468 -752
rect 48268 -940 48468 -928
rect 48268 -974 48280 -940
rect 48456 -974 48468 -940
rect 48268 -986 48468 -974
rect 48268 -1028 48468 -1016
rect 48268 -1062 48280 -1028
rect 48456 -1062 48468 -1028
rect 48268 -1074 48468 -1062
rect 53258 -630 53458 -618
rect 53258 -664 53270 -630
rect 53446 -664 53458 -630
rect 53258 -676 53458 -664
rect 53258 -718 53458 -706
rect 53258 -752 53270 -718
rect 53446 -752 53458 -718
rect 53258 -764 53458 -752
rect 53258 -940 53458 -928
rect 53258 -974 53270 -940
rect 53446 -974 53458 -940
rect 53258 -986 53458 -974
rect 53258 -1028 53458 -1016
rect 53258 -1062 53270 -1028
rect 53446 -1062 53458 -1028
rect 53258 -1074 53458 -1062
rect 58248 -630 58448 -618
rect 58248 -664 58260 -630
rect 58436 -664 58448 -630
rect 58248 -676 58448 -664
rect 58248 -718 58448 -706
rect 58248 -752 58260 -718
rect 58436 -752 58448 -718
rect 58248 -764 58448 -752
rect 58248 -940 58448 -928
rect 58248 -974 58260 -940
rect 58436 -974 58448 -940
rect 58248 -986 58448 -974
rect 58248 -1028 58448 -1016
rect 58248 -1062 58260 -1028
rect 58436 -1062 58448 -1028
rect 58248 -1074 58448 -1062
rect 63238 -630 63438 -618
rect 63238 -664 63250 -630
rect 63426 -664 63438 -630
rect 63238 -676 63438 -664
rect 63238 -718 63438 -706
rect 63238 -752 63250 -718
rect 63426 -752 63438 -718
rect 63238 -764 63438 -752
rect 63238 -940 63438 -928
rect 63238 -974 63250 -940
rect 63426 -974 63438 -940
rect 63238 -986 63438 -974
rect 63238 -1028 63438 -1016
rect 63238 -1062 63250 -1028
rect 63426 -1062 63438 -1028
rect 63238 -1074 63438 -1062
rect 68228 -630 68428 -618
rect 68228 -664 68240 -630
rect 68416 -664 68428 -630
rect 68228 -676 68428 -664
rect 68228 -718 68428 -706
rect 68228 -752 68240 -718
rect 68416 -752 68428 -718
rect 68228 -764 68428 -752
rect 68228 -940 68428 -928
rect 68228 -974 68240 -940
rect 68416 -974 68428 -940
rect 68228 -986 68428 -974
rect 68228 -1028 68428 -1016
rect 68228 -1062 68240 -1028
rect 68416 -1062 68428 -1028
rect 68228 -1074 68428 -1062
rect 73218 -630 73418 -618
rect 73218 -664 73230 -630
rect 73406 -664 73418 -630
rect 73218 -676 73418 -664
rect 73218 -718 73418 -706
rect 73218 -752 73230 -718
rect 73406 -752 73418 -718
rect 73218 -764 73418 -752
rect 73218 -940 73418 -928
rect 73218 -974 73230 -940
rect 73406 -974 73418 -940
rect 73218 -986 73418 -974
rect 73218 -1028 73418 -1016
rect 73218 -1062 73230 -1028
rect 73406 -1062 73418 -1028
rect 73218 -1074 73418 -1062
rect 78208 -630 78408 -618
rect 78208 -664 78220 -630
rect 78396 -664 78408 -630
rect 78208 -676 78408 -664
rect 78208 -718 78408 -706
rect 78208 -752 78220 -718
rect 78396 -752 78408 -718
rect 78208 -764 78408 -752
rect 78208 -940 78408 -928
rect 78208 -974 78220 -940
rect 78396 -974 78408 -940
rect 78208 -986 78408 -974
rect 78208 -1028 78408 -1016
rect 78208 -1062 78220 -1028
rect 78396 -1062 78408 -1028
rect 78208 -1074 78408 -1062
rect 82928 -630 83128 -618
rect 82928 -664 82940 -630
rect 83116 -664 83128 -630
rect 82928 -676 83128 -664
rect 82928 -718 83128 -706
rect 82928 -752 82940 -718
rect 83116 -752 83128 -718
rect 82928 -764 83128 -752
rect 82928 -940 83128 -928
rect 82928 -974 82940 -940
rect 83116 -974 83128 -940
rect 82928 -986 83128 -974
rect 82928 -1028 83128 -1016
rect 82928 -1062 82940 -1028
rect 83116 -1062 83128 -1028
rect 82928 -1074 83128 -1062
<< ndiffc >>
rect 2872 28406 3048 28440
rect 2872 28318 3048 28352
rect 2872 28096 3048 28130
rect 2872 28008 3048 28042
rect 7862 28406 8038 28440
rect 7862 28318 8038 28352
rect 7862 28096 8038 28130
rect 7862 28008 8038 28042
rect 12852 28406 13028 28440
rect 12852 28318 13028 28352
rect 12852 28096 13028 28130
rect 12852 28008 13028 28042
rect 17842 28406 18018 28440
rect 17842 28318 18018 28352
rect 17842 28096 18018 28130
rect 17842 28008 18018 28042
rect 22832 28406 23008 28440
rect 22832 28318 23008 28352
rect 22832 28096 23008 28130
rect 22832 28008 23008 28042
rect 27822 28406 27998 28440
rect 27822 28318 27998 28352
rect 27822 28096 27998 28130
rect 27822 28008 27998 28042
rect 32812 28406 32988 28440
rect 32812 28318 32988 28352
rect 32812 28096 32988 28130
rect 32812 28008 32988 28042
rect 37802 28406 37978 28440
rect 37802 28318 37978 28352
rect 37802 28096 37978 28130
rect 37802 28008 37978 28042
rect 42792 28406 42968 28440
rect 42792 28318 42968 28352
rect 42792 28096 42968 28130
rect 42792 28008 42968 28042
rect 47782 28406 47958 28440
rect 47782 28318 47958 28352
rect 47782 28096 47958 28130
rect 47782 28008 47958 28042
rect 52772 28406 52948 28440
rect 52772 28318 52948 28352
rect 52772 28096 52948 28130
rect 52772 28008 52948 28042
rect 57762 28406 57938 28440
rect 57762 28318 57938 28352
rect 57762 28096 57938 28130
rect 57762 28008 57938 28042
rect 62752 28406 62928 28440
rect 62752 28318 62928 28352
rect 62752 28096 62928 28130
rect 62752 28008 62928 28042
rect 67742 28406 67918 28440
rect 67742 28318 67918 28352
rect 67742 28096 67918 28130
rect 67742 28008 67918 28042
rect 72732 28406 72908 28440
rect 72732 28318 72908 28352
rect 72732 28096 72908 28130
rect 72732 28008 72908 28042
rect 77722 28406 77898 28440
rect 77722 28318 77898 28352
rect 77722 28096 77898 28130
rect 77722 28008 77898 28042
rect 82442 28406 82618 28440
rect 82442 28318 82618 28352
rect 82442 28096 82618 28130
rect 82442 28008 82618 28042
rect 82442 26696 82618 26730
rect 82442 26608 82618 26642
rect 82442 26386 82618 26420
rect 82442 26298 82618 26332
rect 82442 24986 82618 25020
rect 82442 24898 82618 24932
rect 82442 24676 82618 24710
rect 82442 24588 82618 24622
rect -1848 23276 -1672 23310
rect -1848 23188 -1672 23222
rect -1848 22966 -1672 23000
rect -1848 22878 -1672 22912
rect 82442 23276 82618 23310
rect 82442 23188 82618 23222
rect 82442 22966 82618 23000
rect 82442 22878 82618 22912
rect -1848 21566 -1672 21600
rect -1848 21478 -1672 21512
rect -1848 21256 -1672 21290
rect -1848 21168 -1672 21202
rect 82442 21566 82618 21600
rect 82442 21478 82618 21512
rect 82442 21256 82618 21290
rect 82442 21168 82618 21202
rect -1848 19856 -1672 19890
rect -1848 19768 -1672 19802
rect -1848 19546 -1672 19580
rect -1848 19458 -1672 19492
rect 82442 19856 82618 19890
rect 82442 19768 82618 19802
rect 82442 19546 82618 19580
rect 82442 19458 82618 19492
rect -1848 18146 -1672 18180
rect -1848 18058 -1672 18092
rect -1848 17836 -1672 17870
rect -1848 17748 -1672 17782
rect 82442 18146 82618 18180
rect 82442 18058 82618 18092
rect 82442 17836 82618 17870
rect 82442 17748 82618 17782
rect -1848 16436 -1672 16470
rect -1848 16348 -1672 16382
rect -1848 16126 -1672 16160
rect -1848 16038 -1672 16072
rect 82442 16436 82618 16470
rect 82442 16348 82618 16382
rect 82442 16126 82618 16160
rect 82442 16038 82618 16072
rect -1848 14726 -1672 14760
rect -1848 14638 -1672 14672
rect -1848 14416 -1672 14450
rect -1848 14328 -1672 14362
rect 82442 14726 82618 14760
rect 82442 14638 82618 14672
rect 82442 14416 82618 14450
rect 82442 14328 82618 14362
rect -1848 13016 -1672 13050
rect -1848 12928 -1672 12962
rect -1848 12706 -1672 12740
rect -1848 12618 -1672 12652
rect 82442 13016 82618 13050
rect 82442 12928 82618 12962
rect 82442 12706 82618 12740
rect 82442 12618 82618 12652
rect -1848 11306 -1672 11340
rect -1848 11218 -1672 11252
rect -1848 10996 -1672 11030
rect -1848 10908 -1672 10942
rect 82442 11306 82618 11340
rect 82442 11218 82618 11252
rect 82442 10996 82618 11030
rect 82442 10908 82618 10942
rect -1848 9596 -1672 9630
rect -1848 9508 -1672 9542
rect -1848 9286 -1672 9320
rect -1848 9198 -1672 9232
rect 82442 9596 82618 9630
rect 82442 9508 82618 9542
rect 82442 9286 82618 9320
rect 82442 9198 82618 9232
rect -1848 7886 -1672 7920
rect -1848 7798 -1672 7832
rect -1848 7576 -1672 7610
rect -1848 7488 -1672 7522
rect 82442 7886 82618 7920
rect 82442 7798 82618 7832
rect 82442 7576 82618 7610
rect 82442 7488 82618 7522
rect -1848 6176 -1672 6210
rect -1848 6088 -1672 6122
rect -1848 5866 -1672 5900
rect -1848 5778 -1672 5812
rect 82442 6176 82618 6210
rect 82442 6088 82618 6122
rect 82442 5866 82618 5900
rect 82442 5778 82618 5812
rect -1848 4466 -1672 4500
rect -1848 4378 -1672 4412
rect -1848 4156 -1672 4190
rect -1848 4068 -1672 4102
rect 82442 4466 82618 4500
rect 82442 4378 82618 4412
rect 82442 4156 82618 4190
rect 82442 4068 82618 4102
rect -1848 2756 -1672 2790
rect -1848 2668 -1672 2702
rect -1848 2446 -1672 2480
rect -1848 2358 -1672 2392
rect 82442 2756 82618 2790
rect 82442 2668 82618 2702
rect 82442 2446 82618 2480
rect 82442 2358 82618 2392
rect -1848 1046 -1672 1080
rect -1848 958 -1672 992
rect -1848 736 -1672 770
rect -1848 648 -1672 682
rect 82442 1046 82618 1080
rect 82442 958 82618 992
rect 82442 736 82618 770
rect 82442 648 82618 682
rect -1848 -664 -1672 -630
rect -1848 -752 -1672 -718
rect -1848 -974 -1672 -940
rect -1848 -1062 -1672 -1028
rect 2872 -664 3048 -630
rect 2872 -752 3048 -718
rect 2872 -974 3048 -940
rect 2872 -1062 3048 -1028
rect 7862 -664 8038 -630
rect 7862 -752 8038 -718
rect 7862 -974 8038 -940
rect 7862 -1062 8038 -1028
rect 12852 -664 13028 -630
rect 12852 -752 13028 -718
rect 12852 -974 13028 -940
rect 12852 -1062 13028 -1028
rect 17842 -664 18018 -630
rect 17842 -752 18018 -718
rect 17842 -974 18018 -940
rect 17842 -1062 18018 -1028
rect 22832 -664 23008 -630
rect 22832 -752 23008 -718
rect 22832 -974 23008 -940
rect 22832 -1062 23008 -1028
rect 27822 -664 27998 -630
rect 27822 -752 27998 -718
rect 27822 -974 27998 -940
rect 27822 -1062 27998 -1028
rect 32812 -664 32988 -630
rect 32812 -752 32988 -718
rect 32812 -974 32988 -940
rect 32812 -1062 32988 -1028
rect 37802 -664 37978 -630
rect 37802 -752 37978 -718
rect 37802 -974 37978 -940
rect 37802 -1062 37978 -1028
rect 42792 -664 42968 -630
rect 42792 -752 42968 -718
rect 42792 -974 42968 -940
rect 42792 -1062 42968 -1028
rect 47782 -664 47958 -630
rect 47782 -752 47958 -718
rect 47782 -974 47958 -940
rect 47782 -1062 47958 -1028
rect 52772 -664 52948 -630
rect 52772 -752 52948 -718
rect 52772 -974 52948 -940
rect 52772 -1062 52948 -1028
rect 57762 -664 57938 -630
rect 57762 -752 57938 -718
rect 57762 -974 57938 -940
rect 57762 -1062 57938 -1028
rect 62752 -664 62928 -630
rect 62752 -752 62928 -718
rect 62752 -974 62928 -940
rect 62752 -1062 62928 -1028
rect 67742 -664 67918 -630
rect 67742 -752 67918 -718
rect 67742 -974 67918 -940
rect 67742 -1062 67918 -1028
rect 72732 -664 72908 -630
rect 72732 -752 72908 -718
rect 72732 -974 72908 -940
rect 72732 -1062 72908 -1028
rect 77722 -664 77898 -630
rect 77722 -752 77898 -718
rect 77722 -974 77898 -940
rect 77722 -1062 77898 -1028
rect 82442 -664 82618 -630
rect 82442 -752 82618 -718
rect 82442 -974 82618 -940
rect 82442 -1062 82618 -1028
<< pdiffc >>
rect 3370 28406 3546 28440
rect 3370 28318 3546 28352
rect 3370 28096 3546 28130
rect 3370 28008 3546 28042
rect 8360 28406 8536 28440
rect 8360 28318 8536 28352
rect 8360 28096 8536 28130
rect 8360 28008 8536 28042
rect 13350 28406 13526 28440
rect 13350 28318 13526 28352
rect 13350 28096 13526 28130
rect 13350 28008 13526 28042
rect 18340 28406 18516 28440
rect 18340 28318 18516 28352
rect 18340 28096 18516 28130
rect 18340 28008 18516 28042
rect 23330 28406 23506 28440
rect 23330 28318 23506 28352
rect 23330 28096 23506 28130
rect 23330 28008 23506 28042
rect 28320 28406 28496 28440
rect 28320 28318 28496 28352
rect 28320 28096 28496 28130
rect 28320 28008 28496 28042
rect 33310 28406 33486 28440
rect 33310 28318 33486 28352
rect 33310 28096 33486 28130
rect 33310 28008 33486 28042
rect 38300 28406 38476 28440
rect 38300 28318 38476 28352
rect 38300 28096 38476 28130
rect 38300 28008 38476 28042
rect 43290 28406 43466 28440
rect 43290 28318 43466 28352
rect 43290 28096 43466 28130
rect 43290 28008 43466 28042
rect 48280 28406 48456 28440
rect 48280 28318 48456 28352
rect 48280 28096 48456 28130
rect 48280 28008 48456 28042
rect 53270 28406 53446 28440
rect 53270 28318 53446 28352
rect 53270 28096 53446 28130
rect 53270 28008 53446 28042
rect 58260 28406 58436 28440
rect 58260 28318 58436 28352
rect 58260 28096 58436 28130
rect 58260 28008 58436 28042
rect 63250 28406 63426 28440
rect 63250 28318 63426 28352
rect 63250 28096 63426 28130
rect 63250 28008 63426 28042
rect 68240 28406 68416 28440
rect 68240 28318 68416 28352
rect 68240 28096 68416 28130
rect 68240 28008 68416 28042
rect 73230 28406 73406 28440
rect 73230 28318 73406 28352
rect 73230 28096 73406 28130
rect 73230 28008 73406 28042
rect 78220 28406 78396 28440
rect 78220 28318 78396 28352
rect 78220 28096 78396 28130
rect 78220 28008 78396 28042
rect 82940 28406 83116 28440
rect 82940 28318 83116 28352
rect 82940 28096 83116 28130
rect 82940 28008 83116 28042
rect 82940 26696 83116 26730
rect 82940 26608 83116 26642
rect 82940 26386 83116 26420
rect 82940 26298 83116 26332
rect 82940 24986 83116 25020
rect 82940 24898 83116 24932
rect 82940 24676 83116 24710
rect 82940 24588 83116 24622
rect -1350 23276 -1174 23310
rect -1350 23188 -1174 23222
rect -1350 22966 -1174 23000
rect -1350 22878 -1174 22912
rect 82940 23276 83116 23310
rect 82940 23188 83116 23222
rect 82940 22966 83116 23000
rect 82940 22878 83116 22912
rect -1350 21566 -1174 21600
rect -1350 21478 -1174 21512
rect -1350 21256 -1174 21290
rect -1350 21168 -1174 21202
rect 82940 21566 83116 21600
rect 82940 21478 83116 21512
rect 82940 21256 83116 21290
rect 82940 21168 83116 21202
rect -1350 19856 -1174 19890
rect -1350 19768 -1174 19802
rect -1350 19546 -1174 19580
rect -1350 19458 -1174 19492
rect 82940 19856 83116 19890
rect 82940 19768 83116 19802
rect 82940 19546 83116 19580
rect 82940 19458 83116 19492
rect -1350 18146 -1174 18180
rect -1350 18058 -1174 18092
rect -1350 17836 -1174 17870
rect -1350 17748 -1174 17782
rect 82940 18146 83116 18180
rect 82940 18058 83116 18092
rect 82940 17836 83116 17870
rect 82940 17748 83116 17782
rect -1350 16436 -1174 16470
rect -1350 16348 -1174 16382
rect -1350 16126 -1174 16160
rect -1350 16038 -1174 16072
rect 82940 16436 83116 16470
rect 82940 16348 83116 16382
rect 82940 16126 83116 16160
rect 82940 16038 83116 16072
rect -1350 14726 -1174 14760
rect -1350 14638 -1174 14672
rect -1350 14416 -1174 14450
rect -1350 14328 -1174 14362
rect 82940 14726 83116 14760
rect 82940 14638 83116 14672
rect 82940 14416 83116 14450
rect 82940 14328 83116 14362
rect -1350 13016 -1174 13050
rect -1350 12928 -1174 12962
rect -1350 12706 -1174 12740
rect -1350 12618 -1174 12652
rect 82940 13016 83116 13050
rect 82940 12928 83116 12962
rect 82940 12706 83116 12740
rect 82940 12618 83116 12652
rect -1350 11306 -1174 11340
rect -1350 11218 -1174 11252
rect -1350 10996 -1174 11030
rect -1350 10908 -1174 10942
rect 82940 11306 83116 11340
rect 82940 11218 83116 11252
rect 82940 10996 83116 11030
rect 82940 10908 83116 10942
rect -1350 9596 -1174 9630
rect -1350 9508 -1174 9542
rect -1350 9286 -1174 9320
rect -1350 9198 -1174 9232
rect 82940 9596 83116 9630
rect 82940 9508 83116 9542
rect 82940 9286 83116 9320
rect 82940 9198 83116 9232
rect -1350 7886 -1174 7920
rect -1350 7798 -1174 7832
rect -1350 7576 -1174 7610
rect -1350 7488 -1174 7522
rect 82940 7886 83116 7920
rect 82940 7798 83116 7832
rect 82940 7576 83116 7610
rect 82940 7488 83116 7522
rect -1350 6176 -1174 6210
rect -1350 6088 -1174 6122
rect -1350 5866 -1174 5900
rect -1350 5778 -1174 5812
rect 82940 6176 83116 6210
rect 82940 6088 83116 6122
rect 82940 5866 83116 5900
rect 82940 5778 83116 5812
rect -1350 4466 -1174 4500
rect -1350 4378 -1174 4412
rect -1350 4156 -1174 4190
rect -1350 4068 -1174 4102
rect 82940 4466 83116 4500
rect 82940 4378 83116 4412
rect 82940 4156 83116 4190
rect 82940 4068 83116 4102
rect -1350 2756 -1174 2790
rect -1350 2668 -1174 2702
rect -1350 2446 -1174 2480
rect -1350 2358 -1174 2392
rect 82940 2756 83116 2790
rect 82940 2668 83116 2702
rect 82940 2446 83116 2480
rect 82940 2358 83116 2392
rect -1350 1046 -1174 1080
rect -1350 958 -1174 992
rect -1350 736 -1174 770
rect -1350 648 -1174 682
rect 82940 1046 83116 1080
rect 82940 958 83116 992
rect 82940 736 83116 770
rect 82940 648 83116 682
rect -1350 -664 -1174 -630
rect -1350 -752 -1174 -718
rect -1350 -974 -1174 -940
rect -1350 -1062 -1174 -1028
rect 3370 -664 3546 -630
rect 3370 -752 3546 -718
rect 3370 -974 3546 -940
rect 3370 -1062 3546 -1028
rect 8360 -664 8536 -630
rect 8360 -752 8536 -718
rect 8360 -974 8536 -940
rect 8360 -1062 8536 -1028
rect 13350 -664 13526 -630
rect 13350 -752 13526 -718
rect 13350 -974 13526 -940
rect 13350 -1062 13526 -1028
rect 18340 -664 18516 -630
rect 18340 -752 18516 -718
rect 18340 -974 18516 -940
rect 18340 -1062 18516 -1028
rect 23330 -664 23506 -630
rect 23330 -752 23506 -718
rect 23330 -974 23506 -940
rect 23330 -1062 23506 -1028
rect 28320 -664 28496 -630
rect 28320 -752 28496 -718
rect 28320 -974 28496 -940
rect 28320 -1062 28496 -1028
rect 33310 -664 33486 -630
rect 33310 -752 33486 -718
rect 33310 -974 33486 -940
rect 33310 -1062 33486 -1028
rect 38300 -664 38476 -630
rect 38300 -752 38476 -718
rect 38300 -974 38476 -940
rect 38300 -1062 38476 -1028
rect 43290 -664 43466 -630
rect 43290 -752 43466 -718
rect 43290 -974 43466 -940
rect 43290 -1062 43466 -1028
rect 48280 -664 48456 -630
rect 48280 -752 48456 -718
rect 48280 -974 48456 -940
rect 48280 -1062 48456 -1028
rect 53270 -664 53446 -630
rect 53270 -752 53446 -718
rect 53270 -974 53446 -940
rect 53270 -1062 53446 -1028
rect 58260 -664 58436 -630
rect 58260 -752 58436 -718
rect 58260 -974 58436 -940
rect 58260 -1062 58436 -1028
rect 63250 -664 63426 -630
rect 63250 -752 63426 -718
rect 63250 -974 63426 -940
rect 63250 -1062 63426 -1028
rect 68240 -664 68416 -630
rect 68240 -752 68416 -718
rect 68240 -974 68416 -940
rect 68240 -1062 68416 -1028
rect 73230 -664 73406 -630
rect 73230 -752 73406 -718
rect 73230 -974 73406 -940
rect 73230 -1062 73406 -1028
rect 78220 -664 78396 -630
rect 78220 -752 78396 -718
rect 78220 -974 78396 -940
rect 78220 -1062 78396 -1028
rect 82940 -664 83116 -630
rect 82940 -752 83116 -718
rect 82940 -974 83116 -940
rect 82940 -1062 83116 -1028
<< psubdiff >>
rect 2686 28520 3172 28554
rect 2686 28458 2720 28520
rect 2686 28244 2720 28300
rect 3138 28244 3172 28520
rect 2686 28204 3172 28244
rect 2686 28148 2720 28204
rect 2686 27928 2720 27990
rect 3138 27928 3172 28204
rect 2686 27894 3172 27928
rect 7676 28520 8162 28554
rect 7676 28458 7710 28520
rect 7676 28244 7710 28300
rect 8128 28244 8162 28520
rect 7676 28204 8162 28244
rect 7676 28148 7710 28204
rect 7676 27928 7710 27990
rect 8128 27928 8162 28204
rect 7676 27894 8162 27928
rect 12666 28520 13152 28554
rect 12666 28458 12700 28520
rect 12666 28244 12700 28300
rect 13118 28244 13152 28520
rect 12666 28204 13152 28244
rect 12666 28148 12700 28204
rect 12666 27928 12700 27990
rect 13118 27928 13152 28204
rect 12666 27894 13152 27928
rect 17656 28520 18142 28554
rect 17656 28458 17690 28520
rect 17656 28244 17690 28300
rect 18108 28244 18142 28520
rect 17656 28204 18142 28244
rect 17656 28148 17690 28204
rect 17656 27928 17690 27990
rect 18108 27928 18142 28204
rect 17656 27894 18142 27928
rect 22646 28520 23132 28554
rect 22646 28458 22680 28520
rect 22646 28244 22680 28300
rect 23098 28244 23132 28520
rect 22646 28204 23132 28244
rect 22646 28148 22680 28204
rect 22646 27928 22680 27990
rect 23098 27928 23132 28204
rect 22646 27894 23132 27928
rect 27636 28520 28122 28554
rect 27636 28458 27670 28520
rect 27636 28244 27670 28300
rect 28088 28244 28122 28520
rect 27636 28204 28122 28244
rect 27636 28148 27670 28204
rect 27636 27928 27670 27990
rect 28088 27928 28122 28204
rect 27636 27894 28122 27928
rect 32626 28520 33112 28554
rect 32626 28458 32660 28520
rect 32626 28244 32660 28300
rect 33078 28244 33112 28520
rect 32626 28204 33112 28244
rect 32626 28148 32660 28204
rect 32626 27928 32660 27990
rect 33078 27928 33112 28204
rect 32626 27894 33112 27928
rect 37616 28520 38102 28554
rect 37616 28458 37650 28520
rect 37616 28244 37650 28300
rect 38068 28244 38102 28520
rect 37616 28204 38102 28244
rect 37616 28148 37650 28204
rect 37616 27928 37650 27990
rect 38068 27928 38102 28204
rect 37616 27894 38102 27928
rect 42606 28520 43092 28554
rect 42606 28458 42640 28520
rect 42606 28244 42640 28300
rect 43058 28244 43092 28520
rect 42606 28204 43092 28244
rect 42606 28148 42640 28204
rect 42606 27928 42640 27990
rect 43058 27928 43092 28204
rect 42606 27894 43092 27928
rect 47596 28520 48082 28554
rect 47596 28458 47630 28520
rect 47596 28244 47630 28300
rect 48048 28244 48082 28520
rect 47596 28204 48082 28244
rect 47596 28148 47630 28204
rect 47596 27928 47630 27990
rect 48048 27928 48082 28204
rect 47596 27894 48082 27928
rect 52586 28520 53072 28554
rect 52586 28458 52620 28520
rect 52586 28244 52620 28300
rect 53038 28244 53072 28520
rect 52586 28204 53072 28244
rect 52586 28148 52620 28204
rect 52586 27928 52620 27990
rect 53038 27928 53072 28204
rect 52586 27894 53072 27928
rect 57576 28520 58062 28554
rect 57576 28458 57610 28520
rect 57576 28244 57610 28300
rect 58028 28244 58062 28520
rect 57576 28204 58062 28244
rect 57576 28148 57610 28204
rect 57576 27928 57610 27990
rect 58028 27928 58062 28204
rect 57576 27894 58062 27928
rect 62566 28520 63052 28554
rect 62566 28458 62600 28520
rect 62566 28244 62600 28300
rect 63018 28244 63052 28520
rect 62566 28204 63052 28244
rect 62566 28148 62600 28204
rect 62566 27928 62600 27990
rect 63018 27928 63052 28204
rect 62566 27894 63052 27928
rect 67556 28520 68042 28554
rect 67556 28458 67590 28520
rect 67556 28244 67590 28300
rect 68008 28244 68042 28520
rect 67556 28204 68042 28244
rect 67556 28148 67590 28204
rect 67556 27928 67590 27990
rect 68008 27928 68042 28204
rect 67556 27894 68042 27928
rect 72546 28520 73032 28554
rect 72546 28458 72580 28520
rect 72546 28244 72580 28300
rect 72998 28244 73032 28520
rect 72546 28204 73032 28244
rect 72546 28148 72580 28204
rect 72546 27928 72580 27990
rect 72998 27928 73032 28204
rect 72546 27894 73032 27928
rect 77536 28520 78022 28554
rect 77536 28458 77570 28520
rect 77536 28244 77570 28300
rect 77988 28244 78022 28520
rect 77536 28204 78022 28244
rect 77536 28148 77570 28204
rect 77536 27928 77570 27990
rect 77988 27928 78022 28204
rect 77536 27894 78022 27928
rect 82256 28520 82742 28554
rect 82256 28458 82290 28520
rect 82256 28244 82290 28300
rect 82708 28244 82742 28520
rect 82256 28204 82742 28244
rect 82256 28148 82290 28204
rect 82256 27928 82290 27990
rect 82708 27928 82742 28204
rect 82256 27894 82742 27928
rect 82256 26810 82742 26844
rect 82256 26748 82290 26810
rect 82256 26534 82290 26590
rect 82708 26534 82742 26810
rect 82256 26494 82742 26534
rect 82256 26438 82290 26494
rect 82256 26218 82290 26280
rect 82708 26218 82742 26494
rect 82256 26184 82742 26218
rect 82256 25100 82742 25134
rect 82256 25038 82290 25100
rect 82256 24824 82290 24880
rect 82708 24824 82742 25100
rect 82256 24784 82742 24824
rect 82256 24728 82290 24784
rect 82256 24508 82290 24570
rect 82708 24508 82742 24784
rect 82256 24474 82742 24508
rect -2034 23390 -1548 23424
rect -2034 23328 -2000 23390
rect -2034 23114 -2000 23170
rect -1582 23114 -1548 23390
rect -2034 23074 -1548 23114
rect -2034 23018 -2000 23074
rect -2034 22798 -2000 22860
rect -1582 22798 -1548 23074
rect -2034 22764 -1548 22798
rect 82256 23390 82742 23424
rect 82256 23328 82290 23390
rect 82256 23114 82290 23170
rect 82708 23114 82742 23390
rect 82256 23074 82742 23114
rect 82256 23018 82290 23074
rect 82256 22798 82290 22860
rect 82708 22798 82742 23074
rect 82256 22764 82742 22798
rect -2034 21680 -1548 21714
rect -2034 21618 -2000 21680
rect -2034 21404 -2000 21460
rect -1582 21404 -1548 21680
rect -2034 21364 -1548 21404
rect -2034 21308 -2000 21364
rect -2034 21088 -2000 21150
rect -1582 21088 -1548 21364
rect -2034 21054 -1548 21088
rect 82256 21680 82742 21714
rect 82256 21618 82290 21680
rect 82256 21404 82290 21460
rect 82708 21404 82742 21680
rect 82256 21364 82742 21404
rect 82256 21308 82290 21364
rect 82256 21088 82290 21150
rect 82708 21088 82742 21364
rect 82256 21054 82742 21088
rect -2034 19970 -1548 20004
rect -2034 19908 -2000 19970
rect -2034 19694 -2000 19750
rect -1582 19694 -1548 19970
rect -2034 19654 -1548 19694
rect -2034 19598 -2000 19654
rect -2034 19378 -2000 19440
rect -1582 19378 -1548 19654
rect -2034 19344 -1548 19378
rect 82256 19970 82742 20004
rect 82256 19908 82290 19970
rect 82256 19694 82290 19750
rect 82708 19694 82742 19970
rect 82256 19654 82742 19694
rect 82256 19598 82290 19654
rect 82256 19378 82290 19440
rect 82708 19378 82742 19654
rect 82256 19344 82742 19378
rect -2034 18260 -1548 18294
rect -2034 18198 -2000 18260
rect -2034 17984 -2000 18040
rect -1582 17984 -1548 18260
rect -2034 17944 -1548 17984
rect -2034 17888 -2000 17944
rect -2034 17668 -2000 17730
rect -1582 17668 -1548 17944
rect -2034 17634 -1548 17668
rect 82256 18260 82742 18294
rect 82256 18198 82290 18260
rect 82256 17984 82290 18040
rect 82708 17984 82742 18260
rect 82256 17944 82742 17984
rect 82256 17888 82290 17944
rect 82256 17668 82290 17730
rect 82708 17668 82742 17944
rect 82256 17634 82742 17668
rect -2034 16550 -1548 16584
rect -2034 16488 -2000 16550
rect -2034 16274 -2000 16330
rect -1582 16274 -1548 16550
rect -2034 16234 -1548 16274
rect -2034 16178 -2000 16234
rect -2034 15958 -2000 16020
rect -1582 15958 -1548 16234
rect -2034 15924 -1548 15958
rect 82256 16550 82742 16584
rect 82256 16488 82290 16550
rect 82256 16274 82290 16330
rect 82708 16274 82742 16550
rect 82256 16234 82742 16274
rect 82256 16178 82290 16234
rect 82256 15958 82290 16020
rect 82708 15958 82742 16234
rect 82256 15924 82742 15958
rect -2034 14840 -1548 14874
rect -2034 14778 -2000 14840
rect -2034 14564 -2000 14620
rect -1582 14564 -1548 14840
rect -2034 14524 -1548 14564
rect -2034 14468 -2000 14524
rect -2034 14248 -2000 14310
rect -1582 14248 -1548 14524
rect -2034 14214 -1548 14248
rect 82256 14840 82742 14874
rect 82256 14778 82290 14840
rect 82256 14564 82290 14620
rect 82708 14564 82742 14840
rect 82256 14524 82742 14564
rect 82256 14468 82290 14524
rect 82256 14248 82290 14310
rect 82708 14248 82742 14524
rect 82256 14214 82742 14248
rect -2034 13130 -1548 13164
rect -2034 13068 -2000 13130
rect -2034 12854 -2000 12910
rect -1582 12854 -1548 13130
rect -2034 12814 -1548 12854
rect -2034 12758 -2000 12814
rect -2034 12538 -2000 12600
rect -1582 12538 -1548 12814
rect -2034 12504 -1548 12538
rect 82256 13130 82742 13164
rect 82256 13068 82290 13130
rect 82256 12854 82290 12910
rect 82708 12854 82742 13130
rect 82256 12814 82742 12854
rect 82256 12758 82290 12814
rect 82256 12538 82290 12600
rect 82708 12538 82742 12814
rect 82256 12504 82742 12538
rect -2034 11420 -1548 11454
rect -2034 11358 -2000 11420
rect -2034 11144 -2000 11200
rect -1582 11144 -1548 11420
rect -2034 11104 -1548 11144
rect -2034 11048 -2000 11104
rect -2034 10828 -2000 10890
rect -1582 10828 -1548 11104
rect -2034 10794 -1548 10828
rect 82256 11420 82742 11454
rect 82256 11358 82290 11420
rect 82256 11144 82290 11200
rect 82708 11144 82742 11420
rect 82256 11104 82742 11144
rect 82256 11048 82290 11104
rect 82256 10828 82290 10890
rect 82708 10828 82742 11104
rect 82256 10794 82742 10828
rect -2034 9710 -1548 9744
rect -2034 9648 -2000 9710
rect -2034 9434 -2000 9490
rect -1582 9434 -1548 9710
rect -2034 9394 -1548 9434
rect -2034 9338 -2000 9394
rect -2034 9118 -2000 9180
rect -1582 9118 -1548 9394
rect -2034 9084 -1548 9118
rect 82256 9710 82742 9744
rect 82256 9648 82290 9710
rect 82256 9434 82290 9490
rect 82708 9434 82742 9710
rect 82256 9394 82742 9434
rect 82256 9338 82290 9394
rect 82256 9118 82290 9180
rect 82708 9118 82742 9394
rect 82256 9084 82742 9118
rect -2034 8000 -1548 8034
rect -2034 7938 -2000 8000
rect -2034 7724 -2000 7780
rect -1582 7724 -1548 8000
rect -2034 7684 -1548 7724
rect -2034 7628 -2000 7684
rect -2034 7408 -2000 7470
rect -1582 7408 -1548 7684
rect -2034 7374 -1548 7408
rect 82256 8000 82742 8034
rect 82256 7938 82290 8000
rect 82256 7724 82290 7780
rect 82708 7724 82742 8000
rect 82256 7684 82742 7724
rect 82256 7628 82290 7684
rect 82256 7408 82290 7470
rect 82708 7408 82742 7684
rect 82256 7374 82742 7408
rect -2034 6290 -1548 6324
rect -2034 6228 -2000 6290
rect -2034 6014 -2000 6070
rect -1582 6014 -1548 6290
rect -2034 5974 -1548 6014
rect -2034 5918 -2000 5974
rect -2034 5698 -2000 5760
rect -1582 5698 -1548 5974
rect -2034 5664 -1548 5698
rect 82256 6290 82742 6324
rect 82256 6228 82290 6290
rect 82256 6014 82290 6070
rect 82708 6014 82742 6290
rect 82256 5974 82742 6014
rect 82256 5918 82290 5974
rect 82256 5698 82290 5760
rect 82708 5698 82742 5974
rect 82256 5664 82742 5698
rect -2034 4580 -1548 4614
rect -2034 4518 -2000 4580
rect -2034 4304 -2000 4360
rect -1582 4304 -1548 4580
rect -2034 4264 -1548 4304
rect -2034 4208 -2000 4264
rect -2034 3988 -2000 4050
rect -1582 3988 -1548 4264
rect -2034 3954 -1548 3988
rect 82256 4580 82742 4614
rect 82256 4518 82290 4580
rect 82256 4304 82290 4360
rect 82708 4304 82742 4580
rect 82256 4264 82742 4304
rect 82256 4208 82290 4264
rect 82256 3988 82290 4050
rect 82708 3988 82742 4264
rect 82256 3954 82742 3988
rect -2034 2870 -1548 2904
rect -2034 2808 -2000 2870
rect -2034 2594 -2000 2650
rect -1582 2594 -1548 2870
rect -2034 2554 -1548 2594
rect -2034 2498 -2000 2554
rect -2034 2278 -2000 2340
rect -1582 2278 -1548 2554
rect -2034 2244 -1548 2278
rect 82256 2870 82742 2904
rect 82256 2808 82290 2870
rect 82256 2594 82290 2650
rect 82708 2594 82742 2870
rect 82256 2554 82742 2594
rect 82256 2498 82290 2554
rect 82256 2278 82290 2340
rect 82708 2278 82742 2554
rect 82256 2244 82742 2278
rect -2034 1160 -1548 1194
rect -2034 1098 -2000 1160
rect -2034 884 -2000 940
rect -1582 884 -1548 1160
rect -2034 844 -1548 884
rect -2034 788 -2000 844
rect -2034 568 -2000 630
rect -1582 568 -1548 844
rect -2034 534 -1548 568
rect 82256 1160 82742 1194
rect 82256 1098 82290 1160
rect 82256 884 82290 940
rect 82708 884 82742 1160
rect 82256 844 82742 884
rect 82256 788 82290 844
rect 82256 568 82290 630
rect 82708 568 82742 844
rect 82256 534 82742 568
rect -2034 -550 -1548 -516
rect -2034 -612 -2000 -550
rect -2034 -826 -2000 -770
rect -1582 -826 -1548 -550
rect -2034 -866 -1548 -826
rect -2034 -922 -2000 -866
rect -2034 -1142 -2000 -1080
rect -1582 -1142 -1548 -866
rect -2034 -1176 -1548 -1142
rect 2686 -550 3172 -516
rect 2686 -612 2720 -550
rect 2686 -826 2720 -770
rect 3138 -826 3172 -550
rect 2686 -866 3172 -826
rect 2686 -922 2720 -866
rect 2686 -1142 2720 -1080
rect 3138 -1142 3172 -866
rect 2686 -1176 3172 -1142
rect 7676 -550 8162 -516
rect 7676 -612 7710 -550
rect 7676 -826 7710 -770
rect 8128 -826 8162 -550
rect 7676 -866 8162 -826
rect 7676 -922 7710 -866
rect 7676 -1142 7710 -1080
rect 8128 -1142 8162 -866
rect 7676 -1176 8162 -1142
rect 12666 -550 13152 -516
rect 12666 -612 12700 -550
rect 12666 -826 12700 -770
rect 13118 -826 13152 -550
rect 12666 -866 13152 -826
rect 12666 -922 12700 -866
rect 12666 -1142 12700 -1080
rect 13118 -1142 13152 -866
rect 12666 -1176 13152 -1142
rect 17656 -550 18142 -516
rect 17656 -612 17690 -550
rect 17656 -826 17690 -770
rect 18108 -826 18142 -550
rect 17656 -866 18142 -826
rect 17656 -922 17690 -866
rect 17656 -1142 17690 -1080
rect 18108 -1142 18142 -866
rect 17656 -1176 18142 -1142
rect 22646 -550 23132 -516
rect 22646 -612 22680 -550
rect 22646 -826 22680 -770
rect 23098 -826 23132 -550
rect 22646 -866 23132 -826
rect 22646 -922 22680 -866
rect 22646 -1142 22680 -1080
rect 23098 -1142 23132 -866
rect 22646 -1176 23132 -1142
rect 27636 -550 28122 -516
rect 27636 -612 27670 -550
rect 27636 -826 27670 -770
rect 28088 -826 28122 -550
rect 27636 -866 28122 -826
rect 27636 -922 27670 -866
rect 27636 -1142 27670 -1080
rect 28088 -1142 28122 -866
rect 27636 -1176 28122 -1142
rect 32626 -550 33112 -516
rect 32626 -612 32660 -550
rect 32626 -826 32660 -770
rect 33078 -826 33112 -550
rect 32626 -866 33112 -826
rect 32626 -922 32660 -866
rect 32626 -1142 32660 -1080
rect 33078 -1142 33112 -866
rect 32626 -1176 33112 -1142
rect 37616 -550 38102 -516
rect 37616 -612 37650 -550
rect 37616 -826 37650 -770
rect 38068 -826 38102 -550
rect 37616 -866 38102 -826
rect 37616 -922 37650 -866
rect 37616 -1142 37650 -1080
rect 38068 -1142 38102 -866
rect 37616 -1176 38102 -1142
rect 42606 -550 43092 -516
rect 42606 -612 42640 -550
rect 42606 -826 42640 -770
rect 43058 -826 43092 -550
rect 42606 -866 43092 -826
rect 42606 -922 42640 -866
rect 42606 -1142 42640 -1080
rect 43058 -1142 43092 -866
rect 42606 -1176 43092 -1142
rect 47596 -550 48082 -516
rect 47596 -612 47630 -550
rect 47596 -826 47630 -770
rect 48048 -826 48082 -550
rect 47596 -866 48082 -826
rect 47596 -922 47630 -866
rect 47596 -1142 47630 -1080
rect 48048 -1142 48082 -866
rect 47596 -1176 48082 -1142
rect 52586 -550 53072 -516
rect 52586 -612 52620 -550
rect 52586 -826 52620 -770
rect 53038 -826 53072 -550
rect 52586 -866 53072 -826
rect 52586 -922 52620 -866
rect 52586 -1142 52620 -1080
rect 53038 -1142 53072 -866
rect 52586 -1176 53072 -1142
rect 57576 -550 58062 -516
rect 57576 -612 57610 -550
rect 57576 -826 57610 -770
rect 58028 -826 58062 -550
rect 57576 -866 58062 -826
rect 57576 -922 57610 -866
rect 57576 -1142 57610 -1080
rect 58028 -1142 58062 -866
rect 57576 -1176 58062 -1142
rect 62566 -550 63052 -516
rect 62566 -612 62600 -550
rect 62566 -826 62600 -770
rect 63018 -826 63052 -550
rect 62566 -866 63052 -826
rect 62566 -922 62600 -866
rect 62566 -1142 62600 -1080
rect 63018 -1142 63052 -866
rect 62566 -1176 63052 -1142
rect 67556 -550 68042 -516
rect 67556 -612 67590 -550
rect 67556 -826 67590 -770
rect 68008 -826 68042 -550
rect 67556 -866 68042 -826
rect 67556 -922 67590 -866
rect 67556 -1142 67590 -1080
rect 68008 -1142 68042 -866
rect 67556 -1176 68042 -1142
rect 72546 -550 73032 -516
rect 72546 -612 72580 -550
rect 72546 -826 72580 -770
rect 72998 -826 73032 -550
rect 72546 -866 73032 -826
rect 72546 -922 72580 -866
rect 72546 -1142 72580 -1080
rect 72998 -1142 73032 -866
rect 72546 -1176 73032 -1142
rect 77536 -550 78022 -516
rect 77536 -612 77570 -550
rect 77536 -826 77570 -770
rect 77988 -826 78022 -550
rect 77536 -866 78022 -826
rect 77536 -922 77570 -866
rect 77536 -1142 77570 -1080
rect 77988 -1142 78022 -866
rect 77536 -1176 78022 -1142
rect 82256 -550 82742 -516
rect 82256 -612 82290 -550
rect 82256 -826 82290 -770
rect 82708 -826 82742 -550
rect 82256 -866 82742 -826
rect 82256 -922 82290 -866
rect 82256 -1142 82290 -1080
rect 82708 -1142 82742 -866
rect 82256 -1176 82742 -1142
<< nsubdiff >>
rect 3246 28520 3742 28554
rect 3246 28244 3280 28520
rect 3708 28458 3742 28520
rect 3708 28244 3742 28300
rect 3246 28204 3742 28244
rect 3246 27928 3280 28204
rect 3708 28148 3742 28204
rect 3708 27928 3742 27990
rect 3246 27894 3742 27928
rect 8236 28520 8732 28554
rect 8236 28244 8270 28520
rect 8698 28458 8732 28520
rect 8698 28244 8732 28300
rect 8236 28204 8732 28244
rect 8236 27928 8270 28204
rect 8698 28148 8732 28204
rect 8698 27928 8732 27990
rect 8236 27894 8732 27928
rect 13226 28520 13722 28554
rect 13226 28244 13260 28520
rect 13688 28458 13722 28520
rect 13688 28244 13722 28300
rect 13226 28204 13722 28244
rect 13226 27928 13260 28204
rect 13688 28148 13722 28204
rect 13688 27928 13722 27990
rect 13226 27894 13722 27928
rect 18216 28520 18712 28554
rect 18216 28244 18250 28520
rect 18678 28458 18712 28520
rect 18678 28244 18712 28300
rect 18216 28204 18712 28244
rect 18216 27928 18250 28204
rect 18678 28148 18712 28204
rect 18678 27928 18712 27990
rect 18216 27894 18712 27928
rect 23206 28520 23702 28554
rect 23206 28244 23240 28520
rect 23668 28458 23702 28520
rect 23668 28244 23702 28300
rect 23206 28204 23702 28244
rect 23206 27928 23240 28204
rect 23668 28148 23702 28204
rect 23668 27928 23702 27990
rect 23206 27894 23702 27928
rect 28196 28520 28692 28554
rect 28196 28244 28230 28520
rect 28658 28458 28692 28520
rect 28658 28244 28692 28300
rect 28196 28204 28692 28244
rect 28196 27928 28230 28204
rect 28658 28148 28692 28204
rect 28658 27928 28692 27990
rect 28196 27894 28692 27928
rect 33186 28520 33682 28554
rect 33186 28244 33220 28520
rect 33648 28458 33682 28520
rect 33648 28244 33682 28300
rect 33186 28204 33682 28244
rect 33186 27928 33220 28204
rect 33648 28148 33682 28204
rect 33648 27928 33682 27990
rect 33186 27894 33682 27928
rect 38176 28520 38672 28554
rect 38176 28244 38210 28520
rect 38638 28458 38672 28520
rect 38638 28244 38672 28300
rect 38176 28204 38672 28244
rect 38176 27928 38210 28204
rect 38638 28148 38672 28204
rect 38638 27928 38672 27990
rect 38176 27894 38672 27928
rect 43166 28520 43662 28554
rect 43166 28244 43200 28520
rect 43628 28458 43662 28520
rect 43628 28244 43662 28300
rect 43166 28204 43662 28244
rect 43166 27928 43200 28204
rect 43628 28148 43662 28204
rect 43628 27928 43662 27990
rect 43166 27894 43662 27928
rect 48156 28520 48652 28554
rect 48156 28244 48190 28520
rect 48618 28458 48652 28520
rect 48618 28244 48652 28300
rect 48156 28204 48652 28244
rect 48156 27928 48190 28204
rect 48618 28148 48652 28204
rect 48618 27928 48652 27990
rect 48156 27894 48652 27928
rect 53146 28520 53642 28554
rect 53146 28244 53180 28520
rect 53608 28458 53642 28520
rect 53608 28244 53642 28300
rect 53146 28204 53642 28244
rect 53146 27928 53180 28204
rect 53608 28148 53642 28204
rect 53608 27928 53642 27990
rect 53146 27894 53642 27928
rect 58136 28520 58632 28554
rect 58136 28244 58170 28520
rect 58598 28458 58632 28520
rect 58598 28244 58632 28300
rect 58136 28204 58632 28244
rect 58136 27928 58170 28204
rect 58598 28148 58632 28204
rect 58598 27928 58632 27990
rect 58136 27894 58632 27928
rect 63126 28520 63622 28554
rect 63126 28244 63160 28520
rect 63588 28458 63622 28520
rect 63588 28244 63622 28300
rect 63126 28204 63622 28244
rect 63126 27928 63160 28204
rect 63588 28148 63622 28204
rect 63588 27928 63622 27990
rect 63126 27894 63622 27928
rect 68116 28520 68612 28554
rect 68116 28244 68150 28520
rect 68578 28458 68612 28520
rect 68578 28244 68612 28300
rect 68116 28204 68612 28244
rect 68116 27928 68150 28204
rect 68578 28148 68612 28204
rect 68578 27928 68612 27990
rect 68116 27894 68612 27928
rect 73106 28520 73602 28554
rect 73106 28244 73140 28520
rect 73568 28458 73602 28520
rect 73568 28244 73602 28300
rect 73106 28204 73602 28244
rect 73106 27928 73140 28204
rect 73568 28148 73602 28204
rect 73568 27928 73602 27990
rect 73106 27894 73602 27928
rect 78096 28520 78592 28554
rect 78096 28244 78130 28520
rect 78558 28458 78592 28520
rect 78558 28244 78592 28300
rect 78096 28204 78592 28244
rect 78096 27928 78130 28204
rect 78558 28148 78592 28204
rect 78558 27928 78592 27990
rect 78096 27894 78592 27928
rect 82816 28520 83312 28554
rect 82816 28244 82850 28520
rect 83278 28458 83312 28520
rect 83278 28244 83312 28300
rect 82816 28204 83312 28244
rect 82816 27928 82850 28204
rect 83278 28148 83312 28204
rect 83278 27928 83312 27990
rect 82816 27894 83312 27928
rect 82816 26810 83312 26844
rect 82816 26534 82850 26810
rect 83278 26748 83312 26810
rect 83278 26534 83312 26590
rect 82816 26494 83312 26534
rect 82816 26218 82850 26494
rect 83278 26438 83312 26494
rect 83278 26218 83312 26280
rect 82816 26184 83312 26218
rect 82816 25100 83312 25134
rect 82816 24824 82850 25100
rect 83278 25038 83312 25100
rect 83278 24824 83312 24880
rect 82816 24784 83312 24824
rect 82816 24508 82850 24784
rect 83278 24728 83312 24784
rect 83278 24508 83312 24570
rect 82816 24474 83312 24508
rect -1474 23390 -978 23424
rect -1474 23114 -1440 23390
rect -1012 23328 -978 23390
rect -1012 23114 -978 23170
rect -1474 23074 -978 23114
rect -1474 22798 -1440 23074
rect -1012 23018 -978 23074
rect -1012 22798 -978 22860
rect -1474 22764 -978 22798
rect 82816 23390 83312 23424
rect 82816 23114 82850 23390
rect 83278 23328 83312 23390
rect 83278 23114 83312 23170
rect 82816 23074 83312 23114
rect 82816 22798 82850 23074
rect 83278 23018 83312 23074
rect 83278 22798 83312 22860
rect 82816 22764 83312 22798
rect -1474 21680 -978 21714
rect -1474 21404 -1440 21680
rect -1012 21618 -978 21680
rect -1012 21404 -978 21460
rect -1474 21364 -978 21404
rect -1474 21088 -1440 21364
rect -1012 21308 -978 21364
rect -1012 21088 -978 21150
rect -1474 21054 -978 21088
rect 82816 21680 83312 21714
rect 82816 21404 82850 21680
rect 83278 21618 83312 21680
rect 83278 21404 83312 21460
rect 82816 21364 83312 21404
rect 82816 21088 82850 21364
rect 83278 21308 83312 21364
rect 83278 21088 83312 21150
rect 82816 21054 83312 21088
rect -1474 19970 -978 20004
rect -1474 19694 -1440 19970
rect -1012 19908 -978 19970
rect -1012 19694 -978 19750
rect -1474 19654 -978 19694
rect -1474 19378 -1440 19654
rect -1012 19598 -978 19654
rect -1012 19378 -978 19440
rect -1474 19344 -978 19378
rect 82816 19970 83312 20004
rect 82816 19694 82850 19970
rect 83278 19908 83312 19970
rect 83278 19694 83312 19750
rect 82816 19654 83312 19694
rect 82816 19378 82850 19654
rect 83278 19598 83312 19654
rect 83278 19378 83312 19440
rect 82816 19344 83312 19378
rect -1474 18260 -978 18294
rect -1474 17984 -1440 18260
rect -1012 18198 -978 18260
rect -1012 17984 -978 18040
rect -1474 17944 -978 17984
rect -1474 17668 -1440 17944
rect -1012 17888 -978 17944
rect -1012 17668 -978 17730
rect -1474 17634 -978 17668
rect 82816 18260 83312 18294
rect 82816 17984 82850 18260
rect 83278 18198 83312 18260
rect 83278 17984 83312 18040
rect 82816 17944 83312 17984
rect 82816 17668 82850 17944
rect 83278 17888 83312 17944
rect 83278 17668 83312 17730
rect 82816 17634 83312 17668
rect -1474 16550 -978 16584
rect -1474 16274 -1440 16550
rect -1012 16488 -978 16550
rect -1012 16274 -978 16330
rect -1474 16234 -978 16274
rect -1474 15958 -1440 16234
rect -1012 16178 -978 16234
rect -1012 15958 -978 16020
rect -1474 15924 -978 15958
rect 82816 16550 83312 16584
rect 82816 16274 82850 16550
rect 83278 16488 83312 16550
rect 83278 16274 83312 16330
rect 82816 16234 83312 16274
rect 82816 15958 82850 16234
rect 83278 16178 83312 16234
rect 83278 15958 83312 16020
rect 82816 15924 83312 15958
rect -1474 14840 -978 14874
rect -1474 14564 -1440 14840
rect -1012 14778 -978 14840
rect -1012 14564 -978 14620
rect -1474 14524 -978 14564
rect -1474 14248 -1440 14524
rect -1012 14468 -978 14524
rect -1012 14248 -978 14310
rect -1474 14214 -978 14248
rect 82816 14840 83312 14874
rect 82816 14564 82850 14840
rect 83278 14778 83312 14840
rect 83278 14564 83312 14620
rect 82816 14524 83312 14564
rect 82816 14248 82850 14524
rect 83278 14468 83312 14524
rect 83278 14248 83312 14310
rect 82816 14214 83312 14248
rect -1474 13130 -978 13164
rect -1474 12854 -1440 13130
rect -1012 13068 -978 13130
rect -1012 12854 -978 12910
rect -1474 12814 -978 12854
rect -1474 12538 -1440 12814
rect -1012 12758 -978 12814
rect -1012 12538 -978 12600
rect -1474 12504 -978 12538
rect 82816 13130 83312 13164
rect 82816 12854 82850 13130
rect 83278 13068 83312 13130
rect 83278 12854 83312 12910
rect 82816 12814 83312 12854
rect 82816 12538 82850 12814
rect 83278 12758 83312 12814
rect 83278 12538 83312 12600
rect 82816 12504 83312 12538
rect -1474 11420 -978 11454
rect -1474 11144 -1440 11420
rect -1012 11358 -978 11420
rect -1012 11144 -978 11200
rect -1474 11104 -978 11144
rect -1474 10828 -1440 11104
rect -1012 11048 -978 11104
rect -1012 10828 -978 10890
rect -1474 10794 -978 10828
rect 82816 11420 83312 11454
rect 82816 11144 82850 11420
rect 83278 11358 83312 11420
rect 83278 11144 83312 11200
rect 82816 11104 83312 11144
rect 82816 10828 82850 11104
rect 83278 11048 83312 11104
rect 83278 10828 83312 10890
rect 82816 10794 83312 10828
rect -1474 9710 -978 9744
rect -1474 9434 -1440 9710
rect -1012 9648 -978 9710
rect -1012 9434 -978 9490
rect -1474 9394 -978 9434
rect -1474 9118 -1440 9394
rect -1012 9338 -978 9394
rect -1012 9118 -978 9180
rect -1474 9084 -978 9118
rect 82816 9710 83312 9744
rect 82816 9434 82850 9710
rect 83278 9648 83312 9710
rect 83278 9434 83312 9490
rect 82816 9394 83312 9434
rect 82816 9118 82850 9394
rect 83278 9338 83312 9394
rect 83278 9118 83312 9180
rect 82816 9084 83312 9118
rect -1474 8000 -978 8034
rect -1474 7724 -1440 8000
rect -1012 7938 -978 8000
rect -1012 7724 -978 7780
rect -1474 7684 -978 7724
rect -1474 7408 -1440 7684
rect -1012 7628 -978 7684
rect -1012 7408 -978 7470
rect -1474 7374 -978 7408
rect 82816 8000 83312 8034
rect 82816 7724 82850 8000
rect 83278 7938 83312 8000
rect 83278 7724 83312 7780
rect 82816 7684 83312 7724
rect 82816 7408 82850 7684
rect 83278 7628 83312 7684
rect 83278 7408 83312 7470
rect 82816 7374 83312 7408
rect -1474 6290 -978 6324
rect -1474 6014 -1440 6290
rect -1012 6228 -978 6290
rect -1012 6014 -978 6070
rect -1474 5974 -978 6014
rect -1474 5698 -1440 5974
rect -1012 5918 -978 5974
rect -1012 5698 -978 5760
rect -1474 5664 -978 5698
rect 82816 6290 83312 6324
rect 82816 6014 82850 6290
rect 83278 6228 83312 6290
rect 83278 6014 83312 6070
rect 82816 5974 83312 6014
rect 82816 5698 82850 5974
rect 83278 5918 83312 5974
rect 83278 5698 83312 5760
rect 82816 5664 83312 5698
rect -1474 4580 -978 4614
rect -1474 4304 -1440 4580
rect -1012 4518 -978 4580
rect -1012 4304 -978 4360
rect -1474 4264 -978 4304
rect -1474 3988 -1440 4264
rect -1012 4208 -978 4264
rect -1012 3988 -978 4050
rect -1474 3954 -978 3988
rect 82816 4580 83312 4614
rect 82816 4304 82850 4580
rect 83278 4518 83312 4580
rect 83278 4304 83312 4360
rect 82816 4264 83312 4304
rect 82816 3988 82850 4264
rect 83278 4208 83312 4264
rect 83278 3988 83312 4050
rect 82816 3954 83312 3988
rect -1474 2870 -978 2904
rect -1474 2594 -1440 2870
rect -1012 2808 -978 2870
rect -1012 2594 -978 2650
rect -1474 2554 -978 2594
rect -1474 2278 -1440 2554
rect -1012 2498 -978 2554
rect -1012 2278 -978 2340
rect -1474 2244 -978 2278
rect 82816 2870 83312 2904
rect 82816 2594 82850 2870
rect 83278 2808 83312 2870
rect 83278 2594 83312 2650
rect 82816 2554 83312 2594
rect 82816 2278 82850 2554
rect 83278 2498 83312 2554
rect 83278 2278 83312 2340
rect 82816 2244 83312 2278
rect -1474 1160 -978 1194
rect -1474 884 -1440 1160
rect -1012 1098 -978 1160
rect -1012 884 -978 940
rect -1474 844 -978 884
rect -1474 568 -1440 844
rect -1012 788 -978 844
rect -1012 568 -978 630
rect -1474 534 -978 568
rect 82816 1160 83312 1194
rect 82816 884 82850 1160
rect 83278 1098 83312 1160
rect 83278 884 83312 940
rect 82816 844 83312 884
rect 82816 568 82850 844
rect 83278 788 83312 844
rect 83278 568 83312 630
rect 82816 534 83312 568
rect -1474 -550 -978 -516
rect -1474 -826 -1440 -550
rect -1012 -612 -978 -550
rect -1012 -826 -978 -770
rect -1474 -866 -978 -826
rect -1474 -1142 -1440 -866
rect -1012 -922 -978 -866
rect -1012 -1142 -978 -1080
rect -1474 -1176 -978 -1142
rect 3246 -550 3742 -516
rect 3246 -826 3280 -550
rect 3708 -612 3742 -550
rect 3708 -826 3742 -770
rect 3246 -866 3742 -826
rect 3246 -1142 3280 -866
rect 3708 -922 3742 -866
rect 3708 -1142 3742 -1080
rect 3246 -1176 3742 -1142
rect 8236 -550 8732 -516
rect 8236 -826 8270 -550
rect 8698 -612 8732 -550
rect 8698 -826 8732 -770
rect 8236 -866 8732 -826
rect 8236 -1142 8270 -866
rect 8698 -922 8732 -866
rect 8698 -1142 8732 -1080
rect 8236 -1176 8732 -1142
rect 13226 -550 13722 -516
rect 13226 -826 13260 -550
rect 13688 -612 13722 -550
rect 13688 -826 13722 -770
rect 13226 -866 13722 -826
rect 13226 -1142 13260 -866
rect 13688 -922 13722 -866
rect 13688 -1142 13722 -1080
rect 13226 -1176 13722 -1142
rect 18216 -550 18712 -516
rect 18216 -826 18250 -550
rect 18678 -612 18712 -550
rect 18678 -826 18712 -770
rect 18216 -866 18712 -826
rect 18216 -1142 18250 -866
rect 18678 -922 18712 -866
rect 18678 -1142 18712 -1080
rect 18216 -1176 18712 -1142
rect 23206 -550 23702 -516
rect 23206 -826 23240 -550
rect 23668 -612 23702 -550
rect 23668 -826 23702 -770
rect 23206 -866 23702 -826
rect 23206 -1142 23240 -866
rect 23668 -922 23702 -866
rect 23668 -1142 23702 -1080
rect 23206 -1176 23702 -1142
rect 28196 -550 28692 -516
rect 28196 -826 28230 -550
rect 28658 -612 28692 -550
rect 28658 -826 28692 -770
rect 28196 -866 28692 -826
rect 28196 -1142 28230 -866
rect 28658 -922 28692 -866
rect 28658 -1142 28692 -1080
rect 28196 -1176 28692 -1142
rect 33186 -550 33682 -516
rect 33186 -826 33220 -550
rect 33648 -612 33682 -550
rect 33648 -826 33682 -770
rect 33186 -866 33682 -826
rect 33186 -1142 33220 -866
rect 33648 -922 33682 -866
rect 33648 -1142 33682 -1080
rect 33186 -1176 33682 -1142
rect 38176 -550 38672 -516
rect 38176 -826 38210 -550
rect 38638 -612 38672 -550
rect 38638 -826 38672 -770
rect 38176 -866 38672 -826
rect 38176 -1142 38210 -866
rect 38638 -922 38672 -866
rect 38638 -1142 38672 -1080
rect 38176 -1176 38672 -1142
rect 43166 -550 43662 -516
rect 43166 -826 43200 -550
rect 43628 -612 43662 -550
rect 43628 -826 43662 -770
rect 43166 -866 43662 -826
rect 43166 -1142 43200 -866
rect 43628 -922 43662 -866
rect 43628 -1142 43662 -1080
rect 43166 -1176 43662 -1142
rect 48156 -550 48652 -516
rect 48156 -826 48190 -550
rect 48618 -612 48652 -550
rect 48618 -826 48652 -770
rect 48156 -866 48652 -826
rect 48156 -1142 48190 -866
rect 48618 -922 48652 -866
rect 48618 -1142 48652 -1080
rect 48156 -1176 48652 -1142
rect 53146 -550 53642 -516
rect 53146 -826 53180 -550
rect 53608 -612 53642 -550
rect 53608 -826 53642 -770
rect 53146 -866 53642 -826
rect 53146 -1142 53180 -866
rect 53608 -922 53642 -866
rect 53608 -1142 53642 -1080
rect 53146 -1176 53642 -1142
rect 58136 -550 58632 -516
rect 58136 -826 58170 -550
rect 58598 -612 58632 -550
rect 58598 -826 58632 -770
rect 58136 -866 58632 -826
rect 58136 -1142 58170 -866
rect 58598 -922 58632 -866
rect 58598 -1142 58632 -1080
rect 58136 -1176 58632 -1142
rect 63126 -550 63622 -516
rect 63126 -826 63160 -550
rect 63588 -612 63622 -550
rect 63588 -826 63622 -770
rect 63126 -866 63622 -826
rect 63126 -1142 63160 -866
rect 63588 -922 63622 -866
rect 63588 -1142 63622 -1080
rect 63126 -1176 63622 -1142
rect 68116 -550 68612 -516
rect 68116 -826 68150 -550
rect 68578 -612 68612 -550
rect 68578 -826 68612 -770
rect 68116 -866 68612 -826
rect 68116 -1142 68150 -866
rect 68578 -922 68612 -866
rect 68578 -1142 68612 -1080
rect 68116 -1176 68612 -1142
rect 73106 -550 73602 -516
rect 73106 -826 73140 -550
rect 73568 -612 73602 -550
rect 73568 -826 73602 -770
rect 73106 -866 73602 -826
rect 73106 -1142 73140 -866
rect 73568 -922 73602 -866
rect 73568 -1142 73602 -1080
rect 73106 -1176 73602 -1142
rect 78096 -550 78592 -516
rect 78096 -826 78130 -550
rect 78558 -612 78592 -550
rect 78558 -826 78592 -770
rect 78096 -866 78592 -826
rect 78096 -1142 78130 -866
rect 78558 -922 78592 -866
rect 78558 -1142 78592 -1080
rect 78096 -1176 78592 -1142
rect 82816 -550 83312 -516
rect 82816 -826 82850 -550
rect 83278 -612 83312 -550
rect 83278 -826 83312 -770
rect 82816 -866 83312 -826
rect 82816 -1142 82850 -866
rect 83278 -922 83312 -866
rect 83278 -1142 83312 -1080
rect 82816 -1176 83312 -1142
<< psubdiffcont >>
rect 2686 28300 2720 28458
rect 2686 27990 2720 28148
rect 7676 28300 7710 28458
rect 7676 27990 7710 28148
rect 12666 28300 12700 28458
rect 12666 27990 12700 28148
rect 17656 28300 17690 28458
rect 17656 27990 17690 28148
rect 22646 28300 22680 28458
rect 22646 27990 22680 28148
rect 27636 28300 27670 28458
rect 27636 27990 27670 28148
rect 32626 28300 32660 28458
rect 32626 27990 32660 28148
rect 37616 28300 37650 28458
rect 37616 27990 37650 28148
rect 42606 28300 42640 28458
rect 42606 27990 42640 28148
rect 47596 28300 47630 28458
rect 47596 27990 47630 28148
rect 52586 28300 52620 28458
rect 52586 27990 52620 28148
rect 57576 28300 57610 28458
rect 57576 27990 57610 28148
rect 62566 28300 62600 28458
rect 62566 27990 62600 28148
rect 67556 28300 67590 28458
rect 67556 27990 67590 28148
rect 72546 28300 72580 28458
rect 72546 27990 72580 28148
rect 77536 28300 77570 28458
rect 77536 27990 77570 28148
rect 82256 28300 82290 28458
rect 82256 27990 82290 28148
rect 82256 26590 82290 26748
rect 82256 26280 82290 26438
rect 82256 24880 82290 25038
rect 82256 24570 82290 24728
rect -2034 23170 -2000 23328
rect -2034 22860 -2000 23018
rect 82256 23170 82290 23328
rect 82256 22860 82290 23018
rect -2034 21460 -2000 21618
rect -2034 21150 -2000 21308
rect 82256 21460 82290 21618
rect 82256 21150 82290 21308
rect -2034 19750 -2000 19908
rect -2034 19440 -2000 19598
rect 82256 19750 82290 19908
rect 82256 19440 82290 19598
rect -2034 18040 -2000 18198
rect -2034 17730 -2000 17888
rect 82256 18040 82290 18198
rect 82256 17730 82290 17888
rect -2034 16330 -2000 16488
rect -2034 16020 -2000 16178
rect 82256 16330 82290 16488
rect 82256 16020 82290 16178
rect -2034 14620 -2000 14778
rect -2034 14310 -2000 14468
rect 82256 14620 82290 14778
rect 82256 14310 82290 14468
rect -2034 12910 -2000 13068
rect -2034 12600 -2000 12758
rect 82256 12910 82290 13068
rect 82256 12600 82290 12758
rect -2034 11200 -2000 11358
rect -2034 10890 -2000 11048
rect 82256 11200 82290 11358
rect 82256 10890 82290 11048
rect -2034 9490 -2000 9648
rect -2034 9180 -2000 9338
rect 82256 9490 82290 9648
rect 82256 9180 82290 9338
rect -2034 7780 -2000 7938
rect -2034 7470 -2000 7628
rect 82256 7780 82290 7938
rect 82256 7470 82290 7628
rect -2034 6070 -2000 6228
rect -2034 5760 -2000 5918
rect 82256 6070 82290 6228
rect 82256 5760 82290 5918
rect -2034 4360 -2000 4518
rect -2034 4050 -2000 4208
rect 82256 4360 82290 4518
rect 82256 4050 82290 4208
rect -2034 2650 -2000 2808
rect -2034 2340 -2000 2498
rect 82256 2650 82290 2808
rect 82256 2340 82290 2498
rect -2034 940 -2000 1098
rect -2034 630 -2000 788
rect 82256 940 82290 1098
rect 82256 630 82290 788
rect -2034 -770 -2000 -612
rect -2034 -1080 -2000 -922
rect 2686 -770 2720 -612
rect 2686 -1080 2720 -922
rect 7676 -770 7710 -612
rect 7676 -1080 7710 -922
rect 12666 -770 12700 -612
rect 12666 -1080 12700 -922
rect 17656 -770 17690 -612
rect 17656 -1080 17690 -922
rect 22646 -770 22680 -612
rect 22646 -1080 22680 -922
rect 27636 -770 27670 -612
rect 27636 -1080 27670 -922
rect 32626 -770 32660 -612
rect 32626 -1080 32660 -922
rect 37616 -770 37650 -612
rect 37616 -1080 37650 -922
rect 42606 -770 42640 -612
rect 42606 -1080 42640 -922
rect 47596 -770 47630 -612
rect 47596 -1080 47630 -922
rect 52586 -770 52620 -612
rect 52586 -1080 52620 -922
rect 57576 -770 57610 -612
rect 57576 -1080 57610 -922
rect 62566 -770 62600 -612
rect 62566 -1080 62600 -922
rect 67556 -770 67590 -612
rect 67556 -1080 67590 -922
rect 72546 -770 72580 -612
rect 72546 -1080 72580 -922
rect 77536 -770 77570 -612
rect 77536 -1080 77570 -922
rect 82256 -770 82290 -612
rect 82256 -1080 82290 -922
<< nsubdiffcont >>
rect 3708 28300 3742 28458
rect 3708 27990 3742 28148
rect 8698 28300 8732 28458
rect 8698 27990 8732 28148
rect 13688 28300 13722 28458
rect 13688 27990 13722 28148
rect 18678 28300 18712 28458
rect 18678 27990 18712 28148
rect 23668 28300 23702 28458
rect 23668 27990 23702 28148
rect 28658 28300 28692 28458
rect 28658 27990 28692 28148
rect 33648 28300 33682 28458
rect 33648 27990 33682 28148
rect 38638 28300 38672 28458
rect 38638 27990 38672 28148
rect 43628 28300 43662 28458
rect 43628 27990 43662 28148
rect 48618 28300 48652 28458
rect 48618 27990 48652 28148
rect 53608 28300 53642 28458
rect 53608 27990 53642 28148
rect 58598 28300 58632 28458
rect 58598 27990 58632 28148
rect 63588 28300 63622 28458
rect 63588 27990 63622 28148
rect 68578 28300 68612 28458
rect 68578 27990 68612 28148
rect 73568 28300 73602 28458
rect 73568 27990 73602 28148
rect 78558 28300 78592 28458
rect 78558 27990 78592 28148
rect 83278 28300 83312 28458
rect 83278 27990 83312 28148
rect 83278 26590 83312 26748
rect 83278 26280 83312 26438
rect 83278 24880 83312 25038
rect 83278 24570 83312 24728
rect -1012 23170 -978 23328
rect -1012 22860 -978 23018
rect 83278 23170 83312 23328
rect 83278 22860 83312 23018
rect -1012 21460 -978 21618
rect -1012 21150 -978 21308
rect 83278 21460 83312 21618
rect 83278 21150 83312 21308
rect -1012 19750 -978 19908
rect -1012 19440 -978 19598
rect 83278 19750 83312 19908
rect 83278 19440 83312 19598
rect -1012 18040 -978 18198
rect -1012 17730 -978 17888
rect 83278 18040 83312 18198
rect 83278 17730 83312 17888
rect -1012 16330 -978 16488
rect -1012 16020 -978 16178
rect 83278 16330 83312 16488
rect 83278 16020 83312 16178
rect -1012 14620 -978 14778
rect -1012 14310 -978 14468
rect 83278 14620 83312 14778
rect 83278 14310 83312 14468
rect -1012 12910 -978 13068
rect -1012 12600 -978 12758
rect 83278 12910 83312 13068
rect 83278 12600 83312 12758
rect -1012 11200 -978 11358
rect -1012 10890 -978 11048
rect 83278 11200 83312 11358
rect 83278 10890 83312 11048
rect -1012 9490 -978 9648
rect -1012 9180 -978 9338
rect 83278 9490 83312 9648
rect 83278 9180 83312 9338
rect -1012 7780 -978 7938
rect -1012 7470 -978 7628
rect 83278 7780 83312 7938
rect 83278 7470 83312 7628
rect -1012 6070 -978 6228
rect -1012 5760 -978 5918
rect 83278 6070 83312 6228
rect 83278 5760 83312 5918
rect -1012 4360 -978 4518
rect -1012 4050 -978 4208
rect 83278 4360 83312 4518
rect 83278 4050 83312 4208
rect -1012 2650 -978 2808
rect -1012 2340 -978 2498
rect 83278 2650 83312 2808
rect 83278 2340 83312 2498
rect -1012 940 -978 1098
rect -1012 630 -978 788
rect 83278 940 83312 1098
rect 83278 630 83312 788
rect -1012 -770 -978 -612
rect -1012 -1080 -978 -922
rect 3708 -770 3742 -612
rect 3708 -1080 3742 -922
rect 8698 -770 8732 -612
rect 8698 -1080 8732 -922
rect 13688 -770 13722 -612
rect 13688 -1080 13722 -922
rect 18678 -770 18712 -612
rect 18678 -1080 18712 -922
rect 23668 -770 23702 -612
rect 23668 -1080 23702 -922
rect 28658 -770 28692 -612
rect 28658 -1080 28692 -922
rect 33648 -770 33682 -612
rect 33648 -1080 33682 -922
rect 38638 -770 38672 -612
rect 38638 -1080 38672 -922
rect 43628 -770 43662 -612
rect 43628 -1080 43662 -922
rect 48618 -770 48652 -612
rect 48618 -1080 48652 -922
rect 53608 -770 53642 -612
rect 53608 -1080 53642 -922
rect 58598 -770 58632 -612
rect 58598 -1080 58632 -922
rect 63588 -770 63622 -612
rect 63588 -1080 63622 -922
rect 68578 -770 68612 -612
rect 68578 -1080 68612 -922
rect 73568 -770 73602 -612
rect 73568 -1080 73602 -922
rect 78558 -770 78592 -612
rect 78558 -1080 78592 -922
rect 83278 -770 83312 -612
rect 83278 -1080 83312 -922
<< poly >>
rect 2772 28396 2838 28412
rect 2772 28362 2788 28396
rect 2822 28394 2838 28396
rect 2822 28364 2860 28394
rect 3060 28364 3086 28394
rect 2822 28362 2838 28364
rect 2772 28346 2838 28362
rect 2772 28086 2838 28102
rect 2772 28052 2788 28086
rect 2822 28084 2838 28086
rect 2822 28054 2860 28084
rect 3060 28054 3086 28084
rect 2822 28052 2838 28054
rect 2772 28036 2838 28052
rect 3589 28396 3655 28412
rect 3589 28394 3605 28396
rect 3332 28364 3358 28394
rect 3558 28364 3605 28394
rect 3589 28362 3605 28364
rect 3639 28362 3655 28396
rect 3589 28346 3655 28362
rect 3589 28086 3655 28102
rect 3589 28084 3605 28086
rect 3332 28054 3358 28084
rect 3558 28054 3605 28084
rect 3589 28052 3605 28054
rect 3639 28052 3655 28086
rect 3589 28036 3655 28052
rect 7762 28396 7828 28412
rect 7762 28362 7778 28396
rect 7812 28394 7828 28396
rect 7812 28364 7850 28394
rect 8050 28364 8076 28394
rect 7812 28362 7828 28364
rect 7762 28346 7828 28362
rect 7762 28086 7828 28102
rect 7762 28052 7778 28086
rect 7812 28084 7828 28086
rect 7812 28054 7850 28084
rect 8050 28054 8076 28084
rect 7812 28052 7828 28054
rect 7762 28036 7828 28052
rect 8579 28396 8645 28412
rect 8579 28394 8595 28396
rect 8322 28364 8348 28394
rect 8548 28364 8595 28394
rect 8579 28362 8595 28364
rect 8629 28362 8645 28396
rect 8579 28346 8645 28362
rect 8579 28086 8645 28102
rect 8579 28084 8595 28086
rect 8322 28054 8348 28084
rect 8548 28054 8595 28084
rect 8579 28052 8595 28054
rect 8629 28052 8645 28086
rect 8579 28036 8645 28052
rect 12752 28396 12818 28412
rect 12752 28362 12768 28396
rect 12802 28394 12818 28396
rect 12802 28364 12840 28394
rect 13040 28364 13066 28394
rect 12802 28362 12818 28364
rect 12752 28346 12818 28362
rect 12752 28086 12818 28102
rect 12752 28052 12768 28086
rect 12802 28084 12818 28086
rect 12802 28054 12840 28084
rect 13040 28054 13066 28084
rect 12802 28052 12818 28054
rect 12752 28036 12818 28052
rect 13569 28396 13635 28412
rect 13569 28394 13585 28396
rect 13312 28364 13338 28394
rect 13538 28364 13585 28394
rect 13569 28362 13585 28364
rect 13619 28362 13635 28396
rect 13569 28346 13635 28362
rect 13569 28086 13635 28102
rect 13569 28084 13585 28086
rect 13312 28054 13338 28084
rect 13538 28054 13585 28084
rect 13569 28052 13585 28054
rect 13619 28052 13635 28086
rect 13569 28036 13635 28052
rect 17742 28396 17808 28412
rect 17742 28362 17758 28396
rect 17792 28394 17808 28396
rect 17792 28364 17830 28394
rect 18030 28364 18056 28394
rect 17792 28362 17808 28364
rect 17742 28346 17808 28362
rect 17742 28086 17808 28102
rect 17742 28052 17758 28086
rect 17792 28084 17808 28086
rect 17792 28054 17830 28084
rect 18030 28054 18056 28084
rect 17792 28052 17808 28054
rect 17742 28036 17808 28052
rect 18559 28396 18625 28412
rect 18559 28394 18575 28396
rect 18302 28364 18328 28394
rect 18528 28364 18575 28394
rect 18559 28362 18575 28364
rect 18609 28362 18625 28396
rect 18559 28346 18625 28362
rect 18559 28086 18625 28102
rect 18559 28084 18575 28086
rect 18302 28054 18328 28084
rect 18528 28054 18575 28084
rect 18559 28052 18575 28054
rect 18609 28052 18625 28086
rect 18559 28036 18625 28052
rect 22732 28396 22798 28412
rect 22732 28362 22748 28396
rect 22782 28394 22798 28396
rect 22782 28364 22820 28394
rect 23020 28364 23046 28394
rect 22782 28362 22798 28364
rect 22732 28346 22798 28362
rect 22732 28086 22798 28102
rect 22732 28052 22748 28086
rect 22782 28084 22798 28086
rect 22782 28054 22820 28084
rect 23020 28054 23046 28084
rect 22782 28052 22798 28054
rect 22732 28036 22798 28052
rect 23549 28396 23615 28412
rect 23549 28394 23565 28396
rect 23292 28364 23318 28394
rect 23518 28364 23565 28394
rect 23549 28362 23565 28364
rect 23599 28362 23615 28396
rect 23549 28346 23615 28362
rect 23549 28086 23615 28102
rect 23549 28084 23565 28086
rect 23292 28054 23318 28084
rect 23518 28054 23565 28084
rect 23549 28052 23565 28054
rect 23599 28052 23615 28086
rect 23549 28036 23615 28052
rect 27722 28396 27788 28412
rect 27722 28362 27738 28396
rect 27772 28394 27788 28396
rect 27772 28364 27810 28394
rect 28010 28364 28036 28394
rect 27772 28362 27788 28364
rect 27722 28346 27788 28362
rect 27722 28086 27788 28102
rect 27722 28052 27738 28086
rect 27772 28084 27788 28086
rect 27772 28054 27810 28084
rect 28010 28054 28036 28084
rect 27772 28052 27788 28054
rect 27722 28036 27788 28052
rect 28539 28396 28605 28412
rect 28539 28394 28555 28396
rect 28282 28364 28308 28394
rect 28508 28364 28555 28394
rect 28539 28362 28555 28364
rect 28589 28362 28605 28396
rect 28539 28346 28605 28362
rect 28539 28086 28605 28102
rect 28539 28084 28555 28086
rect 28282 28054 28308 28084
rect 28508 28054 28555 28084
rect 28539 28052 28555 28054
rect 28589 28052 28605 28086
rect 28539 28036 28605 28052
rect 32712 28396 32778 28412
rect 32712 28362 32728 28396
rect 32762 28394 32778 28396
rect 32762 28364 32800 28394
rect 33000 28364 33026 28394
rect 32762 28362 32778 28364
rect 32712 28346 32778 28362
rect 32712 28086 32778 28102
rect 32712 28052 32728 28086
rect 32762 28084 32778 28086
rect 32762 28054 32800 28084
rect 33000 28054 33026 28084
rect 32762 28052 32778 28054
rect 32712 28036 32778 28052
rect 33529 28396 33595 28412
rect 33529 28394 33545 28396
rect 33272 28364 33298 28394
rect 33498 28364 33545 28394
rect 33529 28362 33545 28364
rect 33579 28362 33595 28396
rect 33529 28346 33595 28362
rect 33529 28086 33595 28102
rect 33529 28084 33545 28086
rect 33272 28054 33298 28084
rect 33498 28054 33545 28084
rect 33529 28052 33545 28054
rect 33579 28052 33595 28086
rect 33529 28036 33595 28052
rect 37702 28396 37768 28412
rect 37702 28362 37718 28396
rect 37752 28394 37768 28396
rect 37752 28364 37790 28394
rect 37990 28364 38016 28394
rect 37752 28362 37768 28364
rect 37702 28346 37768 28362
rect 37702 28086 37768 28102
rect 37702 28052 37718 28086
rect 37752 28084 37768 28086
rect 37752 28054 37790 28084
rect 37990 28054 38016 28084
rect 37752 28052 37768 28054
rect 37702 28036 37768 28052
rect 38519 28396 38585 28412
rect 38519 28394 38535 28396
rect 38262 28364 38288 28394
rect 38488 28364 38535 28394
rect 38519 28362 38535 28364
rect 38569 28362 38585 28396
rect 38519 28346 38585 28362
rect 38519 28086 38585 28102
rect 38519 28084 38535 28086
rect 38262 28054 38288 28084
rect 38488 28054 38535 28084
rect 38519 28052 38535 28054
rect 38569 28052 38585 28086
rect 38519 28036 38585 28052
rect 42692 28396 42758 28412
rect 42692 28362 42708 28396
rect 42742 28394 42758 28396
rect 42742 28364 42780 28394
rect 42980 28364 43006 28394
rect 42742 28362 42758 28364
rect 42692 28346 42758 28362
rect 42692 28086 42758 28102
rect 42692 28052 42708 28086
rect 42742 28084 42758 28086
rect 42742 28054 42780 28084
rect 42980 28054 43006 28084
rect 42742 28052 42758 28054
rect 42692 28036 42758 28052
rect 43509 28396 43575 28412
rect 43509 28394 43525 28396
rect 43252 28364 43278 28394
rect 43478 28364 43525 28394
rect 43509 28362 43525 28364
rect 43559 28362 43575 28396
rect 43509 28346 43575 28362
rect 43509 28086 43575 28102
rect 43509 28084 43525 28086
rect 43252 28054 43278 28084
rect 43478 28054 43525 28084
rect 43509 28052 43525 28054
rect 43559 28052 43575 28086
rect 43509 28036 43575 28052
rect 47682 28396 47748 28412
rect 47682 28362 47698 28396
rect 47732 28394 47748 28396
rect 47732 28364 47770 28394
rect 47970 28364 47996 28394
rect 47732 28362 47748 28364
rect 47682 28346 47748 28362
rect 47682 28086 47748 28102
rect 47682 28052 47698 28086
rect 47732 28084 47748 28086
rect 47732 28054 47770 28084
rect 47970 28054 47996 28084
rect 47732 28052 47748 28054
rect 47682 28036 47748 28052
rect 48499 28396 48565 28412
rect 48499 28394 48515 28396
rect 48242 28364 48268 28394
rect 48468 28364 48515 28394
rect 48499 28362 48515 28364
rect 48549 28362 48565 28396
rect 48499 28346 48565 28362
rect 48499 28086 48565 28102
rect 48499 28084 48515 28086
rect 48242 28054 48268 28084
rect 48468 28054 48515 28084
rect 48499 28052 48515 28054
rect 48549 28052 48565 28086
rect 48499 28036 48565 28052
rect 52672 28396 52738 28412
rect 52672 28362 52688 28396
rect 52722 28394 52738 28396
rect 52722 28364 52760 28394
rect 52960 28364 52986 28394
rect 52722 28362 52738 28364
rect 52672 28346 52738 28362
rect 52672 28086 52738 28102
rect 52672 28052 52688 28086
rect 52722 28084 52738 28086
rect 52722 28054 52760 28084
rect 52960 28054 52986 28084
rect 52722 28052 52738 28054
rect 52672 28036 52738 28052
rect 53489 28396 53555 28412
rect 53489 28394 53505 28396
rect 53232 28364 53258 28394
rect 53458 28364 53505 28394
rect 53489 28362 53505 28364
rect 53539 28362 53555 28396
rect 53489 28346 53555 28362
rect 53489 28086 53555 28102
rect 53489 28084 53505 28086
rect 53232 28054 53258 28084
rect 53458 28054 53505 28084
rect 53489 28052 53505 28054
rect 53539 28052 53555 28086
rect 53489 28036 53555 28052
rect 57662 28396 57728 28412
rect 57662 28362 57678 28396
rect 57712 28394 57728 28396
rect 57712 28364 57750 28394
rect 57950 28364 57976 28394
rect 57712 28362 57728 28364
rect 57662 28346 57728 28362
rect 57662 28086 57728 28102
rect 57662 28052 57678 28086
rect 57712 28084 57728 28086
rect 57712 28054 57750 28084
rect 57950 28054 57976 28084
rect 57712 28052 57728 28054
rect 57662 28036 57728 28052
rect 58479 28396 58545 28412
rect 58479 28394 58495 28396
rect 58222 28364 58248 28394
rect 58448 28364 58495 28394
rect 58479 28362 58495 28364
rect 58529 28362 58545 28396
rect 58479 28346 58545 28362
rect 58479 28086 58545 28102
rect 58479 28084 58495 28086
rect 58222 28054 58248 28084
rect 58448 28054 58495 28084
rect 58479 28052 58495 28054
rect 58529 28052 58545 28086
rect 58479 28036 58545 28052
rect 62652 28396 62718 28412
rect 62652 28362 62668 28396
rect 62702 28394 62718 28396
rect 62702 28364 62740 28394
rect 62940 28364 62966 28394
rect 62702 28362 62718 28364
rect 62652 28346 62718 28362
rect 62652 28086 62718 28102
rect 62652 28052 62668 28086
rect 62702 28084 62718 28086
rect 62702 28054 62740 28084
rect 62940 28054 62966 28084
rect 62702 28052 62718 28054
rect 62652 28036 62718 28052
rect 63469 28396 63535 28412
rect 63469 28394 63485 28396
rect 63212 28364 63238 28394
rect 63438 28364 63485 28394
rect 63469 28362 63485 28364
rect 63519 28362 63535 28396
rect 63469 28346 63535 28362
rect 63469 28086 63535 28102
rect 63469 28084 63485 28086
rect 63212 28054 63238 28084
rect 63438 28054 63485 28084
rect 63469 28052 63485 28054
rect 63519 28052 63535 28086
rect 63469 28036 63535 28052
rect 67642 28396 67708 28412
rect 67642 28362 67658 28396
rect 67692 28394 67708 28396
rect 67692 28364 67730 28394
rect 67930 28364 67956 28394
rect 67692 28362 67708 28364
rect 67642 28346 67708 28362
rect 67642 28086 67708 28102
rect 67642 28052 67658 28086
rect 67692 28084 67708 28086
rect 67692 28054 67730 28084
rect 67930 28054 67956 28084
rect 67692 28052 67708 28054
rect 67642 28036 67708 28052
rect 68459 28396 68525 28412
rect 68459 28394 68475 28396
rect 68202 28364 68228 28394
rect 68428 28364 68475 28394
rect 68459 28362 68475 28364
rect 68509 28362 68525 28396
rect 68459 28346 68525 28362
rect 68459 28086 68525 28102
rect 68459 28084 68475 28086
rect 68202 28054 68228 28084
rect 68428 28054 68475 28084
rect 68459 28052 68475 28054
rect 68509 28052 68525 28086
rect 68459 28036 68525 28052
rect 72632 28396 72698 28412
rect 72632 28362 72648 28396
rect 72682 28394 72698 28396
rect 72682 28364 72720 28394
rect 72920 28364 72946 28394
rect 72682 28362 72698 28364
rect 72632 28346 72698 28362
rect 72632 28086 72698 28102
rect 72632 28052 72648 28086
rect 72682 28084 72698 28086
rect 72682 28054 72720 28084
rect 72920 28054 72946 28084
rect 72682 28052 72698 28054
rect 72632 28036 72698 28052
rect 73449 28396 73515 28412
rect 73449 28394 73465 28396
rect 73192 28364 73218 28394
rect 73418 28364 73465 28394
rect 73449 28362 73465 28364
rect 73499 28362 73515 28396
rect 73449 28346 73515 28362
rect 73449 28086 73515 28102
rect 73449 28084 73465 28086
rect 73192 28054 73218 28084
rect 73418 28054 73465 28084
rect 73449 28052 73465 28054
rect 73499 28052 73515 28086
rect 73449 28036 73515 28052
rect 77622 28396 77688 28412
rect 77622 28362 77638 28396
rect 77672 28394 77688 28396
rect 77672 28364 77710 28394
rect 77910 28364 77936 28394
rect 77672 28362 77688 28364
rect 77622 28346 77688 28362
rect 77622 28086 77688 28102
rect 77622 28052 77638 28086
rect 77672 28084 77688 28086
rect 77672 28054 77710 28084
rect 77910 28054 77936 28084
rect 77672 28052 77688 28054
rect 77622 28036 77688 28052
rect 78439 28396 78505 28412
rect 78439 28394 78455 28396
rect 78182 28364 78208 28394
rect 78408 28364 78455 28394
rect 78439 28362 78455 28364
rect 78489 28362 78505 28396
rect 78439 28346 78505 28362
rect 78439 28086 78505 28102
rect 78439 28084 78455 28086
rect 78182 28054 78208 28084
rect 78408 28054 78455 28084
rect 78439 28052 78455 28054
rect 78489 28052 78505 28086
rect 78439 28036 78505 28052
rect 82342 28396 82408 28412
rect 82342 28362 82358 28396
rect 82392 28394 82408 28396
rect 82392 28364 82430 28394
rect 82630 28364 82656 28394
rect 82392 28362 82408 28364
rect 82342 28346 82408 28362
rect 82342 28086 82408 28102
rect 82342 28052 82358 28086
rect 82392 28084 82408 28086
rect 82392 28054 82430 28084
rect 82630 28054 82656 28084
rect 82392 28052 82408 28054
rect 82342 28036 82408 28052
rect 83159 28396 83225 28412
rect 83159 28394 83175 28396
rect 82902 28364 82928 28394
rect 83128 28364 83175 28394
rect 83159 28362 83175 28364
rect 83209 28362 83225 28396
rect 83159 28346 83225 28362
rect 83159 28086 83225 28102
rect 83159 28084 83175 28086
rect 82902 28054 82928 28084
rect 83128 28054 83175 28084
rect 83159 28052 83175 28054
rect 83209 28052 83225 28086
rect 83159 28036 83225 28052
rect 82342 26686 82408 26702
rect 82342 26652 82358 26686
rect 82392 26684 82408 26686
rect 82392 26654 82430 26684
rect 82630 26654 82656 26684
rect 82392 26652 82408 26654
rect 82342 26636 82408 26652
rect 82342 26376 82408 26392
rect 82342 26342 82358 26376
rect 82392 26374 82408 26376
rect 82392 26344 82430 26374
rect 82630 26344 82656 26374
rect 82392 26342 82408 26344
rect 82342 26326 82408 26342
rect 83159 26686 83225 26702
rect 83159 26684 83175 26686
rect 82902 26654 82928 26684
rect 83128 26654 83175 26684
rect 83159 26652 83175 26654
rect 83209 26652 83225 26686
rect 83159 26636 83225 26652
rect 83159 26376 83225 26392
rect 83159 26374 83175 26376
rect 82902 26344 82928 26374
rect 83128 26344 83175 26374
rect 83159 26342 83175 26344
rect 83209 26342 83225 26376
rect 83159 26326 83225 26342
rect 82342 24976 82408 24992
rect 82342 24942 82358 24976
rect 82392 24974 82408 24976
rect 82392 24944 82430 24974
rect 82630 24944 82656 24974
rect 82392 24942 82408 24944
rect 82342 24926 82408 24942
rect 82342 24666 82408 24682
rect 82342 24632 82358 24666
rect 82392 24664 82408 24666
rect 82392 24634 82430 24664
rect 82630 24634 82656 24664
rect 82392 24632 82408 24634
rect 82342 24616 82408 24632
rect 83159 24976 83225 24992
rect 83159 24974 83175 24976
rect 82902 24944 82928 24974
rect 83128 24944 83175 24974
rect 83159 24942 83175 24944
rect 83209 24942 83225 24976
rect 83159 24926 83225 24942
rect 83159 24666 83225 24682
rect 83159 24664 83175 24666
rect 82902 24634 82928 24664
rect 83128 24634 83175 24664
rect 83159 24632 83175 24634
rect 83209 24632 83225 24666
rect 83159 24616 83225 24632
rect -1948 23266 -1882 23282
rect -1948 23232 -1932 23266
rect -1898 23264 -1882 23266
rect -1898 23234 -1860 23264
rect -1660 23234 -1634 23264
rect -1898 23232 -1882 23234
rect -1948 23216 -1882 23232
rect -1948 22956 -1882 22972
rect -1948 22922 -1932 22956
rect -1898 22954 -1882 22956
rect -1898 22924 -1860 22954
rect -1660 22924 -1634 22954
rect -1898 22922 -1882 22924
rect -1948 22906 -1882 22922
rect -1131 23266 -1065 23282
rect -1131 23264 -1115 23266
rect -1388 23234 -1362 23264
rect -1162 23234 -1115 23264
rect -1131 23232 -1115 23234
rect -1081 23232 -1065 23266
rect -1131 23216 -1065 23232
rect -1131 22956 -1065 22972
rect -1131 22954 -1115 22956
rect -1388 22924 -1362 22954
rect -1162 22924 -1115 22954
rect -1131 22922 -1115 22924
rect -1081 22922 -1065 22956
rect -1131 22906 -1065 22922
rect 82342 23266 82408 23282
rect 82342 23232 82358 23266
rect 82392 23264 82408 23266
rect 82392 23234 82430 23264
rect 82630 23234 82656 23264
rect 82392 23232 82408 23234
rect 82342 23216 82408 23232
rect 82342 22956 82408 22972
rect 82342 22922 82358 22956
rect 82392 22954 82408 22956
rect 82392 22924 82430 22954
rect 82630 22924 82656 22954
rect 82392 22922 82408 22924
rect 82342 22906 82408 22922
rect 83159 23266 83225 23282
rect 83159 23264 83175 23266
rect 82902 23234 82928 23264
rect 83128 23234 83175 23264
rect 83159 23232 83175 23234
rect 83209 23232 83225 23266
rect 83159 23216 83225 23232
rect 83159 22956 83225 22972
rect 83159 22954 83175 22956
rect 82902 22924 82928 22954
rect 83128 22924 83175 22954
rect 83159 22922 83175 22924
rect 83209 22922 83225 22956
rect 83159 22906 83225 22922
rect -1948 21556 -1882 21572
rect -1948 21522 -1932 21556
rect -1898 21554 -1882 21556
rect -1898 21524 -1860 21554
rect -1660 21524 -1634 21554
rect -1898 21522 -1882 21524
rect -1948 21506 -1882 21522
rect -1948 21246 -1882 21262
rect -1948 21212 -1932 21246
rect -1898 21244 -1882 21246
rect -1898 21214 -1860 21244
rect -1660 21214 -1634 21244
rect -1898 21212 -1882 21214
rect -1948 21196 -1882 21212
rect -1131 21556 -1065 21572
rect -1131 21554 -1115 21556
rect -1388 21524 -1362 21554
rect -1162 21524 -1115 21554
rect -1131 21522 -1115 21524
rect -1081 21522 -1065 21556
rect -1131 21506 -1065 21522
rect -1131 21246 -1065 21262
rect -1131 21244 -1115 21246
rect -1388 21214 -1362 21244
rect -1162 21214 -1115 21244
rect -1131 21212 -1115 21214
rect -1081 21212 -1065 21246
rect -1131 21196 -1065 21212
rect 82342 21556 82408 21572
rect 82342 21522 82358 21556
rect 82392 21554 82408 21556
rect 82392 21524 82430 21554
rect 82630 21524 82656 21554
rect 82392 21522 82408 21524
rect 82342 21506 82408 21522
rect 82342 21246 82408 21262
rect 82342 21212 82358 21246
rect 82392 21244 82408 21246
rect 82392 21214 82430 21244
rect 82630 21214 82656 21244
rect 82392 21212 82408 21214
rect 82342 21196 82408 21212
rect 83159 21556 83225 21572
rect 83159 21554 83175 21556
rect 82902 21524 82928 21554
rect 83128 21524 83175 21554
rect 83159 21522 83175 21524
rect 83209 21522 83225 21556
rect 83159 21506 83225 21522
rect 83159 21246 83225 21262
rect 83159 21244 83175 21246
rect 82902 21214 82928 21244
rect 83128 21214 83175 21244
rect 83159 21212 83175 21214
rect 83209 21212 83225 21246
rect 83159 21196 83225 21212
rect -1948 19846 -1882 19862
rect -1948 19812 -1932 19846
rect -1898 19844 -1882 19846
rect -1898 19814 -1860 19844
rect -1660 19814 -1634 19844
rect -1898 19812 -1882 19814
rect -1948 19796 -1882 19812
rect -1948 19536 -1882 19552
rect -1948 19502 -1932 19536
rect -1898 19534 -1882 19536
rect -1898 19504 -1860 19534
rect -1660 19504 -1634 19534
rect -1898 19502 -1882 19504
rect -1948 19486 -1882 19502
rect -1131 19846 -1065 19862
rect -1131 19844 -1115 19846
rect -1388 19814 -1362 19844
rect -1162 19814 -1115 19844
rect -1131 19812 -1115 19814
rect -1081 19812 -1065 19846
rect -1131 19796 -1065 19812
rect -1131 19536 -1065 19552
rect -1131 19534 -1115 19536
rect -1388 19504 -1362 19534
rect -1162 19504 -1115 19534
rect -1131 19502 -1115 19504
rect -1081 19502 -1065 19536
rect -1131 19486 -1065 19502
rect 82342 19846 82408 19862
rect 82342 19812 82358 19846
rect 82392 19844 82408 19846
rect 82392 19814 82430 19844
rect 82630 19814 82656 19844
rect 82392 19812 82408 19814
rect 82342 19796 82408 19812
rect 82342 19536 82408 19552
rect 82342 19502 82358 19536
rect 82392 19534 82408 19536
rect 82392 19504 82430 19534
rect 82630 19504 82656 19534
rect 82392 19502 82408 19504
rect 82342 19486 82408 19502
rect 83159 19846 83225 19862
rect 83159 19844 83175 19846
rect 82902 19814 82928 19844
rect 83128 19814 83175 19844
rect 83159 19812 83175 19814
rect 83209 19812 83225 19846
rect 83159 19796 83225 19812
rect 83159 19536 83225 19552
rect 83159 19534 83175 19536
rect 82902 19504 82928 19534
rect 83128 19504 83175 19534
rect 83159 19502 83175 19504
rect 83209 19502 83225 19536
rect 83159 19486 83225 19502
rect -1948 18136 -1882 18152
rect -1948 18102 -1932 18136
rect -1898 18134 -1882 18136
rect -1898 18104 -1860 18134
rect -1660 18104 -1634 18134
rect -1898 18102 -1882 18104
rect -1948 18086 -1882 18102
rect -1948 17826 -1882 17842
rect -1948 17792 -1932 17826
rect -1898 17824 -1882 17826
rect -1898 17794 -1860 17824
rect -1660 17794 -1634 17824
rect -1898 17792 -1882 17794
rect -1948 17776 -1882 17792
rect -1131 18136 -1065 18152
rect -1131 18134 -1115 18136
rect -1388 18104 -1362 18134
rect -1162 18104 -1115 18134
rect -1131 18102 -1115 18104
rect -1081 18102 -1065 18136
rect -1131 18086 -1065 18102
rect -1131 17826 -1065 17842
rect -1131 17824 -1115 17826
rect -1388 17794 -1362 17824
rect -1162 17794 -1115 17824
rect -1131 17792 -1115 17794
rect -1081 17792 -1065 17826
rect -1131 17776 -1065 17792
rect 82342 18136 82408 18152
rect 82342 18102 82358 18136
rect 82392 18134 82408 18136
rect 82392 18104 82430 18134
rect 82630 18104 82656 18134
rect 82392 18102 82408 18104
rect 82342 18086 82408 18102
rect 82342 17826 82408 17842
rect 82342 17792 82358 17826
rect 82392 17824 82408 17826
rect 82392 17794 82430 17824
rect 82630 17794 82656 17824
rect 82392 17792 82408 17794
rect 82342 17776 82408 17792
rect 83159 18136 83225 18152
rect 83159 18134 83175 18136
rect 82902 18104 82928 18134
rect 83128 18104 83175 18134
rect 83159 18102 83175 18104
rect 83209 18102 83225 18136
rect 83159 18086 83225 18102
rect 83159 17826 83225 17842
rect 83159 17824 83175 17826
rect 82902 17794 82928 17824
rect 83128 17794 83175 17824
rect 83159 17792 83175 17794
rect 83209 17792 83225 17826
rect 83159 17776 83225 17792
rect -1948 16426 -1882 16442
rect -1948 16392 -1932 16426
rect -1898 16424 -1882 16426
rect -1898 16394 -1860 16424
rect -1660 16394 -1634 16424
rect -1898 16392 -1882 16394
rect -1948 16376 -1882 16392
rect -1948 16116 -1882 16132
rect -1948 16082 -1932 16116
rect -1898 16114 -1882 16116
rect -1898 16084 -1860 16114
rect -1660 16084 -1634 16114
rect -1898 16082 -1882 16084
rect -1948 16066 -1882 16082
rect -1131 16426 -1065 16442
rect -1131 16424 -1115 16426
rect -1388 16394 -1362 16424
rect -1162 16394 -1115 16424
rect -1131 16392 -1115 16394
rect -1081 16392 -1065 16426
rect -1131 16376 -1065 16392
rect -1131 16116 -1065 16132
rect -1131 16114 -1115 16116
rect -1388 16084 -1362 16114
rect -1162 16084 -1115 16114
rect -1131 16082 -1115 16084
rect -1081 16082 -1065 16116
rect -1131 16066 -1065 16082
rect 82342 16426 82408 16442
rect 82342 16392 82358 16426
rect 82392 16424 82408 16426
rect 82392 16394 82430 16424
rect 82630 16394 82656 16424
rect 82392 16392 82408 16394
rect 82342 16376 82408 16392
rect 82342 16116 82408 16132
rect 82342 16082 82358 16116
rect 82392 16114 82408 16116
rect 82392 16084 82430 16114
rect 82630 16084 82656 16114
rect 82392 16082 82408 16084
rect 82342 16066 82408 16082
rect 83159 16426 83225 16442
rect 83159 16424 83175 16426
rect 82902 16394 82928 16424
rect 83128 16394 83175 16424
rect 83159 16392 83175 16394
rect 83209 16392 83225 16426
rect 83159 16376 83225 16392
rect 83159 16116 83225 16132
rect 83159 16114 83175 16116
rect 82902 16084 82928 16114
rect 83128 16084 83175 16114
rect 83159 16082 83175 16084
rect 83209 16082 83225 16116
rect 83159 16066 83225 16082
rect -1948 14716 -1882 14732
rect -1948 14682 -1932 14716
rect -1898 14714 -1882 14716
rect -1898 14684 -1860 14714
rect -1660 14684 -1634 14714
rect -1898 14682 -1882 14684
rect -1948 14666 -1882 14682
rect -1948 14406 -1882 14422
rect -1948 14372 -1932 14406
rect -1898 14404 -1882 14406
rect -1898 14374 -1860 14404
rect -1660 14374 -1634 14404
rect -1898 14372 -1882 14374
rect -1948 14356 -1882 14372
rect -1131 14716 -1065 14732
rect -1131 14714 -1115 14716
rect -1388 14684 -1362 14714
rect -1162 14684 -1115 14714
rect -1131 14682 -1115 14684
rect -1081 14682 -1065 14716
rect -1131 14666 -1065 14682
rect -1131 14406 -1065 14422
rect -1131 14404 -1115 14406
rect -1388 14374 -1362 14404
rect -1162 14374 -1115 14404
rect -1131 14372 -1115 14374
rect -1081 14372 -1065 14406
rect -1131 14356 -1065 14372
rect 82342 14716 82408 14732
rect 82342 14682 82358 14716
rect 82392 14714 82408 14716
rect 82392 14684 82430 14714
rect 82630 14684 82656 14714
rect 82392 14682 82408 14684
rect 82342 14666 82408 14682
rect 82342 14406 82408 14422
rect 82342 14372 82358 14406
rect 82392 14404 82408 14406
rect 82392 14374 82430 14404
rect 82630 14374 82656 14404
rect 82392 14372 82408 14374
rect 82342 14356 82408 14372
rect 83159 14716 83225 14732
rect 83159 14714 83175 14716
rect 82902 14684 82928 14714
rect 83128 14684 83175 14714
rect 83159 14682 83175 14684
rect 83209 14682 83225 14716
rect 83159 14666 83225 14682
rect 83159 14406 83225 14422
rect 83159 14404 83175 14406
rect 82902 14374 82928 14404
rect 83128 14374 83175 14404
rect 83159 14372 83175 14374
rect 83209 14372 83225 14406
rect 83159 14356 83225 14372
rect -1948 13006 -1882 13022
rect -1948 12972 -1932 13006
rect -1898 13004 -1882 13006
rect -1898 12974 -1860 13004
rect -1660 12974 -1634 13004
rect -1898 12972 -1882 12974
rect -1948 12956 -1882 12972
rect -1948 12696 -1882 12712
rect -1948 12662 -1932 12696
rect -1898 12694 -1882 12696
rect -1898 12664 -1860 12694
rect -1660 12664 -1634 12694
rect -1898 12662 -1882 12664
rect -1948 12646 -1882 12662
rect -1131 13006 -1065 13022
rect -1131 13004 -1115 13006
rect -1388 12974 -1362 13004
rect -1162 12974 -1115 13004
rect -1131 12972 -1115 12974
rect -1081 12972 -1065 13006
rect -1131 12956 -1065 12972
rect -1131 12696 -1065 12712
rect -1131 12694 -1115 12696
rect -1388 12664 -1362 12694
rect -1162 12664 -1115 12694
rect -1131 12662 -1115 12664
rect -1081 12662 -1065 12696
rect -1131 12646 -1065 12662
rect 82342 13006 82408 13022
rect 82342 12972 82358 13006
rect 82392 13004 82408 13006
rect 82392 12974 82430 13004
rect 82630 12974 82656 13004
rect 82392 12972 82408 12974
rect 82342 12956 82408 12972
rect 82342 12696 82408 12712
rect 82342 12662 82358 12696
rect 82392 12694 82408 12696
rect 82392 12664 82430 12694
rect 82630 12664 82656 12694
rect 82392 12662 82408 12664
rect 82342 12646 82408 12662
rect 83159 13006 83225 13022
rect 83159 13004 83175 13006
rect 82902 12974 82928 13004
rect 83128 12974 83175 13004
rect 83159 12972 83175 12974
rect 83209 12972 83225 13006
rect 83159 12956 83225 12972
rect 83159 12696 83225 12712
rect 83159 12694 83175 12696
rect 82902 12664 82928 12694
rect 83128 12664 83175 12694
rect 83159 12662 83175 12664
rect 83209 12662 83225 12696
rect 83159 12646 83225 12662
rect -1948 11296 -1882 11312
rect -1948 11262 -1932 11296
rect -1898 11294 -1882 11296
rect -1898 11264 -1860 11294
rect -1660 11264 -1634 11294
rect -1898 11262 -1882 11264
rect -1948 11246 -1882 11262
rect -1948 10986 -1882 11002
rect -1948 10952 -1932 10986
rect -1898 10984 -1882 10986
rect -1898 10954 -1860 10984
rect -1660 10954 -1634 10984
rect -1898 10952 -1882 10954
rect -1948 10936 -1882 10952
rect -1131 11296 -1065 11312
rect -1131 11294 -1115 11296
rect -1388 11264 -1362 11294
rect -1162 11264 -1115 11294
rect -1131 11262 -1115 11264
rect -1081 11262 -1065 11296
rect -1131 11246 -1065 11262
rect -1131 10986 -1065 11002
rect -1131 10984 -1115 10986
rect -1388 10954 -1362 10984
rect -1162 10954 -1115 10984
rect -1131 10952 -1115 10954
rect -1081 10952 -1065 10986
rect -1131 10936 -1065 10952
rect 82342 11296 82408 11312
rect 82342 11262 82358 11296
rect 82392 11294 82408 11296
rect 82392 11264 82430 11294
rect 82630 11264 82656 11294
rect 82392 11262 82408 11264
rect 82342 11246 82408 11262
rect 82342 10986 82408 11002
rect 82342 10952 82358 10986
rect 82392 10984 82408 10986
rect 82392 10954 82430 10984
rect 82630 10954 82656 10984
rect 82392 10952 82408 10954
rect 82342 10936 82408 10952
rect 83159 11296 83225 11312
rect 83159 11294 83175 11296
rect 82902 11264 82928 11294
rect 83128 11264 83175 11294
rect 83159 11262 83175 11264
rect 83209 11262 83225 11296
rect 83159 11246 83225 11262
rect 83159 10986 83225 11002
rect 83159 10984 83175 10986
rect 82902 10954 82928 10984
rect 83128 10954 83175 10984
rect 83159 10952 83175 10954
rect 83209 10952 83225 10986
rect 83159 10936 83225 10952
rect -1948 9586 -1882 9602
rect -1948 9552 -1932 9586
rect -1898 9584 -1882 9586
rect -1898 9554 -1860 9584
rect -1660 9554 -1634 9584
rect -1898 9552 -1882 9554
rect -1948 9536 -1882 9552
rect -1948 9276 -1882 9292
rect -1948 9242 -1932 9276
rect -1898 9274 -1882 9276
rect -1898 9244 -1860 9274
rect -1660 9244 -1634 9274
rect -1898 9242 -1882 9244
rect -1948 9226 -1882 9242
rect -1131 9586 -1065 9602
rect -1131 9584 -1115 9586
rect -1388 9554 -1362 9584
rect -1162 9554 -1115 9584
rect -1131 9552 -1115 9554
rect -1081 9552 -1065 9586
rect -1131 9536 -1065 9552
rect -1131 9276 -1065 9292
rect -1131 9274 -1115 9276
rect -1388 9244 -1362 9274
rect -1162 9244 -1115 9274
rect -1131 9242 -1115 9244
rect -1081 9242 -1065 9276
rect -1131 9226 -1065 9242
rect 82342 9586 82408 9602
rect 82342 9552 82358 9586
rect 82392 9584 82408 9586
rect 82392 9554 82430 9584
rect 82630 9554 82656 9584
rect 82392 9552 82408 9554
rect 82342 9536 82408 9552
rect 82342 9276 82408 9292
rect 82342 9242 82358 9276
rect 82392 9274 82408 9276
rect 82392 9244 82430 9274
rect 82630 9244 82656 9274
rect 82392 9242 82408 9244
rect 82342 9226 82408 9242
rect 83159 9586 83225 9602
rect 83159 9584 83175 9586
rect 82902 9554 82928 9584
rect 83128 9554 83175 9584
rect 83159 9552 83175 9554
rect 83209 9552 83225 9586
rect 83159 9536 83225 9552
rect 83159 9276 83225 9292
rect 83159 9274 83175 9276
rect 82902 9244 82928 9274
rect 83128 9244 83175 9274
rect 83159 9242 83175 9244
rect 83209 9242 83225 9276
rect 83159 9226 83225 9242
rect -1948 7876 -1882 7892
rect -1948 7842 -1932 7876
rect -1898 7874 -1882 7876
rect -1898 7844 -1860 7874
rect -1660 7844 -1634 7874
rect -1898 7842 -1882 7844
rect -1948 7826 -1882 7842
rect -1948 7566 -1882 7582
rect -1948 7532 -1932 7566
rect -1898 7564 -1882 7566
rect -1898 7534 -1860 7564
rect -1660 7534 -1634 7564
rect -1898 7532 -1882 7534
rect -1948 7516 -1882 7532
rect -1131 7876 -1065 7892
rect -1131 7874 -1115 7876
rect -1388 7844 -1362 7874
rect -1162 7844 -1115 7874
rect -1131 7842 -1115 7844
rect -1081 7842 -1065 7876
rect -1131 7826 -1065 7842
rect -1131 7566 -1065 7582
rect -1131 7564 -1115 7566
rect -1388 7534 -1362 7564
rect -1162 7534 -1115 7564
rect -1131 7532 -1115 7534
rect -1081 7532 -1065 7566
rect -1131 7516 -1065 7532
rect 82342 7876 82408 7892
rect 82342 7842 82358 7876
rect 82392 7874 82408 7876
rect 82392 7844 82430 7874
rect 82630 7844 82656 7874
rect 82392 7842 82408 7844
rect 82342 7826 82408 7842
rect 82342 7566 82408 7582
rect 82342 7532 82358 7566
rect 82392 7564 82408 7566
rect 82392 7534 82430 7564
rect 82630 7534 82656 7564
rect 82392 7532 82408 7534
rect 82342 7516 82408 7532
rect 83159 7876 83225 7892
rect 83159 7874 83175 7876
rect 82902 7844 82928 7874
rect 83128 7844 83175 7874
rect 83159 7842 83175 7844
rect 83209 7842 83225 7876
rect 83159 7826 83225 7842
rect 83159 7566 83225 7582
rect 83159 7564 83175 7566
rect 82902 7534 82928 7564
rect 83128 7534 83175 7564
rect 83159 7532 83175 7534
rect 83209 7532 83225 7566
rect 83159 7516 83225 7532
rect -1948 6166 -1882 6182
rect -1948 6132 -1932 6166
rect -1898 6164 -1882 6166
rect -1898 6134 -1860 6164
rect -1660 6134 -1634 6164
rect -1898 6132 -1882 6134
rect -1948 6116 -1882 6132
rect -1948 5856 -1882 5872
rect -1948 5822 -1932 5856
rect -1898 5854 -1882 5856
rect -1898 5824 -1860 5854
rect -1660 5824 -1634 5854
rect -1898 5822 -1882 5824
rect -1948 5806 -1882 5822
rect -1131 6166 -1065 6182
rect -1131 6164 -1115 6166
rect -1388 6134 -1362 6164
rect -1162 6134 -1115 6164
rect -1131 6132 -1115 6134
rect -1081 6132 -1065 6166
rect -1131 6116 -1065 6132
rect -1131 5856 -1065 5872
rect -1131 5854 -1115 5856
rect -1388 5824 -1362 5854
rect -1162 5824 -1115 5854
rect -1131 5822 -1115 5824
rect -1081 5822 -1065 5856
rect -1131 5806 -1065 5822
rect 82342 6166 82408 6182
rect 82342 6132 82358 6166
rect 82392 6164 82408 6166
rect 82392 6134 82430 6164
rect 82630 6134 82656 6164
rect 82392 6132 82408 6134
rect 82342 6116 82408 6132
rect 82342 5856 82408 5872
rect 82342 5822 82358 5856
rect 82392 5854 82408 5856
rect 82392 5824 82430 5854
rect 82630 5824 82656 5854
rect 82392 5822 82408 5824
rect 82342 5806 82408 5822
rect 83159 6166 83225 6182
rect 83159 6164 83175 6166
rect 82902 6134 82928 6164
rect 83128 6134 83175 6164
rect 83159 6132 83175 6134
rect 83209 6132 83225 6166
rect 83159 6116 83225 6132
rect 83159 5856 83225 5872
rect 83159 5854 83175 5856
rect 82902 5824 82928 5854
rect 83128 5824 83175 5854
rect 83159 5822 83175 5824
rect 83209 5822 83225 5856
rect 83159 5806 83225 5822
rect -1948 4456 -1882 4472
rect -1948 4422 -1932 4456
rect -1898 4454 -1882 4456
rect -1898 4424 -1860 4454
rect -1660 4424 -1634 4454
rect -1898 4422 -1882 4424
rect -1948 4406 -1882 4422
rect -1948 4146 -1882 4162
rect -1948 4112 -1932 4146
rect -1898 4144 -1882 4146
rect -1898 4114 -1860 4144
rect -1660 4114 -1634 4144
rect -1898 4112 -1882 4114
rect -1948 4096 -1882 4112
rect -1131 4456 -1065 4472
rect -1131 4454 -1115 4456
rect -1388 4424 -1362 4454
rect -1162 4424 -1115 4454
rect -1131 4422 -1115 4424
rect -1081 4422 -1065 4456
rect -1131 4406 -1065 4422
rect -1131 4146 -1065 4162
rect -1131 4144 -1115 4146
rect -1388 4114 -1362 4144
rect -1162 4114 -1115 4144
rect -1131 4112 -1115 4114
rect -1081 4112 -1065 4146
rect -1131 4096 -1065 4112
rect 82342 4456 82408 4472
rect 82342 4422 82358 4456
rect 82392 4454 82408 4456
rect 82392 4424 82430 4454
rect 82630 4424 82656 4454
rect 82392 4422 82408 4424
rect 82342 4406 82408 4422
rect 82342 4146 82408 4162
rect 82342 4112 82358 4146
rect 82392 4144 82408 4146
rect 82392 4114 82430 4144
rect 82630 4114 82656 4144
rect 82392 4112 82408 4114
rect 82342 4096 82408 4112
rect 83159 4456 83225 4472
rect 83159 4454 83175 4456
rect 82902 4424 82928 4454
rect 83128 4424 83175 4454
rect 83159 4422 83175 4424
rect 83209 4422 83225 4456
rect 83159 4406 83225 4422
rect 83159 4146 83225 4162
rect 83159 4144 83175 4146
rect 82902 4114 82928 4144
rect 83128 4114 83175 4144
rect 83159 4112 83175 4114
rect 83209 4112 83225 4146
rect 83159 4096 83225 4112
rect -1948 2746 -1882 2762
rect -1948 2712 -1932 2746
rect -1898 2744 -1882 2746
rect -1898 2714 -1860 2744
rect -1660 2714 -1634 2744
rect -1898 2712 -1882 2714
rect -1948 2696 -1882 2712
rect -1948 2436 -1882 2452
rect -1948 2402 -1932 2436
rect -1898 2434 -1882 2436
rect -1898 2404 -1860 2434
rect -1660 2404 -1634 2434
rect -1898 2402 -1882 2404
rect -1948 2386 -1882 2402
rect -1131 2746 -1065 2762
rect -1131 2744 -1115 2746
rect -1388 2714 -1362 2744
rect -1162 2714 -1115 2744
rect -1131 2712 -1115 2714
rect -1081 2712 -1065 2746
rect -1131 2696 -1065 2712
rect -1131 2436 -1065 2452
rect -1131 2434 -1115 2436
rect -1388 2404 -1362 2434
rect -1162 2404 -1115 2434
rect -1131 2402 -1115 2404
rect -1081 2402 -1065 2436
rect -1131 2386 -1065 2402
rect 82342 2746 82408 2762
rect 82342 2712 82358 2746
rect 82392 2744 82408 2746
rect 82392 2714 82430 2744
rect 82630 2714 82656 2744
rect 82392 2712 82408 2714
rect 82342 2696 82408 2712
rect 82342 2436 82408 2452
rect 82342 2402 82358 2436
rect 82392 2434 82408 2436
rect 82392 2404 82430 2434
rect 82630 2404 82656 2434
rect 82392 2402 82408 2404
rect 82342 2386 82408 2402
rect 83159 2746 83225 2762
rect 83159 2744 83175 2746
rect 82902 2714 82928 2744
rect 83128 2714 83175 2744
rect 83159 2712 83175 2714
rect 83209 2712 83225 2746
rect 83159 2696 83225 2712
rect 83159 2436 83225 2452
rect 83159 2434 83175 2436
rect 82902 2404 82928 2434
rect 83128 2404 83175 2434
rect 83159 2402 83175 2404
rect 83209 2402 83225 2436
rect 83159 2386 83225 2402
rect -1948 1036 -1882 1052
rect -1948 1002 -1932 1036
rect -1898 1034 -1882 1036
rect -1898 1004 -1860 1034
rect -1660 1004 -1634 1034
rect -1898 1002 -1882 1004
rect -1948 986 -1882 1002
rect -1948 726 -1882 742
rect -1948 692 -1932 726
rect -1898 724 -1882 726
rect -1898 694 -1860 724
rect -1660 694 -1634 724
rect -1898 692 -1882 694
rect -1948 676 -1882 692
rect -1131 1036 -1065 1052
rect -1131 1034 -1115 1036
rect -1388 1004 -1362 1034
rect -1162 1004 -1115 1034
rect -1131 1002 -1115 1004
rect -1081 1002 -1065 1036
rect -1131 986 -1065 1002
rect -1131 726 -1065 742
rect -1131 724 -1115 726
rect -1388 694 -1362 724
rect -1162 694 -1115 724
rect -1131 692 -1115 694
rect -1081 692 -1065 726
rect -1131 676 -1065 692
rect 82342 1036 82408 1052
rect 82342 1002 82358 1036
rect 82392 1034 82408 1036
rect 82392 1004 82430 1034
rect 82630 1004 82656 1034
rect 82392 1002 82408 1004
rect 82342 986 82408 1002
rect 82342 726 82408 742
rect 82342 692 82358 726
rect 82392 724 82408 726
rect 82392 694 82430 724
rect 82630 694 82656 724
rect 82392 692 82408 694
rect 82342 676 82408 692
rect 83159 1036 83225 1052
rect 83159 1034 83175 1036
rect 82902 1004 82928 1034
rect 83128 1004 83175 1034
rect 83159 1002 83175 1004
rect 83209 1002 83225 1036
rect 83159 986 83225 1002
rect 83159 726 83225 742
rect 83159 724 83175 726
rect 82902 694 82928 724
rect 83128 694 83175 724
rect 83159 692 83175 694
rect 83209 692 83225 726
rect 83159 676 83225 692
rect -1948 -674 -1882 -658
rect -1948 -708 -1932 -674
rect -1898 -676 -1882 -674
rect -1898 -706 -1860 -676
rect -1660 -706 -1634 -676
rect -1898 -708 -1882 -706
rect -1948 -724 -1882 -708
rect -1948 -984 -1882 -968
rect -1948 -1018 -1932 -984
rect -1898 -986 -1882 -984
rect -1898 -1016 -1860 -986
rect -1660 -1016 -1634 -986
rect -1898 -1018 -1882 -1016
rect -1948 -1034 -1882 -1018
rect -1131 -674 -1065 -658
rect -1131 -676 -1115 -674
rect -1388 -706 -1362 -676
rect -1162 -706 -1115 -676
rect -1131 -708 -1115 -706
rect -1081 -708 -1065 -674
rect -1131 -724 -1065 -708
rect -1131 -984 -1065 -968
rect -1131 -986 -1115 -984
rect -1388 -1016 -1362 -986
rect -1162 -1016 -1115 -986
rect -1131 -1018 -1115 -1016
rect -1081 -1018 -1065 -984
rect -1131 -1034 -1065 -1018
rect 2772 -674 2838 -658
rect 2772 -708 2788 -674
rect 2822 -676 2838 -674
rect 2822 -706 2860 -676
rect 3060 -706 3086 -676
rect 2822 -708 2838 -706
rect 2772 -724 2838 -708
rect 2772 -984 2838 -968
rect 2772 -1018 2788 -984
rect 2822 -986 2838 -984
rect 2822 -1016 2860 -986
rect 3060 -1016 3086 -986
rect 2822 -1018 2838 -1016
rect 2772 -1034 2838 -1018
rect 3589 -674 3655 -658
rect 3589 -676 3605 -674
rect 3332 -706 3358 -676
rect 3558 -706 3605 -676
rect 3589 -708 3605 -706
rect 3639 -708 3655 -674
rect 3589 -724 3655 -708
rect 3589 -984 3655 -968
rect 3589 -986 3605 -984
rect 3332 -1016 3358 -986
rect 3558 -1016 3605 -986
rect 3589 -1018 3605 -1016
rect 3639 -1018 3655 -984
rect 3589 -1034 3655 -1018
rect 7762 -674 7828 -658
rect 7762 -708 7778 -674
rect 7812 -676 7828 -674
rect 7812 -706 7850 -676
rect 8050 -706 8076 -676
rect 7812 -708 7828 -706
rect 7762 -724 7828 -708
rect 7762 -984 7828 -968
rect 7762 -1018 7778 -984
rect 7812 -986 7828 -984
rect 7812 -1016 7850 -986
rect 8050 -1016 8076 -986
rect 7812 -1018 7828 -1016
rect 7762 -1034 7828 -1018
rect 8579 -674 8645 -658
rect 8579 -676 8595 -674
rect 8322 -706 8348 -676
rect 8548 -706 8595 -676
rect 8579 -708 8595 -706
rect 8629 -708 8645 -674
rect 8579 -724 8645 -708
rect 8579 -984 8645 -968
rect 8579 -986 8595 -984
rect 8322 -1016 8348 -986
rect 8548 -1016 8595 -986
rect 8579 -1018 8595 -1016
rect 8629 -1018 8645 -984
rect 8579 -1034 8645 -1018
rect 12752 -674 12818 -658
rect 12752 -708 12768 -674
rect 12802 -676 12818 -674
rect 12802 -706 12840 -676
rect 13040 -706 13066 -676
rect 12802 -708 12818 -706
rect 12752 -724 12818 -708
rect 12752 -984 12818 -968
rect 12752 -1018 12768 -984
rect 12802 -986 12818 -984
rect 12802 -1016 12840 -986
rect 13040 -1016 13066 -986
rect 12802 -1018 12818 -1016
rect 12752 -1034 12818 -1018
rect 13569 -674 13635 -658
rect 13569 -676 13585 -674
rect 13312 -706 13338 -676
rect 13538 -706 13585 -676
rect 13569 -708 13585 -706
rect 13619 -708 13635 -674
rect 13569 -724 13635 -708
rect 13569 -984 13635 -968
rect 13569 -986 13585 -984
rect 13312 -1016 13338 -986
rect 13538 -1016 13585 -986
rect 13569 -1018 13585 -1016
rect 13619 -1018 13635 -984
rect 13569 -1034 13635 -1018
rect 17742 -674 17808 -658
rect 17742 -708 17758 -674
rect 17792 -676 17808 -674
rect 17792 -706 17830 -676
rect 18030 -706 18056 -676
rect 17792 -708 17808 -706
rect 17742 -724 17808 -708
rect 17742 -984 17808 -968
rect 17742 -1018 17758 -984
rect 17792 -986 17808 -984
rect 17792 -1016 17830 -986
rect 18030 -1016 18056 -986
rect 17792 -1018 17808 -1016
rect 17742 -1034 17808 -1018
rect 18559 -674 18625 -658
rect 18559 -676 18575 -674
rect 18302 -706 18328 -676
rect 18528 -706 18575 -676
rect 18559 -708 18575 -706
rect 18609 -708 18625 -674
rect 18559 -724 18625 -708
rect 18559 -984 18625 -968
rect 18559 -986 18575 -984
rect 18302 -1016 18328 -986
rect 18528 -1016 18575 -986
rect 18559 -1018 18575 -1016
rect 18609 -1018 18625 -984
rect 18559 -1034 18625 -1018
rect 22732 -674 22798 -658
rect 22732 -708 22748 -674
rect 22782 -676 22798 -674
rect 22782 -706 22820 -676
rect 23020 -706 23046 -676
rect 22782 -708 22798 -706
rect 22732 -724 22798 -708
rect 22732 -984 22798 -968
rect 22732 -1018 22748 -984
rect 22782 -986 22798 -984
rect 22782 -1016 22820 -986
rect 23020 -1016 23046 -986
rect 22782 -1018 22798 -1016
rect 22732 -1034 22798 -1018
rect 23549 -674 23615 -658
rect 23549 -676 23565 -674
rect 23292 -706 23318 -676
rect 23518 -706 23565 -676
rect 23549 -708 23565 -706
rect 23599 -708 23615 -674
rect 23549 -724 23615 -708
rect 23549 -984 23615 -968
rect 23549 -986 23565 -984
rect 23292 -1016 23318 -986
rect 23518 -1016 23565 -986
rect 23549 -1018 23565 -1016
rect 23599 -1018 23615 -984
rect 23549 -1034 23615 -1018
rect 27722 -674 27788 -658
rect 27722 -708 27738 -674
rect 27772 -676 27788 -674
rect 27772 -706 27810 -676
rect 28010 -706 28036 -676
rect 27772 -708 27788 -706
rect 27722 -724 27788 -708
rect 27722 -984 27788 -968
rect 27722 -1018 27738 -984
rect 27772 -986 27788 -984
rect 27772 -1016 27810 -986
rect 28010 -1016 28036 -986
rect 27772 -1018 27788 -1016
rect 27722 -1034 27788 -1018
rect 28539 -674 28605 -658
rect 28539 -676 28555 -674
rect 28282 -706 28308 -676
rect 28508 -706 28555 -676
rect 28539 -708 28555 -706
rect 28589 -708 28605 -674
rect 28539 -724 28605 -708
rect 28539 -984 28605 -968
rect 28539 -986 28555 -984
rect 28282 -1016 28308 -986
rect 28508 -1016 28555 -986
rect 28539 -1018 28555 -1016
rect 28589 -1018 28605 -984
rect 28539 -1034 28605 -1018
rect 32712 -674 32778 -658
rect 32712 -708 32728 -674
rect 32762 -676 32778 -674
rect 32762 -706 32800 -676
rect 33000 -706 33026 -676
rect 32762 -708 32778 -706
rect 32712 -724 32778 -708
rect 32712 -984 32778 -968
rect 32712 -1018 32728 -984
rect 32762 -986 32778 -984
rect 32762 -1016 32800 -986
rect 33000 -1016 33026 -986
rect 32762 -1018 32778 -1016
rect 32712 -1034 32778 -1018
rect 33529 -674 33595 -658
rect 33529 -676 33545 -674
rect 33272 -706 33298 -676
rect 33498 -706 33545 -676
rect 33529 -708 33545 -706
rect 33579 -708 33595 -674
rect 33529 -724 33595 -708
rect 33529 -984 33595 -968
rect 33529 -986 33545 -984
rect 33272 -1016 33298 -986
rect 33498 -1016 33545 -986
rect 33529 -1018 33545 -1016
rect 33579 -1018 33595 -984
rect 33529 -1034 33595 -1018
rect 37702 -674 37768 -658
rect 37702 -708 37718 -674
rect 37752 -676 37768 -674
rect 37752 -706 37790 -676
rect 37990 -706 38016 -676
rect 37752 -708 37768 -706
rect 37702 -724 37768 -708
rect 37702 -984 37768 -968
rect 37702 -1018 37718 -984
rect 37752 -986 37768 -984
rect 37752 -1016 37790 -986
rect 37990 -1016 38016 -986
rect 37752 -1018 37768 -1016
rect 37702 -1034 37768 -1018
rect 38519 -674 38585 -658
rect 38519 -676 38535 -674
rect 38262 -706 38288 -676
rect 38488 -706 38535 -676
rect 38519 -708 38535 -706
rect 38569 -708 38585 -674
rect 38519 -724 38585 -708
rect 38519 -984 38585 -968
rect 38519 -986 38535 -984
rect 38262 -1016 38288 -986
rect 38488 -1016 38535 -986
rect 38519 -1018 38535 -1016
rect 38569 -1018 38585 -984
rect 38519 -1034 38585 -1018
rect 42692 -674 42758 -658
rect 42692 -708 42708 -674
rect 42742 -676 42758 -674
rect 42742 -706 42780 -676
rect 42980 -706 43006 -676
rect 42742 -708 42758 -706
rect 42692 -724 42758 -708
rect 42692 -984 42758 -968
rect 42692 -1018 42708 -984
rect 42742 -986 42758 -984
rect 42742 -1016 42780 -986
rect 42980 -1016 43006 -986
rect 42742 -1018 42758 -1016
rect 42692 -1034 42758 -1018
rect 43509 -674 43575 -658
rect 43509 -676 43525 -674
rect 43252 -706 43278 -676
rect 43478 -706 43525 -676
rect 43509 -708 43525 -706
rect 43559 -708 43575 -674
rect 43509 -724 43575 -708
rect 43509 -984 43575 -968
rect 43509 -986 43525 -984
rect 43252 -1016 43278 -986
rect 43478 -1016 43525 -986
rect 43509 -1018 43525 -1016
rect 43559 -1018 43575 -984
rect 43509 -1034 43575 -1018
rect 47682 -674 47748 -658
rect 47682 -708 47698 -674
rect 47732 -676 47748 -674
rect 47732 -706 47770 -676
rect 47970 -706 47996 -676
rect 47732 -708 47748 -706
rect 47682 -724 47748 -708
rect 47682 -984 47748 -968
rect 47682 -1018 47698 -984
rect 47732 -986 47748 -984
rect 47732 -1016 47770 -986
rect 47970 -1016 47996 -986
rect 47732 -1018 47748 -1016
rect 47682 -1034 47748 -1018
rect 48499 -674 48565 -658
rect 48499 -676 48515 -674
rect 48242 -706 48268 -676
rect 48468 -706 48515 -676
rect 48499 -708 48515 -706
rect 48549 -708 48565 -674
rect 48499 -724 48565 -708
rect 48499 -984 48565 -968
rect 48499 -986 48515 -984
rect 48242 -1016 48268 -986
rect 48468 -1016 48515 -986
rect 48499 -1018 48515 -1016
rect 48549 -1018 48565 -984
rect 48499 -1034 48565 -1018
rect 52672 -674 52738 -658
rect 52672 -708 52688 -674
rect 52722 -676 52738 -674
rect 52722 -706 52760 -676
rect 52960 -706 52986 -676
rect 52722 -708 52738 -706
rect 52672 -724 52738 -708
rect 52672 -984 52738 -968
rect 52672 -1018 52688 -984
rect 52722 -986 52738 -984
rect 52722 -1016 52760 -986
rect 52960 -1016 52986 -986
rect 52722 -1018 52738 -1016
rect 52672 -1034 52738 -1018
rect 53489 -674 53555 -658
rect 53489 -676 53505 -674
rect 53232 -706 53258 -676
rect 53458 -706 53505 -676
rect 53489 -708 53505 -706
rect 53539 -708 53555 -674
rect 53489 -724 53555 -708
rect 53489 -984 53555 -968
rect 53489 -986 53505 -984
rect 53232 -1016 53258 -986
rect 53458 -1016 53505 -986
rect 53489 -1018 53505 -1016
rect 53539 -1018 53555 -984
rect 53489 -1034 53555 -1018
rect 57662 -674 57728 -658
rect 57662 -708 57678 -674
rect 57712 -676 57728 -674
rect 57712 -706 57750 -676
rect 57950 -706 57976 -676
rect 57712 -708 57728 -706
rect 57662 -724 57728 -708
rect 57662 -984 57728 -968
rect 57662 -1018 57678 -984
rect 57712 -986 57728 -984
rect 57712 -1016 57750 -986
rect 57950 -1016 57976 -986
rect 57712 -1018 57728 -1016
rect 57662 -1034 57728 -1018
rect 58479 -674 58545 -658
rect 58479 -676 58495 -674
rect 58222 -706 58248 -676
rect 58448 -706 58495 -676
rect 58479 -708 58495 -706
rect 58529 -708 58545 -674
rect 58479 -724 58545 -708
rect 58479 -984 58545 -968
rect 58479 -986 58495 -984
rect 58222 -1016 58248 -986
rect 58448 -1016 58495 -986
rect 58479 -1018 58495 -1016
rect 58529 -1018 58545 -984
rect 58479 -1034 58545 -1018
rect 62652 -674 62718 -658
rect 62652 -708 62668 -674
rect 62702 -676 62718 -674
rect 62702 -706 62740 -676
rect 62940 -706 62966 -676
rect 62702 -708 62718 -706
rect 62652 -724 62718 -708
rect 62652 -984 62718 -968
rect 62652 -1018 62668 -984
rect 62702 -986 62718 -984
rect 62702 -1016 62740 -986
rect 62940 -1016 62966 -986
rect 62702 -1018 62718 -1016
rect 62652 -1034 62718 -1018
rect 63469 -674 63535 -658
rect 63469 -676 63485 -674
rect 63212 -706 63238 -676
rect 63438 -706 63485 -676
rect 63469 -708 63485 -706
rect 63519 -708 63535 -674
rect 63469 -724 63535 -708
rect 63469 -984 63535 -968
rect 63469 -986 63485 -984
rect 63212 -1016 63238 -986
rect 63438 -1016 63485 -986
rect 63469 -1018 63485 -1016
rect 63519 -1018 63535 -984
rect 63469 -1034 63535 -1018
rect 67642 -674 67708 -658
rect 67642 -708 67658 -674
rect 67692 -676 67708 -674
rect 67692 -706 67730 -676
rect 67930 -706 67956 -676
rect 67692 -708 67708 -706
rect 67642 -724 67708 -708
rect 67642 -984 67708 -968
rect 67642 -1018 67658 -984
rect 67692 -986 67708 -984
rect 67692 -1016 67730 -986
rect 67930 -1016 67956 -986
rect 67692 -1018 67708 -1016
rect 67642 -1034 67708 -1018
rect 68459 -674 68525 -658
rect 68459 -676 68475 -674
rect 68202 -706 68228 -676
rect 68428 -706 68475 -676
rect 68459 -708 68475 -706
rect 68509 -708 68525 -674
rect 68459 -724 68525 -708
rect 68459 -984 68525 -968
rect 68459 -986 68475 -984
rect 68202 -1016 68228 -986
rect 68428 -1016 68475 -986
rect 68459 -1018 68475 -1016
rect 68509 -1018 68525 -984
rect 68459 -1034 68525 -1018
rect 72632 -674 72698 -658
rect 72632 -708 72648 -674
rect 72682 -676 72698 -674
rect 72682 -706 72720 -676
rect 72920 -706 72946 -676
rect 72682 -708 72698 -706
rect 72632 -724 72698 -708
rect 72632 -984 72698 -968
rect 72632 -1018 72648 -984
rect 72682 -986 72698 -984
rect 72682 -1016 72720 -986
rect 72920 -1016 72946 -986
rect 72682 -1018 72698 -1016
rect 72632 -1034 72698 -1018
rect 73449 -674 73515 -658
rect 73449 -676 73465 -674
rect 73192 -706 73218 -676
rect 73418 -706 73465 -676
rect 73449 -708 73465 -706
rect 73499 -708 73515 -674
rect 73449 -724 73515 -708
rect 73449 -984 73515 -968
rect 73449 -986 73465 -984
rect 73192 -1016 73218 -986
rect 73418 -1016 73465 -986
rect 73449 -1018 73465 -1016
rect 73499 -1018 73515 -984
rect 73449 -1034 73515 -1018
rect 77622 -674 77688 -658
rect 77622 -708 77638 -674
rect 77672 -676 77688 -674
rect 77672 -706 77710 -676
rect 77910 -706 77936 -676
rect 77672 -708 77688 -706
rect 77622 -724 77688 -708
rect 77622 -984 77688 -968
rect 77622 -1018 77638 -984
rect 77672 -986 77688 -984
rect 77672 -1016 77710 -986
rect 77910 -1016 77936 -986
rect 77672 -1018 77688 -1016
rect 77622 -1034 77688 -1018
rect 78439 -674 78505 -658
rect 78439 -676 78455 -674
rect 78182 -706 78208 -676
rect 78408 -706 78455 -676
rect 78439 -708 78455 -706
rect 78489 -708 78505 -674
rect 78439 -724 78505 -708
rect 78439 -984 78505 -968
rect 78439 -986 78455 -984
rect 78182 -1016 78208 -986
rect 78408 -1016 78455 -986
rect 78439 -1018 78455 -1016
rect 78489 -1018 78505 -984
rect 78439 -1034 78505 -1018
rect 82342 -674 82408 -658
rect 82342 -708 82358 -674
rect 82392 -676 82408 -674
rect 82392 -706 82430 -676
rect 82630 -706 82656 -676
rect 82392 -708 82408 -706
rect 82342 -724 82408 -708
rect 82342 -984 82408 -968
rect 82342 -1018 82358 -984
rect 82392 -986 82408 -984
rect 82392 -1016 82430 -986
rect 82630 -1016 82656 -986
rect 82392 -1018 82408 -1016
rect 82342 -1034 82408 -1018
rect 83159 -674 83225 -658
rect 83159 -676 83175 -674
rect 82902 -706 82928 -676
rect 83128 -706 83175 -676
rect 83159 -708 83175 -706
rect 83209 -708 83225 -674
rect 83159 -724 83225 -708
rect 83159 -984 83225 -968
rect 83159 -986 83175 -984
rect 82902 -1016 82928 -986
rect 83128 -1016 83175 -986
rect 83159 -1018 83175 -1016
rect 83209 -1018 83225 -984
rect 83159 -1034 83225 -1018
<< polycont >>
rect 2788 28362 2822 28396
rect 2788 28052 2822 28086
rect 3605 28362 3639 28396
rect 3605 28052 3639 28086
rect 7778 28362 7812 28396
rect 7778 28052 7812 28086
rect 8595 28362 8629 28396
rect 8595 28052 8629 28086
rect 12768 28362 12802 28396
rect 12768 28052 12802 28086
rect 13585 28362 13619 28396
rect 13585 28052 13619 28086
rect 17758 28362 17792 28396
rect 17758 28052 17792 28086
rect 18575 28362 18609 28396
rect 18575 28052 18609 28086
rect 22748 28362 22782 28396
rect 22748 28052 22782 28086
rect 23565 28362 23599 28396
rect 23565 28052 23599 28086
rect 27738 28362 27772 28396
rect 27738 28052 27772 28086
rect 28555 28362 28589 28396
rect 28555 28052 28589 28086
rect 32728 28362 32762 28396
rect 32728 28052 32762 28086
rect 33545 28362 33579 28396
rect 33545 28052 33579 28086
rect 37718 28362 37752 28396
rect 37718 28052 37752 28086
rect 38535 28362 38569 28396
rect 38535 28052 38569 28086
rect 42708 28362 42742 28396
rect 42708 28052 42742 28086
rect 43525 28362 43559 28396
rect 43525 28052 43559 28086
rect 47698 28362 47732 28396
rect 47698 28052 47732 28086
rect 48515 28362 48549 28396
rect 48515 28052 48549 28086
rect 52688 28362 52722 28396
rect 52688 28052 52722 28086
rect 53505 28362 53539 28396
rect 53505 28052 53539 28086
rect 57678 28362 57712 28396
rect 57678 28052 57712 28086
rect 58495 28362 58529 28396
rect 58495 28052 58529 28086
rect 62668 28362 62702 28396
rect 62668 28052 62702 28086
rect 63485 28362 63519 28396
rect 63485 28052 63519 28086
rect 67658 28362 67692 28396
rect 67658 28052 67692 28086
rect 68475 28362 68509 28396
rect 68475 28052 68509 28086
rect 72648 28362 72682 28396
rect 72648 28052 72682 28086
rect 73465 28362 73499 28396
rect 73465 28052 73499 28086
rect 77638 28362 77672 28396
rect 77638 28052 77672 28086
rect 78455 28362 78489 28396
rect 78455 28052 78489 28086
rect 82358 28362 82392 28396
rect 82358 28052 82392 28086
rect 83175 28362 83209 28396
rect 83175 28052 83209 28086
rect 82358 26652 82392 26686
rect 82358 26342 82392 26376
rect 83175 26652 83209 26686
rect 83175 26342 83209 26376
rect 82358 24942 82392 24976
rect 82358 24632 82392 24666
rect 83175 24942 83209 24976
rect 83175 24632 83209 24666
rect -1932 23232 -1898 23266
rect -1932 22922 -1898 22956
rect -1115 23232 -1081 23266
rect -1115 22922 -1081 22956
rect 82358 23232 82392 23266
rect 82358 22922 82392 22956
rect 83175 23232 83209 23266
rect 83175 22922 83209 22956
rect -1932 21522 -1898 21556
rect -1932 21212 -1898 21246
rect -1115 21522 -1081 21556
rect -1115 21212 -1081 21246
rect 82358 21522 82392 21556
rect 82358 21212 82392 21246
rect 83175 21522 83209 21556
rect 83175 21212 83209 21246
rect -1932 19812 -1898 19846
rect -1932 19502 -1898 19536
rect -1115 19812 -1081 19846
rect -1115 19502 -1081 19536
rect 82358 19812 82392 19846
rect 82358 19502 82392 19536
rect 83175 19812 83209 19846
rect 83175 19502 83209 19536
rect -1932 18102 -1898 18136
rect -1932 17792 -1898 17826
rect -1115 18102 -1081 18136
rect -1115 17792 -1081 17826
rect 82358 18102 82392 18136
rect 82358 17792 82392 17826
rect 83175 18102 83209 18136
rect 83175 17792 83209 17826
rect -1932 16392 -1898 16426
rect -1932 16082 -1898 16116
rect -1115 16392 -1081 16426
rect -1115 16082 -1081 16116
rect 82358 16392 82392 16426
rect 82358 16082 82392 16116
rect 83175 16392 83209 16426
rect 83175 16082 83209 16116
rect -1932 14682 -1898 14716
rect -1932 14372 -1898 14406
rect -1115 14682 -1081 14716
rect -1115 14372 -1081 14406
rect 82358 14682 82392 14716
rect 82358 14372 82392 14406
rect 83175 14682 83209 14716
rect 83175 14372 83209 14406
rect -1932 12972 -1898 13006
rect -1932 12662 -1898 12696
rect -1115 12972 -1081 13006
rect -1115 12662 -1081 12696
rect 82358 12972 82392 13006
rect 82358 12662 82392 12696
rect 83175 12972 83209 13006
rect 83175 12662 83209 12696
rect -1932 11262 -1898 11296
rect -1932 10952 -1898 10986
rect -1115 11262 -1081 11296
rect -1115 10952 -1081 10986
rect 82358 11262 82392 11296
rect 82358 10952 82392 10986
rect 83175 11262 83209 11296
rect 83175 10952 83209 10986
rect -1932 9552 -1898 9586
rect -1932 9242 -1898 9276
rect -1115 9552 -1081 9586
rect -1115 9242 -1081 9276
rect 82358 9552 82392 9586
rect 82358 9242 82392 9276
rect 83175 9552 83209 9586
rect 83175 9242 83209 9276
rect -1932 7842 -1898 7876
rect -1932 7532 -1898 7566
rect -1115 7842 -1081 7876
rect -1115 7532 -1081 7566
rect 82358 7842 82392 7876
rect 82358 7532 82392 7566
rect 83175 7842 83209 7876
rect 83175 7532 83209 7566
rect -1932 6132 -1898 6166
rect -1932 5822 -1898 5856
rect -1115 6132 -1081 6166
rect -1115 5822 -1081 5856
rect 82358 6132 82392 6166
rect 82358 5822 82392 5856
rect 83175 6132 83209 6166
rect 83175 5822 83209 5856
rect -1932 4422 -1898 4456
rect -1932 4112 -1898 4146
rect -1115 4422 -1081 4456
rect -1115 4112 -1081 4146
rect 82358 4422 82392 4456
rect 82358 4112 82392 4146
rect 83175 4422 83209 4456
rect 83175 4112 83209 4146
rect -1932 2712 -1898 2746
rect -1932 2402 -1898 2436
rect -1115 2712 -1081 2746
rect -1115 2402 -1081 2436
rect 82358 2712 82392 2746
rect 82358 2402 82392 2436
rect 83175 2712 83209 2746
rect 83175 2402 83209 2436
rect -1932 1002 -1898 1036
rect -1932 692 -1898 726
rect -1115 1002 -1081 1036
rect -1115 692 -1081 726
rect 82358 1002 82392 1036
rect 82358 692 82392 726
rect 83175 1002 83209 1036
rect 83175 692 83209 726
rect -1932 -708 -1898 -674
rect -1932 -1018 -1898 -984
rect -1115 -708 -1081 -674
rect -1115 -1018 -1081 -984
rect 2788 -708 2822 -674
rect 2788 -1018 2822 -984
rect 3605 -708 3639 -674
rect 3605 -1018 3639 -984
rect 7778 -708 7812 -674
rect 7778 -1018 7812 -984
rect 8595 -708 8629 -674
rect 8595 -1018 8629 -984
rect 12768 -708 12802 -674
rect 12768 -1018 12802 -984
rect 13585 -708 13619 -674
rect 13585 -1018 13619 -984
rect 17758 -708 17792 -674
rect 17758 -1018 17792 -984
rect 18575 -708 18609 -674
rect 18575 -1018 18609 -984
rect 22748 -708 22782 -674
rect 22748 -1018 22782 -984
rect 23565 -708 23599 -674
rect 23565 -1018 23599 -984
rect 27738 -708 27772 -674
rect 27738 -1018 27772 -984
rect 28555 -708 28589 -674
rect 28555 -1018 28589 -984
rect 32728 -708 32762 -674
rect 32728 -1018 32762 -984
rect 33545 -708 33579 -674
rect 33545 -1018 33579 -984
rect 37718 -708 37752 -674
rect 37718 -1018 37752 -984
rect 38535 -708 38569 -674
rect 38535 -1018 38569 -984
rect 42708 -708 42742 -674
rect 42708 -1018 42742 -984
rect 43525 -708 43559 -674
rect 43525 -1018 43559 -984
rect 47698 -708 47732 -674
rect 47698 -1018 47732 -984
rect 48515 -708 48549 -674
rect 48515 -1018 48549 -984
rect 52688 -708 52722 -674
rect 52688 -1018 52722 -984
rect 53505 -708 53539 -674
rect 53505 -1018 53539 -984
rect 57678 -708 57712 -674
rect 57678 -1018 57712 -984
rect 58495 -708 58529 -674
rect 58495 -1018 58529 -984
rect 62668 -708 62702 -674
rect 62668 -1018 62702 -984
rect 63485 -708 63519 -674
rect 63485 -1018 63519 -984
rect 67658 -708 67692 -674
rect 67658 -1018 67692 -984
rect 68475 -708 68509 -674
rect 68475 -1018 68509 -984
rect 72648 -708 72682 -674
rect 72648 -1018 72682 -984
rect 73465 -708 73499 -674
rect 73465 -1018 73499 -984
rect 77638 -708 77672 -674
rect 77638 -1018 77672 -984
rect 78455 -708 78489 -674
rect 78455 -1018 78489 -984
rect 82358 -708 82392 -674
rect 82358 -1018 82392 -984
rect 83175 -708 83209 -674
rect 83175 -1018 83209 -984
<< locali >>
rect 2640 28500 2730 28630
rect 2640 28260 2660 28500
rect 2700 28458 2730 28500
rect 2720 28300 2730 28458
rect 3700 28500 3790 28630
rect 3700 28458 3730 28500
rect 2788 28396 2822 28412
rect 2856 28406 2872 28440
rect 3048 28406 3064 28440
rect 3354 28406 3370 28440
rect 3546 28406 3562 28440
rect 2788 28346 2822 28362
rect 3605 28396 3639 28412
rect 2856 28318 2872 28352
rect 3048 28318 3064 28352
rect 3354 28318 3370 28352
rect 3546 28318 3562 28352
rect 3605 28346 3639 28362
rect 2700 28260 2730 28300
rect 2640 28200 2730 28260
rect 2640 27940 2660 28200
rect 2700 28148 2730 28200
rect 2720 27990 2730 28148
rect 3700 28300 3708 28458
rect 3700 28260 3730 28300
rect 3770 28260 3790 28500
rect 3700 28180 3790 28260
rect 3700 28148 3730 28180
rect 2788 28086 2822 28102
rect 2856 28096 2872 28130
rect 3048 28096 3064 28130
rect 3354 28096 3370 28130
rect 3546 28096 3562 28130
rect 2788 28036 2822 28052
rect 3605 28086 3639 28102
rect 2856 28008 2872 28042
rect 3048 28008 3064 28042
rect 3354 28008 3370 28042
rect 3546 28008 3562 28042
rect 3605 28036 3639 28052
rect 2700 27940 2730 27990
rect 2640 27820 2730 27940
rect 3700 27990 3708 28148
rect 3700 27940 3730 27990
rect 3770 27940 3790 28180
rect 3700 27820 3790 27940
rect 7630 28500 7720 28630
rect 7630 28260 7650 28500
rect 7690 28458 7720 28500
rect 7710 28300 7720 28458
rect 8690 28500 8780 28630
rect 8690 28458 8720 28500
rect 7778 28396 7812 28412
rect 7846 28406 7862 28440
rect 8038 28406 8054 28440
rect 8344 28406 8360 28440
rect 8536 28406 8552 28440
rect 7778 28346 7812 28362
rect 8595 28396 8629 28412
rect 7846 28318 7862 28352
rect 8038 28318 8054 28352
rect 8344 28318 8360 28352
rect 8536 28318 8552 28352
rect 8595 28346 8629 28362
rect 7690 28260 7720 28300
rect 7630 28200 7720 28260
rect 7630 27940 7650 28200
rect 7690 28148 7720 28200
rect 7710 27990 7720 28148
rect 8690 28300 8698 28458
rect 8690 28260 8720 28300
rect 8760 28260 8780 28500
rect 8690 28180 8780 28260
rect 8690 28148 8720 28180
rect 7778 28086 7812 28102
rect 7846 28096 7862 28130
rect 8038 28096 8054 28130
rect 8344 28096 8360 28130
rect 8536 28096 8552 28130
rect 7778 28036 7812 28052
rect 8595 28086 8629 28102
rect 7846 28008 7862 28042
rect 8038 28008 8054 28042
rect 8344 28008 8360 28042
rect 8536 28008 8552 28042
rect 8595 28036 8629 28052
rect 7690 27940 7720 27990
rect 7630 27820 7720 27940
rect 8690 27990 8698 28148
rect 8690 27940 8720 27990
rect 8760 27940 8780 28180
rect 8690 27820 8780 27940
rect 12620 28500 12710 28630
rect 12620 28260 12640 28500
rect 12680 28458 12710 28500
rect 12700 28300 12710 28458
rect 13680 28500 13770 28630
rect 13680 28458 13710 28500
rect 12768 28396 12802 28412
rect 12836 28406 12852 28440
rect 13028 28406 13044 28440
rect 13334 28406 13350 28440
rect 13526 28406 13542 28440
rect 12768 28346 12802 28362
rect 13585 28396 13619 28412
rect 12836 28318 12852 28352
rect 13028 28318 13044 28352
rect 13334 28318 13350 28352
rect 13526 28318 13542 28352
rect 13585 28346 13619 28362
rect 12680 28260 12710 28300
rect 12620 28200 12710 28260
rect 12620 27940 12640 28200
rect 12680 28148 12710 28200
rect 12700 27990 12710 28148
rect 13680 28300 13688 28458
rect 13680 28260 13710 28300
rect 13750 28260 13770 28500
rect 13680 28180 13770 28260
rect 13680 28148 13710 28180
rect 12768 28086 12802 28102
rect 12836 28096 12852 28130
rect 13028 28096 13044 28130
rect 13334 28096 13350 28130
rect 13526 28096 13542 28130
rect 12768 28036 12802 28052
rect 13585 28086 13619 28102
rect 12836 28008 12852 28042
rect 13028 28008 13044 28042
rect 13334 28008 13350 28042
rect 13526 28008 13542 28042
rect 13585 28036 13619 28052
rect 12680 27940 12710 27990
rect 12620 27820 12710 27940
rect 13680 27990 13688 28148
rect 13680 27940 13710 27990
rect 13750 27940 13770 28180
rect 13680 27820 13770 27940
rect 17610 28500 17700 28630
rect 17610 28260 17630 28500
rect 17670 28458 17700 28500
rect 17690 28300 17700 28458
rect 18670 28500 18760 28630
rect 18670 28458 18700 28500
rect 17758 28396 17792 28412
rect 17826 28406 17842 28440
rect 18018 28406 18034 28440
rect 18324 28406 18340 28440
rect 18516 28406 18532 28440
rect 17758 28346 17792 28362
rect 18575 28396 18609 28412
rect 17826 28318 17842 28352
rect 18018 28318 18034 28352
rect 18324 28318 18340 28352
rect 18516 28318 18532 28352
rect 18575 28346 18609 28362
rect 17670 28260 17700 28300
rect 17610 28200 17700 28260
rect 17610 27940 17630 28200
rect 17670 28148 17700 28200
rect 17690 27990 17700 28148
rect 18670 28300 18678 28458
rect 18670 28260 18700 28300
rect 18740 28260 18760 28500
rect 18670 28180 18760 28260
rect 18670 28148 18700 28180
rect 17758 28086 17792 28102
rect 17826 28096 17842 28130
rect 18018 28096 18034 28130
rect 18324 28096 18340 28130
rect 18516 28096 18532 28130
rect 17758 28036 17792 28052
rect 18575 28086 18609 28102
rect 17826 28008 17842 28042
rect 18018 28008 18034 28042
rect 18324 28008 18340 28042
rect 18516 28008 18532 28042
rect 18575 28036 18609 28052
rect 17670 27940 17700 27990
rect 17610 27820 17700 27940
rect 18670 27990 18678 28148
rect 18670 27940 18700 27990
rect 18740 27940 18760 28180
rect 18670 27820 18760 27940
rect 22600 28500 22690 28630
rect 22600 28260 22620 28500
rect 22660 28458 22690 28500
rect 22680 28300 22690 28458
rect 23660 28500 23750 28630
rect 23660 28458 23690 28500
rect 22748 28396 22782 28412
rect 22816 28406 22832 28440
rect 23008 28406 23024 28440
rect 23314 28406 23330 28440
rect 23506 28406 23522 28440
rect 22748 28346 22782 28362
rect 23565 28396 23599 28412
rect 22816 28318 22832 28352
rect 23008 28318 23024 28352
rect 23314 28318 23330 28352
rect 23506 28318 23522 28352
rect 23565 28346 23599 28362
rect 22660 28260 22690 28300
rect 22600 28200 22690 28260
rect 22600 27940 22620 28200
rect 22660 28148 22690 28200
rect 22680 27990 22690 28148
rect 23660 28300 23668 28458
rect 23660 28260 23690 28300
rect 23730 28260 23750 28500
rect 23660 28180 23750 28260
rect 23660 28148 23690 28180
rect 22748 28086 22782 28102
rect 22816 28096 22832 28130
rect 23008 28096 23024 28130
rect 23314 28096 23330 28130
rect 23506 28096 23522 28130
rect 22748 28036 22782 28052
rect 23565 28086 23599 28102
rect 22816 28008 22832 28042
rect 23008 28008 23024 28042
rect 23314 28008 23330 28042
rect 23506 28008 23522 28042
rect 23565 28036 23599 28052
rect 22660 27940 22690 27990
rect 22600 27820 22690 27940
rect 23660 27990 23668 28148
rect 23660 27940 23690 27990
rect 23730 27940 23750 28180
rect 23660 27820 23750 27940
rect 27590 28500 27680 28630
rect 27590 28260 27610 28500
rect 27650 28458 27680 28500
rect 27670 28300 27680 28458
rect 28650 28500 28740 28630
rect 28650 28458 28680 28500
rect 27738 28396 27772 28412
rect 27806 28406 27822 28440
rect 27998 28406 28014 28440
rect 28304 28406 28320 28440
rect 28496 28406 28512 28440
rect 27738 28346 27772 28362
rect 28555 28396 28589 28412
rect 27806 28318 27822 28352
rect 27998 28318 28014 28352
rect 28304 28318 28320 28352
rect 28496 28318 28512 28352
rect 28555 28346 28589 28362
rect 27650 28260 27680 28300
rect 27590 28200 27680 28260
rect 27590 27940 27610 28200
rect 27650 28148 27680 28200
rect 27670 27990 27680 28148
rect 28650 28300 28658 28458
rect 28650 28260 28680 28300
rect 28720 28260 28740 28500
rect 28650 28180 28740 28260
rect 28650 28148 28680 28180
rect 27738 28086 27772 28102
rect 27806 28096 27822 28130
rect 27998 28096 28014 28130
rect 28304 28096 28320 28130
rect 28496 28096 28512 28130
rect 27738 28036 27772 28052
rect 28555 28086 28589 28102
rect 27806 28008 27822 28042
rect 27998 28008 28014 28042
rect 28304 28008 28320 28042
rect 28496 28008 28512 28042
rect 28555 28036 28589 28052
rect 27650 27940 27680 27990
rect 27590 27820 27680 27940
rect 28650 27990 28658 28148
rect 28650 27940 28680 27990
rect 28720 27940 28740 28180
rect 28650 27820 28740 27940
rect 32580 28500 32670 28630
rect 32580 28260 32600 28500
rect 32640 28458 32670 28500
rect 32660 28300 32670 28458
rect 33640 28500 33730 28630
rect 33640 28458 33670 28500
rect 32728 28396 32762 28412
rect 32796 28406 32812 28440
rect 32988 28406 33004 28440
rect 33294 28406 33310 28440
rect 33486 28406 33502 28440
rect 32728 28346 32762 28362
rect 33545 28396 33579 28412
rect 32796 28318 32812 28352
rect 32988 28318 33004 28352
rect 33294 28318 33310 28352
rect 33486 28318 33502 28352
rect 33545 28346 33579 28362
rect 32640 28260 32670 28300
rect 32580 28200 32670 28260
rect 32580 27940 32600 28200
rect 32640 28148 32670 28200
rect 32660 27990 32670 28148
rect 33640 28300 33648 28458
rect 33640 28260 33670 28300
rect 33710 28260 33730 28500
rect 33640 28180 33730 28260
rect 33640 28148 33670 28180
rect 32728 28086 32762 28102
rect 32796 28096 32812 28130
rect 32988 28096 33004 28130
rect 33294 28096 33310 28130
rect 33486 28096 33502 28130
rect 32728 28036 32762 28052
rect 33545 28086 33579 28102
rect 32796 28008 32812 28042
rect 32988 28008 33004 28042
rect 33294 28008 33310 28042
rect 33486 28008 33502 28042
rect 33545 28036 33579 28052
rect 32640 27940 32670 27990
rect 32580 27820 32670 27940
rect 33640 27990 33648 28148
rect 33640 27940 33670 27990
rect 33710 27940 33730 28180
rect 33640 27820 33730 27940
rect 37570 28500 37660 28630
rect 37570 28260 37590 28500
rect 37630 28458 37660 28500
rect 37650 28300 37660 28458
rect 38630 28500 38720 28630
rect 38630 28458 38660 28500
rect 37718 28396 37752 28412
rect 37786 28406 37802 28440
rect 37978 28406 37994 28440
rect 38284 28406 38300 28440
rect 38476 28406 38492 28440
rect 37718 28346 37752 28362
rect 38535 28396 38569 28412
rect 37786 28318 37802 28352
rect 37978 28318 37994 28352
rect 38284 28318 38300 28352
rect 38476 28318 38492 28352
rect 38535 28346 38569 28362
rect 37630 28260 37660 28300
rect 37570 28200 37660 28260
rect 37570 27940 37590 28200
rect 37630 28148 37660 28200
rect 37650 27990 37660 28148
rect 38630 28300 38638 28458
rect 38630 28260 38660 28300
rect 38700 28260 38720 28500
rect 38630 28180 38720 28260
rect 38630 28148 38660 28180
rect 37718 28086 37752 28102
rect 37786 28096 37802 28130
rect 37978 28096 37994 28130
rect 38284 28096 38300 28130
rect 38476 28096 38492 28130
rect 37718 28036 37752 28052
rect 38535 28086 38569 28102
rect 37786 28008 37802 28042
rect 37978 28008 37994 28042
rect 38284 28008 38300 28042
rect 38476 28008 38492 28042
rect 38535 28036 38569 28052
rect 37630 27940 37660 27990
rect 37570 27820 37660 27940
rect 38630 27990 38638 28148
rect 38630 27940 38660 27990
rect 38700 27940 38720 28180
rect 38630 27820 38720 27940
rect 42560 28500 42650 28630
rect 42560 28260 42580 28500
rect 42620 28458 42650 28500
rect 42640 28300 42650 28458
rect 43620 28500 43710 28630
rect 43620 28458 43650 28500
rect 42708 28396 42742 28412
rect 42776 28406 42792 28440
rect 42968 28406 42984 28440
rect 43274 28406 43290 28440
rect 43466 28406 43482 28440
rect 42708 28346 42742 28362
rect 43525 28396 43559 28412
rect 42776 28318 42792 28352
rect 42968 28318 42984 28352
rect 43274 28318 43290 28352
rect 43466 28318 43482 28352
rect 43525 28346 43559 28362
rect 42620 28260 42650 28300
rect 42560 28200 42650 28260
rect 42560 27940 42580 28200
rect 42620 28148 42650 28200
rect 42640 27990 42650 28148
rect 43620 28300 43628 28458
rect 43620 28260 43650 28300
rect 43690 28260 43710 28500
rect 43620 28180 43710 28260
rect 43620 28148 43650 28180
rect 42708 28086 42742 28102
rect 42776 28096 42792 28130
rect 42968 28096 42984 28130
rect 43274 28096 43290 28130
rect 43466 28096 43482 28130
rect 42708 28036 42742 28052
rect 43525 28086 43559 28102
rect 42776 28008 42792 28042
rect 42968 28008 42984 28042
rect 43274 28008 43290 28042
rect 43466 28008 43482 28042
rect 43525 28036 43559 28052
rect 42620 27940 42650 27990
rect 42560 27820 42650 27940
rect 43620 27990 43628 28148
rect 43620 27940 43650 27990
rect 43690 27940 43710 28180
rect 43620 27820 43710 27940
rect 47550 28500 47640 28630
rect 47550 28260 47570 28500
rect 47610 28458 47640 28500
rect 47630 28300 47640 28458
rect 48610 28500 48700 28630
rect 48610 28458 48640 28500
rect 47698 28396 47732 28412
rect 47766 28406 47782 28440
rect 47958 28406 47974 28440
rect 48264 28406 48280 28440
rect 48456 28406 48472 28440
rect 47698 28346 47732 28362
rect 48515 28396 48549 28412
rect 47766 28318 47782 28352
rect 47958 28318 47974 28352
rect 48264 28318 48280 28352
rect 48456 28318 48472 28352
rect 48515 28346 48549 28362
rect 47610 28260 47640 28300
rect 47550 28200 47640 28260
rect 47550 27940 47570 28200
rect 47610 28148 47640 28200
rect 47630 27990 47640 28148
rect 48610 28300 48618 28458
rect 48610 28260 48640 28300
rect 48680 28260 48700 28500
rect 48610 28180 48700 28260
rect 48610 28148 48640 28180
rect 47698 28086 47732 28102
rect 47766 28096 47782 28130
rect 47958 28096 47974 28130
rect 48264 28096 48280 28130
rect 48456 28096 48472 28130
rect 47698 28036 47732 28052
rect 48515 28086 48549 28102
rect 47766 28008 47782 28042
rect 47958 28008 47974 28042
rect 48264 28008 48280 28042
rect 48456 28008 48472 28042
rect 48515 28036 48549 28052
rect 47610 27940 47640 27990
rect 47550 27820 47640 27940
rect 48610 27990 48618 28148
rect 48610 27940 48640 27990
rect 48680 27940 48700 28180
rect 48610 27820 48700 27940
rect 52540 28500 52630 28630
rect 52540 28260 52560 28500
rect 52600 28458 52630 28500
rect 52620 28300 52630 28458
rect 53600 28500 53690 28630
rect 53600 28458 53630 28500
rect 52688 28396 52722 28412
rect 52756 28406 52772 28440
rect 52948 28406 52964 28440
rect 53254 28406 53270 28440
rect 53446 28406 53462 28440
rect 52688 28346 52722 28362
rect 53505 28396 53539 28412
rect 52756 28318 52772 28352
rect 52948 28318 52964 28352
rect 53254 28318 53270 28352
rect 53446 28318 53462 28352
rect 53505 28346 53539 28362
rect 52600 28260 52630 28300
rect 52540 28200 52630 28260
rect 52540 27940 52560 28200
rect 52600 28148 52630 28200
rect 52620 27990 52630 28148
rect 53600 28300 53608 28458
rect 53600 28260 53630 28300
rect 53670 28260 53690 28500
rect 53600 28180 53690 28260
rect 53600 28148 53630 28180
rect 52688 28086 52722 28102
rect 52756 28096 52772 28130
rect 52948 28096 52964 28130
rect 53254 28096 53270 28130
rect 53446 28096 53462 28130
rect 52688 28036 52722 28052
rect 53505 28086 53539 28102
rect 52756 28008 52772 28042
rect 52948 28008 52964 28042
rect 53254 28008 53270 28042
rect 53446 28008 53462 28042
rect 53505 28036 53539 28052
rect 52600 27940 52630 27990
rect 52540 27820 52630 27940
rect 53600 27990 53608 28148
rect 53600 27940 53630 27990
rect 53670 27940 53690 28180
rect 53600 27820 53690 27940
rect 57530 28500 57620 28630
rect 57530 28260 57550 28500
rect 57590 28458 57620 28500
rect 57610 28300 57620 28458
rect 58590 28500 58680 28630
rect 58590 28458 58620 28500
rect 57678 28396 57712 28412
rect 57746 28406 57762 28440
rect 57938 28406 57954 28440
rect 58244 28406 58260 28440
rect 58436 28406 58452 28440
rect 57678 28346 57712 28362
rect 58495 28396 58529 28412
rect 57746 28318 57762 28352
rect 57938 28318 57954 28352
rect 58244 28318 58260 28352
rect 58436 28318 58452 28352
rect 58495 28346 58529 28362
rect 57590 28260 57620 28300
rect 57530 28200 57620 28260
rect 57530 27940 57550 28200
rect 57590 28148 57620 28200
rect 57610 27990 57620 28148
rect 58590 28300 58598 28458
rect 58590 28260 58620 28300
rect 58660 28260 58680 28500
rect 58590 28180 58680 28260
rect 58590 28148 58620 28180
rect 57678 28086 57712 28102
rect 57746 28096 57762 28130
rect 57938 28096 57954 28130
rect 58244 28096 58260 28130
rect 58436 28096 58452 28130
rect 57678 28036 57712 28052
rect 58495 28086 58529 28102
rect 57746 28008 57762 28042
rect 57938 28008 57954 28042
rect 58244 28008 58260 28042
rect 58436 28008 58452 28042
rect 58495 28036 58529 28052
rect 57590 27940 57620 27990
rect 57530 27820 57620 27940
rect 58590 27990 58598 28148
rect 58590 27940 58620 27990
rect 58660 27940 58680 28180
rect 58590 27820 58680 27940
rect 62520 28500 62610 28630
rect 62520 28260 62540 28500
rect 62580 28458 62610 28500
rect 62600 28300 62610 28458
rect 63580 28500 63670 28630
rect 63580 28458 63610 28500
rect 62668 28396 62702 28412
rect 62736 28406 62752 28440
rect 62928 28406 62944 28440
rect 63234 28406 63250 28440
rect 63426 28406 63442 28440
rect 62668 28346 62702 28362
rect 63485 28396 63519 28412
rect 62736 28318 62752 28352
rect 62928 28318 62944 28352
rect 63234 28318 63250 28352
rect 63426 28318 63442 28352
rect 63485 28346 63519 28362
rect 62580 28260 62610 28300
rect 62520 28200 62610 28260
rect 62520 27940 62540 28200
rect 62580 28148 62610 28200
rect 62600 27990 62610 28148
rect 63580 28300 63588 28458
rect 63580 28260 63610 28300
rect 63650 28260 63670 28500
rect 63580 28180 63670 28260
rect 63580 28148 63610 28180
rect 62668 28086 62702 28102
rect 62736 28096 62752 28130
rect 62928 28096 62944 28130
rect 63234 28096 63250 28130
rect 63426 28096 63442 28130
rect 62668 28036 62702 28052
rect 63485 28086 63519 28102
rect 62736 28008 62752 28042
rect 62928 28008 62944 28042
rect 63234 28008 63250 28042
rect 63426 28008 63442 28042
rect 63485 28036 63519 28052
rect 62580 27940 62610 27990
rect 62520 27820 62610 27940
rect 63580 27990 63588 28148
rect 63580 27940 63610 27990
rect 63650 27940 63670 28180
rect 63580 27820 63670 27940
rect 67510 28500 67600 28630
rect 67510 28260 67530 28500
rect 67570 28458 67600 28500
rect 67590 28300 67600 28458
rect 68570 28500 68660 28630
rect 68570 28458 68600 28500
rect 67658 28396 67692 28412
rect 67726 28406 67742 28440
rect 67918 28406 67934 28440
rect 68224 28406 68240 28440
rect 68416 28406 68432 28440
rect 67658 28346 67692 28362
rect 68475 28396 68509 28412
rect 67726 28318 67742 28352
rect 67918 28318 67934 28352
rect 68224 28318 68240 28352
rect 68416 28318 68432 28352
rect 68475 28346 68509 28362
rect 67570 28260 67600 28300
rect 67510 28200 67600 28260
rect 67510 27940 67530 28200
rect 67570 28148 67600 28200
rect 67590 27990 67600 28148
rect 68570 28300 68578 28458
rect 68570 28260 68600 28300
rect 68640 28260 68660 28500
rect 68570 28180 68660 28260
rect 68570 28148 68600 28180
rect 67658 28086 67692 28102
rect 67726 28096 67742 28130
rect 67918 28096 67934 28130
rect 68224 28096 68240 28130
rect 68416 28096 68432 28130
rect 67658 28036 67692 28052
rect 68475 28086 68509 28102
rect 67726 28008 67742 28042
rect 67918 28008 67934 28042
rect 68224 28008 68240 28042
rect 68416 28008 68432 28042
rect 68475 28036 68509 28052
rect 67570 27940 67600 27990
rect 67510 27820 67600 27940
rect 68570 27990 68578 28148
rect 68570 27940 68600 27990
rect 68640 27940 68660 28180
rect 68570 27820 68660 27940
rect 72500 28500 72590 28630
rect 72500 28260 72520 28500
rect 72560 28458 72590 28500
rect 72580 28300 72590 28458
rect 73560 28500 73650 28630
rect 73560 28458 73590 28500
rect 72648 28396 72682 28412
rect 72716 28406 72732 28440
rect 72908 28406 72924 28440
rect 73214 28406 73230 28440
rect 73406 28406 73422 28440
rect 72648 28346 72682 28362
rect 73465 28396 73499 28412
rect 72716 28318 72732 28352
rect 72908 28318 72924 28352
rect 73214 28318 73230 28352
rect 73406 28318 73422 28352
rect 73465 28346 73499 28362
rect 72560 28260 72590 28300
rect 72500 28200 72590 28260
rect 72500 27940 72520 28200
rect 72560 28148 72590 28200
rect 72580 27990 72590 28148
rect 73560 28300 73568 28458
rect 73560 28260 73590 28300
rect 73630 28260 73650 28500
rect 73560 28180 73650 28260
rect 73560 28148 73590 28180
rect 72648 28086 72682 28102
rect 72716 28096 72732 28130
rect 72908 28096 72924 28130
rect 73214 28096 73230 28130
rect 73406 28096 73422 28130
rect 72648 28036 72682 28052
rect 73465 28086 73499 28102
rect 72716 28008 72732 28042
rect 72908 28008 72924 28042
rect 73214 28008 73230 28042
rect 73406 28008 73422 28042
rect 73465 28036 73499 28052
rect 72560 27940 72590 27990
rect 72500 27820 72590 27940
rect 73560 27990 73568 28148
rect 73560 27940 73590 27990
rect 73630 27940 73650 28180
rect 73560 27820 73650 27940
rect 77490 28500 77580 28630
rect 77490 28260 77510 28500
rect 77550 28458 77580 28500
rect 77570 28300 77580 28458
rect 78550 28500 78640 28630
rect 78550 28458 78580 28500
rect 77638 28396 77672 28412
rect 77706 28406 77722 28440
rect 77898 28406 77914 28440
rect 78204 28406 78220 28440
rect 78396 28406 78412 28440
rect 77638 28346 77672 28362
rect 78455 28396 78489 28412
rect 77706 28318 77722 28352
rect 77898 28318 77914 28352
rect 78204 28318 78220 28352
rect 78396 28318 78412 28352
rect 78455 28346 78489 28362
rect 77550 28260 77580 28300
rect 77490 28200 77580 28260
rect 77490 27940 77510 28200
rect 77550 28148 77580 28200
rect 77570 27990 77580 28148
rect 78550 28300 78558 28458
rect 78550 28260 78580 28300
rect 78620 28260 78640 28500
rect 78550 28180 78640 28260
rect 78550 28148 78580 28180
rect 77638 28086 77672 28102
rect 77706 28096 77722 28130
rect 77898 28096 77914 28130
rect 78204 28096 78220 28130
rect 78396 28096 78412 28130
rect 77638 28036 77672 28052
rect 78455 28086 78489 28102
rect 77706 28008 77722 28042
rect 77898 28008 77914 28042
rect 78204 28008 78220 28042
rect 78396 28008 78412 28042
rect 78455 28036 78489 28052
rect 77550 27940 77580 27990
rect 77490 27820 77580 27940
rect 78550 27990 78558 28148
rect 78550 27940 78580 27990
rect 78620 27940 78640 28180
rect 78550 27820 78640 27940
rect 82210 28500 82300 28630
rect 82210 28260 82230 28500
rect 82270 28458 82300 28500
rect 82290 28300 82300 28458
rect 83270 28500 83360 28630
rect 83270 28458 83300 28500
rect 82358 28396 82392 28412
rect 82426 28406 82442 28440
rect 82618 28406 82634 28440
rect 82924 28406 82940 28440
rect 83116 28406 83132 28440
rect 82358 28346 82392 28362
rect 83175 28396 83209 28412
rect 82426 28318 82442 28352
rect 82618 28318 82634 28352
rect 82924 28318 82940 28352
rect 83116 28318 83132 28352
rect 83175 28346 83209 28362
rect 82270 28260 82300 28300
rect 82210 28200 82300 28260
rect 82210 27940 82230 28200
rect 82270 28148 82300 28200
rect 82290 27990 82300 28148
rect 83270 28300 83278 28458
rect 83270 28260 83300 28300
rect 83340 28260 83360 28500
rect 83270 28180 83360 28260
rect 83270 28148 83300 28180
rect 82358 28086 82392 28102
rect 82426 28096 82442 28130
rect 82618 28096 82634 28130
rect 82924 28096 82940 28130
rect 83116 28096 83132 28130
rect 82358 28036 82392 28052
rect 83175 28086 83209 28102
rect 82426 28008 82442 28042
rect 82618 28008 82634 28042
rect 82924 28008 82940 28042
rect 83116 28008 83132 28042
rect 83175 28036 83209 28052
rect 82270 27940 82300 27990
rect 82210 27820 82300 27940
rect 83270 27990 83278 28148
rect 83270 27940 83300 27990
rect 83340 27940 83360 28180
rect 83270 27820 83360 27940
rect 82210 26790 82300 26920
rect 82210 26550 82230 26790
rect 82270 26748 82300 26790
rect 82290 26590 82300 26748
rect 83270 26790 83360 26920
rect 83270 26748 83300 26790
rect 82358 26686 82392 26702
rect 82426 26696 82442 26730
rect 82618 26696 82634 26730
rect 82924 26696 82940 26730
rect 83116 26696 83132 26730
rect 82358 26636 82392 26652
rect 83175 26686 83209 26702
rect 82426 26608 82442 26642
rect 82618 26608 82634 26642
rect 82924 26608 82940 26642
rect 83116 26608 83132 26642
rect 83175 26636 83209 26652
rect 82270 26550 82300 26590
rect 82210 26490 82300 26550
rect 82210 26230 82230 26490
rect 82270 26438 82300 26490
rect 82290 26280 82300 26438
rect 83270 26590 83278 26748
rect 83270 26550 83300 26590
rect 83340 26550 83360 26790
rect 83270 26470 83360 26550
rect 83270 26438 83300 26470
rect 82358 26376 82392 26392
rect 82426 26386 82442 26420
rect 82618 26386 82634 26420
rect 82924 26386 82940 26420
rect 83116 26386 83132 26420
rect 82358 26326 82392 26342
rect 83175 26376 83209 26392
rect 82426 26298 82442 26332
rect 82618 26298 82634 26332
rect 82924 26298 82940 26332
rect 83116 26298 83132 26332
rect 83175 26326 83209 26342
rect 82270 26230 82300 26280
rect 82210 26110 82300 26230
rect 83270 26280 83278 26438
rect 83270 26230 83300 26280
rect 83340 26230 83360 26470
rect 83270 26110 83360 26230
rect 82210 25080 82300 25210
rect 82210 24840 82230 25080
rect 82270 25038 82300 25080
rect 82290 24880 82300 25038
rect 83270 25080 83360 25210
rect 83270 25038 83300 25080
rect 82358 24976 82392 24992
rect 82426 24986 82442 25020
rect 82618 24986 82634 25020
rect 82924 24986 82940 25020
rect 83116 24986 83132 25020
rect 82358 24926 82392 24942
rect 83175 24976 83209 24992
rect 82426 24898 82442 24932
rect 82618 24898 82634 24932
rect 82924 24898 82940 24932
rect 83116 24898 83132 24932
rect 83175 24926 83209 24942
rect 82270 24840 82300 24880
rect 82210 24780 82300 24840
rect 82210 24520 82230 24780
rect 82270 24728 82300 24780
rect 82290 24570 82300 24728
rect 83270 24880 83278 25038
rect 83270 24840 83300 24880
rect 83340 24840 83360 25080
rect 83270 24760 83360 24840
rect 83270 24728 83300 24760
rect 82358 24666 82392 24682
rect 82426 24676 82442 24710
rect 82618 24676 82634 24710
rect 82924 24676 82940 24710
rect 83116 24676 83132 24710
rect 82358 24616 82392 24632
rect 83175 24666 83209 24682
rect 82426 24588 82442 24622
rect 82618 24588 82634 24622
rect 82924 24588 82940 24622
rect 83116 24588 83132 24622
rect 83175 24616 83209 24632
rect 82270 24520 82300 24570
rect 82210 24400 82300 24520
rect 83270 24570 83278 24728
rect 83270 24520 83300 24570
rect 83340 24520 83360 24760
rect 83270 24400 83360 24520
rect -2080 23370 -1990 23500
rect -2080 23130 -2060 23370
rect -2020 23328 -1990 23370
rect -2000 23170 -1990 23328
rect -1020 23370 -930 23500
rect -1020 23328 -990 23370
rect -1932 23266 -1898 23282
rect -1864 23276 -1848 23310
rect -1672 23276 -1656 23310
rect -1366 23276 -1350 23310
rect -1174 23276 -1158 23310
rect -1932 23216 -1898 23232
rect -1115 23266 -1081 23282
rect -1864 23188 -1848 23222
rect -1672 23188 -1656 23222
rect -1366 23188 -1350 23222
rect -1174 23188 -1158 23222
rect -1115 23216 -1081 23232
rect -2020 23130 -1990 23170
rect -2080 23070 -1990 23130
rect -2080 22810 -2060 23070
rect -2020 23018 -1990 23070
rect -2000 22860 -1990 23018
rect -1020 23170 -1012 23328
rect -1020 23130 -990 23170
rect -950 23130 -930 23370
rect -1020 23050 -930 23130
rect -1020 23018 -990 23050
rect -1932 22956 -1898 22972
rect -1864 22966 -1848 23000
rect -1672 22966 -1656 23000
rect -1366 22966 -1350 23000
rect -1174 22966 -1158 23000
rect -1932 22906 -1898 22922
rect -1115 22956 -1081 22972
rect -1864 22878 -1848 22912
rect -1672 22878 -1656 22912
rect -1366 22878 -1350 22912
rect -1174 22878 -1158 22912
rect -1115 22906 -1081 22922
rect -2020 22810 -1990 22860
rect -2080 22690 -1990 22810
rect -1020 22860 -1012 23018
rect -1020 22810 -990 22860
rect -950 22810 -930 23050
rect -1020 22690 -930 22810
rect 82210 23370 82300 23500
rect 82210 23130 82230 23370
rect 82270 23328 82300 23370
rect 82290 23170 82300 23328
rect 83270 23370 83360 23500
rect 83270 23328 83300 23370
rect 82358 23266 82392 23282
rect 82426 23276 82442 23310
rect 82618 23276 82634 23310
rect 82924 23276 82940 23310
rect 83116 23276 83132 23310
rect 82358 23216 82392 23232
rect 83175 23266 83209 23282
rect 82426 23188 82442 23222
rect 82618 23188 82634 23222
rect 82924 23188 82940 23222
rect 83116 23188 83132 23222
rect 83175 23216 83209 23232
rect 82270 23130 82300 23170
rect 82210 23070 82300 23130
rect 82210 22810 82230 23070
rect 82270 23018 82300 23070
rect 82290 22860 82300 23018
rect 83270 23170 83278 23328
rect 83270 23130 83300 23170
rect 83340 23130 83360 23370
rect 83270 23050 83360 23130
rect 83270 23018 83300 23050
rect 82358 22956 82392 22972
rect 82426 22966 82442 23000
rect 82618 22966 82634 23000
rect 82924 22966 82940 23000
rect 83116 22966 83132 23000
rect 82358 22906 82392 22922
rect 83175 22956 83209 22972
rect 82426 22878 82442 22912
rect 82618 22878 82634 22912
rect 82924 22878 82940 22912
rect 83116 22878 83132 22912
rect 83175 22906 83209 22922
rect 82270 22810 82300 22860
rect 82210 22690 82300 22810
rect 83270 22860 83278 23018
rect 83270 22810 83300 22860
rect 83340 22810 83360 23050
rect 83270 22690 83360 22810
rect -2080 21660 -1990 21790
rect -2080 21420 -2060 21660
rect -2020 21618 -1990 21660
rect -2000 21460 -1990 21618
rect -1020 21660 -930 21790
rect -1020 21618 -990 21660
rect -1932 21556 -1898 21572
rect -1864 21566 -1848 21600
rect -1672 21566 -1656 21600
rect -1366 21566 -1350 21600
rect -1174 21566 -1158 21600
rect -1932 21506 -1898 21522
rect -1115 21556 -1081 21572
rect -1864 21478 -1848 21512
rect -1672 21478 -1656 21512
rect -1366 21478 -1350 21512
rect -1174 21478 -1158 21512
rect -1115 21506 -1081 21522
rect -2020 21420 -1990 21460
rect -2080 21360 -1990 21420
rect -2080 21100 -2060 21360
rect -2020 21308 -1990 21360
rect -2000 21150 -1990 21308
rect -1020 21460 -1012 21618
rect -1020 21420 -990 21460
rect -950 21420 -930 21660
rect -1020 21340 -930 21420
rect -1020 21308 -990 21340
rect -1932 21246 -1898 21262
rect -1864 21256 -1848 21290
rect -1672 21256 -1656 21290
rect -1366 21256 -1350 21290
rect -1174 21256 -1158 21290
rect -1932 21196 -1898 21212
rect -1115 21246 -1081 21262
rect -1864 21168 -1848 21202
rect -1672 21168 -1656 21202
rect -1366 21168 -1350 21202
rect -1174 21168 -1158 21202
rect -1115 21196 -1081 21212
rect -2020 21100 -1990 21150
rect -2080 20980 -1990 21100
rect -1020 21150 -1012 21308
rect -1020 21100 -990 21150
rect -950 21100 -930 21340
rect -1020 20980 -930 21100
rect 82210 21660 82300 21790
rect 82210 21420 82230 21660
rect 82270 21618 82300 21660
rect 82290 21460 82300 21618
rect 83270 21660 83360 21790
rect 83270 21618 83300 21660
rect 82358 21556 82392 21572
rect 82426 21566 82442 21600
rect 82618 21566 82634 21600
rect 82924 21566 82940 21600
rect 83116 21566 83132 21600
rect 82358 21506 82392 21522
rect 83175 21556 83209 21572
rect 82426 21478 82442 21512
rect 82618 21478 82634 21512
rect 82924 21478 82940 21512
rect 83116 21478 83132 21512
rect 83175 21506 83209 21522
rect 82270 21420 82300 21460
rect 82210 21360 82300 21420
rect 82210 21100 82230 21360
rect 82270 21308 82300 21360
rect 82290 21150 82300 21308
rect 83270 21460 83278 21618
rect 83270 21420 83300 21460
rect 83340 21420 83360 21660
rect 83270 21340 83360 21420
rect 83270 21308 83300 21340
rect 82358 21246 82392 21262
rect 82426 21256 82442 21290
rect 82618 21256 82634 21290
rect 82924 21256 82940 21290
rect 83116 21256 83132 21290
rect 82358 21196 82392 21212
rect 83175 21246 83209 21262
rect 82426 21168 82442 21202
rect 82618 21168 82634 21202
rect 82924 21168 82940 21202
rect 83116 21168 83132 21202
rect 83175 21196 83209 21212
rect 82270 21100 82300 21150
rect 82210 20980 82300 21100
rect 83270 21150 83278 21308
rect 83270 21100 83300 21150
rect 83340 21100 83360 21340
rect 83270 20980 83360 21100
rect -2080 19950 -1990 20080
rect -2080 19710 -2060 19950
rect -2020 19908 -1990 19950
rect -2000 19750 -1990 19908
rect -1020 19950 -930 20080
rect -1020 19908 -990 19950
rect -1932 19846 -1898 19862
rect -1864 19856 -1848 19890
rect -1672 19856 -1656 19890
rect -1366 19856 -1350 19890
rect -1174 19856 -1158 19890
rect -1932 19796 -1898 19812
rect -1115 19846 -1081 19862
rect -1864 19768 -1848 19802
rect -1672 19768 -1656 19802
rect -1366 19768 -1350 19802
rect -1174 19768 -1158 19802
rect -1115 19796 -1081 19812
rect -2020 19710 -1990 19750
rect -2080 19650 -1990 19710
rect -2080 19390 -2060 19650
rect -2020 19598 -1990 19650
rect -2000 19440 -1990 19598
rect -1020 19750 -1012 19908
rect -1020 19710 -990 19750
rect -950 19710 -930 19950
rect -1020 19630 -930 19710
rect -1020 19598 -990 19630
rect -1932 19536 -1898 19552
rect -1864 19546 -1848 19580
rect -1672 19546 -1656 19580
rect -1366 19546 -1350 19580
rect -1174 19546 -1158 19580
rect -1932 19486 -1898 19502
rect -1115 19536 -1081 19552
rect -1864 19458 -1848 19492
rect -1672 19458 -1656 19492
rect -1366 19458 -1350 19492
rect -1174 19458 -1158 19492
rect -1115 19486 -1081 19502
rect -2020 19390 -1990 19440
rect -2080 19270 -1990 19390
rect -1020 19440 -1012 19598
rect -1020 19390 -990 19440
rect -950 19390 -930 19630
rect -1020 19270 -930 19390
rect 82210 19950 82300 20080
rect 82210 19710 82230 19950
rect 82270 19908 82300 19950
rect 82290 19750 82300 19908
rect 83270 19950 83360 20080
rect 83270 19908 83300 19950
rect 82358 19846 82392 19862
rect 82426 19856 82442 19890
rect 82618 19856 82634 19890
rect 82924 19856 82940 19890
rect 83116 19856 83132 19890
rect 82358 19796 82392 19812
rect 83175 19846 83209 19862
rect 82426 19768 82442 19802
rect 82618 19768 82634 19802
rect 82924 19768 82940 19802
rect 83116 19768 83132 19802
rect 83175 19796 83209 19812
rect 82270 19710 82300 19750
rect 82210 19650 82300 19710
rect 82210 19390 82230 19650
rect 82270 19598 82300 19650
rect 82290 19440 82300 19598
rect 83270 19750 83278 19908
rect 83270 19710 83300 19750
rect 83340 19710 83360 19950
rect 83270 19630 83360 19710
rect 83270 19598 83300 19630
rect 82358 19536 82392 19552
rect 82426 19546 82442 19580
rect 82618 19546 82634 19580
rect 82924 19546 82940 19580
rect 83116 19546 83132 19580
rect 82358 19486 82392 19502
rect 83175 19536 83209 19552
rect 82426 19458 82442 19492
rect 82618 19458 82634 19492
rect 82924 19458 82940 19492
rect 83116 19458 83132 19492
rect 83175 19486 83209 19502
rect 82270 19390 82300 19440
rect 82210 19270 82300 19390
rect 83270 19440 83278 19598
rect 83270 19390 83300 19440
rect 83340 19390 83360 19630
rect 83270 19270 83360 19390
rect -2080 18240 -1990 18370
rect -2080 18000 -2060 18240
rect -2020 18198 -1990 18240
rect -2000 18040 -1990 18198
rect -1020 18240 -930 18370
rect -1020 18198 -990 18240
rect -1932 18136 -1898 18152
rect -1864 18146 -1848 18180
rect -1672 18146 -1656 18180
rect -1366 18146 -1350 18180
rect -1174 18146 -1158 18180
rect -1932 18086 -1898 18102
rect -1115 18136 -1081 18152
rect -1864 18058 -1848 18092
rect -1672 18058 -1656 18092
rect -1366 18058 -1350 18092
rect -1174 18058 -1158 18092
rect -1115 18086 -1081 18102
rect -2020 18000 -1990 18040
rect -2080 17940 -1990 18000
rect -2080 17680 -2060 17940
rect -2020 17888 -1990 17940
rect -2000 17730 -1990 17888
rect -1020 18040 -1012 18198
rect -1020 18000 -990 18040
rect -950 18000 -930 18240
rect -1020 17920 -930 18000
rect -1020 17888 -990 17920
rect -1932 17826 -1898 17842
rect -1864 17836 -1848 17870
rect -1672 17836 -1656 17870
rect -1366 17836 -1350 17870
rect -1174 17836 -1158 17870
rect -1932 17776 -1898 17792
rect -1115 17826 -1081 17842
rect -1864 17748 -1848 17782
rect -1672 17748 -1656 17782
rect -1366 17748 -1350 17782
rect -1174 17748 -1158 17782
rect -1115 17776 -1081 17792
rect -2020 17680 -1990 17730
rect -2080 17560 -1990 17680
rect -1020 17730 -1012 17888
rect -1020 17680 -990 17730
rect -950 17680 -930 17920
rect -1020 17560 -930 17680
rect 82210 18240 82300 18370
rect 82210 18000 82230 18240
rect 82270 18198 82300 18240
rect 82290 18040 82300 18198
rect 83270 18240 83360 18370
rect 83270 18198 83300 18240
rect 82358 18136 82392 18152
rect 82426 18146 82442 18180
rect 82618 18146 82634 18180
rect 82924 18146 82940 18180
rect 83116 18146 83132 18180
rect 82358 18086 82392 18102
rect 83175 18136 83209 18152
rect 82426 18058 82442 18092
rect 82618 18058 82634 18092
rect 82924 18058 82940 18092
rect 83116 18058 83132 18092
rect 83175 18086 83209 18102
rect 82270 18000 82300 18040
rect 82210 17940 82300 18000
rect 82210 17680 82230 17940
rect 82270 17888 82300 17940
rect 82290 17730 82300 17888
rect 83270 18040 83278 18198
rect 83270 18000 83300 18040
rect 83340 18000 83360 18240
rect 83270 17920 83360 18000
rect 83270 17888 83300 17920
rect 82358 17826 82392 17842
rect 82426 17836 82442 17870
rect 82618 17836 82634 17870
rect 82924 17836 82940 17870
rect 83116 17836 83132 17870
rect 82358 17776 82392 17792
rect 83175 17826 83209 17842
rect 82426 17748 82442 17782
rect 82618 17748 82634 17782
rect 82924 17748 82940 17782
rect 83116 17748 83132 17782
rect 83175 17776 83209 17792
rect 82270 17680 82300 17730
rect 82210 17560 82300 17680
rect 83270 17730 83278 17888
rect 83270 17680 83300 17730
rect 83340 17680 83360 17920
rect 83270 17560 83360 17680
rect -2080 16530 -1990 16660
rect -2080 16290 -2060 16530
rect -2020 16488 -1990 16530
rect -2000 16330 -1990 16488
rect -1020 16530 -930 16660
rect -1020 16488 -990 16530
rect -1932 16426 -1898 16442
rect -1864 16436 -1848 16470
rect -1672 16436 -1656 16470
rect -1366 16436 -1350 16470
rect -1174 16436 -1158 16470
rect -1932 16376 -1898 16392
rect -1115 16426 -1081 16442
rect -1864 16348 -1848 16382
rect -1672 16348 -1656 16382
rect -1366 16348 -1350 16382
rect -1174 16348 -1158 16382
rect -1115 16376 -1081 16392
rect -2020 16290 -1990 16330
rect -2080 16230 -1990 16290
rect -2080 15970 -2060 16230
rect -2020 16178 -1990 16230
rect -2000 16020 -1990 16178
rect -1020 16330 -1012 16488
rect -1020 16290 -990 16330
rect -950 16290 -930 16530
rect -1020 16210 -930 16290
rect -1020 16178 -990 16210
rect -1932 16116 -1898 16132
rect -1864 16126 -1848 16160
rect -1672 16126 -1656 16160
rect -1366 16126 -1350 16160
rect -1174 16126 -1158 16160
rect -1932 16066 -1898 16082
rect -1115 16116 -1081 16132
rect -1864 16038 -1848 16072
rect -1672 16038 -1656 16072
rect -1366 16038 -1350 16072
rect -1174 16038 -1158 16072
rect -1115 16066 -1081 16082
rect -2020 15970 -1990 16020
rect -2080 15850 -1990 15970
rect -1020 16020 -1012 16178
rect -1020 15970 -990 16020
rect -950 15970 -930 16210
rect -1020 15850 -930 15970
rect 82210 16530 82300 16660
rect 82210 16290 82230 16530
rect 82270 16488 82300 16530
rect 82290 16330 82300 16488
rect 83270 16530 83360 16660
rect 83270 16488 83300 16530
rect 82358 16426 82392 16442
rect 82426 16436 82442 16470
rect 82618 16436 82634 16470
rect 82924 16436 82940 16470
rect 83116 16436 83132 16470
rect 82358 16376 82392 16392
rect 83175 16426 83209 16442
rect 82426 16348 82442 16382
rect 82618 16348 82634 16382
rect 82924 16348 82940 16382
rect 83116 16348 83132 16382
rect 83175 16376 83209 16392
rect 82270 16290 82300 16330
rect 82210 16230 82300 16290
rect 82210 15970 82230 16230
rect 82270 16178 82300 16230
rect 82290 16020 82300 16178
rect 83270 16330 83278 16488
rect 83270 16290 83300 16330
rect 83340 16290 83360 16530
rect 83270 16210 83360 16290
rect 83270 16178 83300 16210
rect 82358 16116 82392 16132
rect 82426 16126 82442 16160
rect 82618 16126 82634 16160
rect 82924 16126 82940 16160
rect 83116 16126 83132 16160
rect 82358 16066 82392 16082
rect 83175 16116 83209 16132
rect 82426 16038 82442 16072
rect 82618 16038 82634 16072
rect 82924 16038 82940 16072
rect 83116 16038 83132 16072
rect 83175 16066 83209 16082
rect 82270 15970 82300 16020
rect 82210 15850 82300 15970
rect 83270 16020 83278 16178
rect 83270 15970 83300 16020
rect 83340 15970 83360 16210
rect 83270 15850 83360 15970
rect -2080 14820 -1990 14950
rect -2080 14580 -2060 14820
rect -2020 14778 -1990 14820
rect -2000 14620 -1990 14778
rect -1020 14820 -930 14950
rect -1020 14778 -990 14820
rect -1932 14716 -1898 14732
rect -1864 14726 -1848 14760
rect -1672 14726 -1656 14760
rect -1366 14726 -1350 14760
rect -1174 14726 -1158 14760
rect -1932 14666 -1898 14682
rect -1115 14716 -1081 14732
rect -1864 14638 -1848 14672
rect -1672 14638 -1656 14672
rect -1366 14638 -1350 14672
rect -1174 14638 -1158 14672
rect -1115 14666 -1081 14682
rect -2020 14580 -1990 14620
rect -2080 14520 -1990 14580
rect -2080 14260 -2060 14520
rect -2020 14468 -1990 14520
rect -2000 14310 -1990 14468
rect -1020 14620 -1012 14778
rect -1020 14580 -990 14620
rect -950 14580 -930 14820
rect -1020 14500 -930 14580
rect -1020 14468 -990 14500
rect -1932 14406 -1898 14422
rect -1864 14416 -1848 14450
rect -1672 14416 -1656 14450
rect -1366 14416 -1350 14450
rect -1174 14416 -1158 14450
rect -1932 14356 -1898 14372
rect -1115 14406 -1081 14422
rect -1864 14328 -1848 14362
rect -1672 14328 -1656 14362
rect -1366 14328 -1350 14362
rect -1174 14328 -1158 14362
rect -1115 14356 -1081 14372
rect -2020 14260 -1990 14310
rect -2080 14140 -1990 14260
rect -1020 14310 -1012 14468
rect -1020 14260 -990 14310
rect -950 14260 -930 14500
rect -1020 14140 -930 14260
rect 82210 14820 82300 14950
rect 82210 14580 82230 14820
rect 82270 14778 82300 14820
rect 82290 14620 82300 14778
rect 83270 14820 83360 14950
rect 83270 14778 83300 14820
rect 82358 14716 82392 14732
rect 82426 14726 82442 14760
rect 82618 14726 82634 14760
rect 82924 14726 82940 14760
rect 83116 14726 83132 14760
rect 82358 14666 82392 14682
rect 83175 14716 83209 14732
rect 82426 14638 82442 14672
rect 82618 14638 82634 14672
rect 82924 14638 82940 14672
rect 83116 14638 83132 14672
rect 83175 14666 83209 14682
rect 82270 14580 82300 14620
rect 82210 14520 82300 14580
rect 82210 14260 82230 14520
rect 82270 14468 82300 14520
rect 82290 14310 82300 14468
rect 83270 14620 83278 14778
rect 83270 14580 83300 14620
rect 83340 14580 83360 14820
rect 83270 14500 83360 14580
rect 83270 14468 83300 14500
rect 82358 14406 82392 14422
rect 82426 14416 82442 14450
rect 82618 14416 82634 14450
rect 82924 14416 82940 14450
rect 83116 14416 83132 14450
rect 82358 14356 82392 14372
rect 83175 14406 83209 14422
rect 82426 14328 82442 14362
rect 82618 14328 82634 14362
rect 82924 14328 82940 14362
rect 83116 14328 83132 14362
rect 83175 14356 83209 14372
rect 82270 14260 82300 14310
rect 82210 14140 82300 14260
rect 83270 14310 83278 14468
rect 83270 14260 83300 14310
rect 83340 14260 83360 14500
rect 83270 14140 83360 14260
rect -2080 13110 -1990 13240
rect -2080 12870 -2060 13110
rect -2020 13068 -1990 13110
rect -2000 12910 -1990 13068
rect -1020 13110 -930 13240
rect -1020 13068 -990 13110
rect -1932 13006 -1898 13022
rect -1864 13016 -1848 13050
rect -1672 13016 -1656 13050
rect -1366 13016 -1350 13050
rect -1174 13016 -1158 13050
rect -1932 12956 -1898 12972
rect -1115 13006 -1081 13022
rect -1864 12928 -1848 12962
rect -1672 12928 -1656 12962
rect -1366 12928 -1350 12962
rect -1174 12928 -1158 12962
rect -1115 12956 -1081 12972
rect -2020 12870 -1990 12910
rect -2080 12810 -1990 12870
rect -2080 12550 -2060 12810
rect -2020 12758 -1990 12810
rect -2000 12600 -1990 12758
rect -1020 12910 -1012 13068
rect -1020 12870 -990 12910
rect -950 12870 -930 13110
rect -1020 12790 -930 12870
rect -1020 12758 -990 12790
rect -1932 12696 -1898 12712
rect -1864 12706 -1848 12740
rect -1672 12706 -1656 12740
rect -1366 12706 -1350 12740
rect -1174 12706 -1158 12740
rect -1932 12646 -1898 12662
rect -1115 12696 -1081 12712
rect -1864 12618 -1848 12652
rect -1672 12618 -1656 12652
rect -1366 12618 -1350 12652
rect -1174 12618 -1158 12652
rect -1115 12646 -1081 12662
rect -2020 12550 -1990 12600
rect -2080 12430 -1990 12550
rect -1020 12600 -1012 12758
rect -1020 12550 -990 12600
rect -950 12550 -930 12790
rect -1020 12430 -930 12550
rect 82210 13110 82300 13240
rect 82210 12870 82230 13110
rect 82270 13068 82300 13110
rect 82290 12910 82300 13068
rect 83270 13110 83360 13240
rect 83270 13068 83300 13110
rect 82358 13006 82392 13022
rect 82426 13016 82442 13050
rect 82618 13016 82634 13050
rect 82924 13016 82940 13050
rect 83116 13016 83132 13050
rect 82358 12956 82392 12972
rect 83175 13006 83209 13022
rect 82426 12928 82442 12962
rect 82618 12928 82634 12962
rect 82924 12928 82940 12962
rect 83116 12928 83132 12962
rect 83175 12956 83209 12972
rect 82270 12870 82300 12910
rect 82210 12810 82300 12870
rect 82210 12550 82230 12810
rect 82270 12758 82300 12810
rect 82290 12600 82300 12758
rect 83270 12910 83278 13068
rect 83270 12870 83300 12910
rect 83340 12870 83360 13110
rect 83270 12790 83360 12870
rect 83270 12758 83300 12790
rect 82358 12696 82392 12712
rect 82426 12706 82442 12740
rect 82618 12706 82634 12740
rect 82924 12706 82940 12740
rect 83116 12706 83132 12740
rect 82358 12646 82392 12662
rect 83175 12696 83209 12712
rect 82426 12618 82442 12652
rect 82618 12618 82634 12652
rect 82924 12618 82940 12652
rect 83116 12618 83132 12652
rect 83175 12646 83209 12662
rect 82270 12550 82300 12600
rect 82210 12430 82300 12550
rect 83270 12600 83278 12758
rect 83270 12550 83300 12600
rect 83340 12550 83360 12790
rect 83270 12430 83360 12550
rect -2080 11400 -1990 11530
rect -2080 11160 -2060 11400
rect -2020 11358 -1990 11400
rect -2000 11200 -1990 11358
rect -1020 11400 -930 11530
rect -1020 11358 -990 11400
rect -1932 11296 -1898 11312
rect -1864 11306 -1848 11340
rect -1672 11306 -1656 11340
rect -1366 11306 -1350 11340
rect -1174 11306 -1158 11340
rect -1932 11246 -1898 11262
rect -1115 11296 -1081 11312
rect -1864 11218 -1848 11252
rect -1672 11218 -1656 11252
rect -1366 11218 -1350 11252
rect -1174 11218 -1158 11252
rect -1115 11246 -1081 11262
rect -2020 11160 -1990 11200
rect -2080 11100 -1990 11160
rect -2080 10840 -2060 11100
rect -2020 11048 -1990 11100
rect -2000 10890 -1990 11048
rect -1020 11200 -1012 11358
rect -1020 11160 -990 11200
rect -950 11160 -930 11400
rect -1020 11080 -930 11160
rect -1020 11048 -990 11080
rect -1932 10986 -1898 11002
rect -1864 10996 -1848 11030
rect -1672 10996 -1656 11030
rect -1366 10996 -1350 11030
rect -1174 10996 -1158 11030
rect -1932 10936 -1898 10952
rect -1115 10986 -1081 11002
rect -1864 10908 -1848 10942
rect -1672 10908 -1656 10942
rect -1366 10908 -1350 10942
rect -1174 10908 -1158 10942
rect -1115 10936 -1081 10952
rect -2020 10840 -1990 10890
rect -2080 10720 -1990 10840
rect -1020 10890 -1012 11048
rect -1020 10840 -990 10890
rect -950 10840 -930 11080
rect -1020 10720 -930 10840
rect 82210 11400 82300 11530
rect 82210 11160 82230 11400
rect 82270 11358 82300 11400
rect 82290 11200 82300 11358
rect 83270 11400 83360 11530
rect 83270 11358 83300 11400
rect 82358 11296 82392 11312
rect 82426 11306 82442 11340
rect 82618 11306 82634 11340
rect 82924 11306 82940 11340
rect 83116 11306 83132 11340
rect 82358 11246 82392 11262
rect 83175 11296 83209 11312
rect 82426 11218 82442 11252
rect 82618 11218 82634 11252
rect 82924 11218 82940 11252
rect 83116 11218 83132 11252
rect 83175 11246 83209 11262
rect 82270 11160 82300 11200
rect 82210 11100 82300 11160
rect 82210 10840 82230 11100
rect 82270 11048 82300 11100
rect 82290 10890 82300 11048
rect 83270 11200 83278 11358
rect 83270 11160 83300 11200
rect 83340 11160 83360 11400
rect 83270 11080 83360 11160
rect 83270 11048 83300 11080
rect 82358 10986 82392 11002
rect 82426 10996 82442 11030
rect 82618 10996 82634 11030
rect 82924 10996 82940 11030
rect 83116 10996 83132 11030
rect 82358 10936 82392 10952
rect 83175 10986 83209 11002
rect 82426 10908 82442 10942
rect 82618 10908 82634 10942
rect 82924 10908 82940 10942
rect 83116 10908 83132 10942
rect 83175 10936 83209 10952
rect 82270 10840 82300 10890
rect 82210 10720 82300 10840
rect 83270 10890 83278 11048
rect 83270 10840 83300 10890
rect 83340 10840 83360 11080
rect 83270 10720 83360 10840
rect -2080 9690 -1990 9820
rect -2080 9450 -2060 9690
rect -2020 9648 -1990 9690
rect -2000 9490 -1990 9648
rect -1020 9690 -930 9820
rect -1020 9648 -990 9690
rect -1932 9586 -1898 9602
rect -1864 9596 -1848 9630
rect -1672 9596 -1656 9630
rect -1366 9596 -1350 9630
rect -1174 9596 -1158 9630
rect -1932 9536 -1898 9552
rect -1115 9586 -1081 9602
rect -1864 9508 -1848 9542
rect -1672 9508 -1656 9542
rect -1366 9508 -1350 9542
rect -1174 9508 -1158 9542
rect -1115 9536 -1081 9552
rect -2020 9450 -1990 9490
rect -2080 9390 -1990 9450
rect -2080 9130 -2060 9390
rect -2020 9338 -1990 9390
rect -2000 9180 -1990 9338
rect -1020 9490 -1012 9648
rect -1020 9450 -990 9490
rect -950 9450 -930 9690
rect -1020 9370 -930 9450
rect -1020 9338 -990 9370
rect -1932 9276 -1898 9292
rect -1864 9286 -1848 9320
rect -1672 9286 -1656 9320
rect -1366 9286 -1350 9320
rect -1174 9286 -1158 9320
rect -1932 9226 -1898 9242
rect -1115 9276 -1081 9292
rect -1864 9198 -1848 9232
rect -1672 9198 -1656 9232
rect -1366 9198 -1350 9232
rect -1174 9198 -1158 9232
rect -1115 9226 -1081 9242
rect -2020 9130 -1990 9180
rect -2080 9010 -1990 9130
rect -1020 9180 -1012 9338
rect -1020 9130 -990 9180
rect -950 9130 -930 9370
rect -1020 9010 -930 9130
rect 82210 9690 82300 9820
rect 82210 9450 82230 9690
rect 82270 9648 82300 9690
rect 82290 9490 82300 9648
rect 83270 9690 83360 9820
rect 83270 9648 83300 9690
rect 82358 9586 82392 9602
rect 82426 9596 82442 9630
rect 82618 9596 82634 9630
rect 82924 9596 82940 9630
rect 83116 9596 83132 9630
rect 82358 9536 82392 9552
rect 83175 9586 83209 9602
rect 82426 9508 82442 9542
rect 82618 9508 82634 9542
rect 82924 9508 82940 9542
rect 83116 9508 83132 9542
rect 83175 9536 83209 9552
rect 82270 9450 82300 9490
rect 82210 9390 82300 9450
rect 82210 9130 82230 9390
rect 82270 9338 82300 9390
rect 82290 9180 82300 9338
rect 83270 9490 83278 9648
rect 83270 9450 83300 9490
rect 83340 9450 83360 9690
rect 83270 9370 83360 9450
rect 83270 9338 83300 9370
rect 82358 9276 82392 9292
rect 82426 9286 82442 9320
rect 82618 9286 82634 9320
rect 82924 9286 82940 9320
rect 83116 9286 83132 9320
rect 82358 9226 82392 9242
rect 83175 9276 83209 9292
rect 82426 9198 82442 9232
rect 82618 9198 82634 9232
rect 82924 9198 82940 9232
rect 83116 9198 83132 9232
rect 83175 9226 83209 9242
rect 82270 9130 82300 9180
rect 82210 9010 82300 9130
rect 83270 9180 83278 9338
rect 83270 9130 83300 9180
rect 83340 9130 83360 9370
rect 83270 9010 83360 9130
rect -2080 7980 -1990 8110
rect -2080 7740 -2060 7980
rect -2020 7938 -1990 7980
rect -2000 7780 -1990 7938
rect -1020 7980 -930 8110
rect -1020 7938 -990 7980
rect -1932 7876 -1898 7892
rect -1864 7886 -1848 7920
rect -1672 7886 -1656 7920
rect -1366 7886 -1350 7920
rect -1174 7886 -1158 7920
rect -1932 7826 -1898 7842
rect -1115 7876 -1081 7892
rect -1864 7798 -1848 7832
rect -1672 7798 -1656 7832
rect -1366 7798 -1350 7832
rect -1174 7798 -1158 7832
rect -1115 7826 -1081 7842
rect -2020 7740 -1990 7780
rect -2080 7680 -1990 7740
rect -2080 7420 -2060 7680
rect -2020 7628 -1990 7680
rect -2000 7470 -1990 7628
rect -1020 7780 -1012 7938
rect -1020 7740 -990 7780
rect -950 7740 -930 7980
rect -1020 7660 -930 7740
rect -1020 7628 -990 7660
rect -1932 7566 -1898 7582
rect -1864 7576 -1848 7610
rect -1672 7576 -1656 7610
rect -1366 7576 -1350 7610
rect -1174 7576 -1158 7610
rect -1932 7516 -1898 7532
rect -1115 7566 -1081 7582
rect -1864 7488 -1848 7522
rect -1672 7488 -1656 7522
rect -1366 7488 -1350 7522
rect -1174 7488 -1158 7522
rect -1115 7516 -1081 7532
rect -2020 7420 -1990 7470
rect -2080 7300 -1990 7420
rect -1020 7470 -1012 7628
rect -1020 7420 -990 7470
rect -950 7420 -930 7660
rect -1020 7300 -930 7420
rect 82210 7980 82300 8110
rect 82210 7740 82230 7980
rect 82270 7938 82300 7980
rect 82290 7780 82300 7938
rect 83270 7980 83360 8110
rect 83270 7938 83300 7980
rect 82358 7876 82392 7892
rect 82426 7886 82442 7920
rect 82618 7886 82634 7920
rect 82924 7886 82940 7920
rect 83116 7886 83132 7920
rect 82358 7826 82392 7842
rect 83175 7876 83209 7892
rect 82426 7798 82442 7832
rect 82618 7798 82634 7832
rect 82924 7798 82940 7832
rect 83116 7798 83132 7832
rect 83175 7826 83209 7842
rect 82270 7740 82300 7780
rect 82210 7680 82300 7740
rect 82210 7420 82230 7680
rect 82270 7628 82300 7680
rect 82290 7470 82300 7628
rect 83270 7780 83278 7938
rect 83270 7740 83300 7780
rect 83340 7740 83360 7980
rect 83270 7660 83360 7740
rect 83270 7628 83300 7660
rect 82358 7566 82392 7582
rect 82426 7576 82442 7610
rect 82618 7576 82634 7610
rect 82924 7576 82940 7610
rect 83116 7576 83132 7610
rect 82358 7516 82392 7532
rect 83175 7566 83209 7582
rect 82426 7488 82442 7522
rect 82618 7488 82634 7522
rect 82924 7488 82940 7522
rect 83116 7488 83132 7522
rect 83175 7516 83209 7532
rect 82270 7420 82300 7470
rect 82210 7300 82300 7420
rect 83270 7470 83278 7628
rect 83270 7420 83300 7470
rect 83340 7420 83360 7660
rect 83270 7300 83360 7420
rect -2080 6270 -1990 6400
rect -2080 6030 -2060 6270
rect -2020 6228 -1990 6270
rect -2000 6070 -1990 6228
rect -1020 6270 -930 6400
rect -1020 6228 -990 6270
rect -1932 6166 -1898 6182
rect -1864 6176 -1848 6210
rect -1672 6176 -1656 6210
rect -1366 6176 -1350 6210
rect -1174 6176 -1158 6210
rect -1932 6116 -1898 6132
rect -1115 6166 -1081 6182
rect -1864 6088 -1848 6122
rect -1672 6088 -1656 6122
rect -1366 6088 -1350 6122
rect -1174 6088 -1158 6122
rect -1115 6116 -1081 6132
rect -2020 6030 -1990 6070
rect -2080 5970 -1990 6030
rect -2080 5710 -2060 5970
rect -2020 5918 -1990 5970
rect -2000 5760 -1990 5918
rect -1020 6070 -1012 6228
rect -1020 6030 -990 6070
rect -950 6030 -930 6270
rect -1020 5950 -930 6030
rect -1020 5918 -990 5950
rect -1932 5856 -1898 5872
rect -1864 5866 -1848 5900
rect -1672 5866 -1656 5900
rect -1366 5866 -1350 5900
rect -1174 5866 -1158 5900
rect -1932 5806 -1898 5822
rect -1115 5856 -1081 5872
rect -1864 5778 -1848 5812
rect -1672 5778 -1656 5812
rect -1366 5778 -1350 5812
rect -1174 5778 -1158 5812
rect -1115 5806 -1081 5822
rect -2020 5710 -1990 5760
rect -2080 5590 -1990 5710
rect -1020 5760 -1012 5918
rect -1020 5710 -990 5760
rect -950 5710 -930 5950
rect -1020 5590 -930 5710
rect 82210 6270 82300 6400
rect 82210 6030 82230 6270
rect 82270 6228 82300 6270
rect 82290 6070 82300 6228
rect 83270 6270 83360 6400
rect 83270 6228 83300 6270
rect 82358 6166 82392 6182
rect 82426 6176 82442 6210
rect 82618 6176 82634 6210
rect 82924 6176 82940 6210
rect 83116 6176 83132 6210
rect 82358 6116 82392 6132
rect 83175 6166 83209 6182
rect 82426 6088 82442 6122
rect 82618 6088 82634 6122
rect 82924 6088 82940 6122
rect 83116 6088 83132 6122
rect 83175 6116 83209 6132
rect 82270 6030 82300 6070
rect 82210 5970 82300 6030
rect 82210 5710 82230 5970
rect 82270 5918 82300 5970
rect 82290 5760 82300 5918
rect 83270 6070 83278 6228
rect 83270 6030 83300 6070
rect 83340 6030 83360 6270
rect 83270 5950 83360 6030
rect 83270 5918 83300 5950
rect 82358 5856 82392 5872
rect 82426 5866 82442 5900
rect 82618 5866 82634 5900
rect 82924 5866 82940 5900
rect 83116 5866 83132 5900
rect 82358 5806 82392 5822
rect 83175 5856 83209 5872
rect 82426 5778 82442 5812
rect 82618 5778 82634 5812
rect 82924 5778 82940 5812
rect 83116 5778 83132 5812
rect 83175 5806 83209 5822
rect 82270 5710 82300 5760
rect 82210 5590 82300 5710
rect 83270 5760 83278 5918
rect 83270 5710 83300 5760
rect 83340 5710 83360 5950
rect 83270 5590 83360 5710
rect -2080 4560 -1990 4690
rect -2080 4320 -2060 4560
rect -2020 4518 -1990 4560
rect -2000 4360 -1990 4518
rect -1020 4560 -930 4690
rect -1020 4518 -990 4560
rect -1932 4456 -1898 4472
rect -1864 4466 -1848 4500
rect -1672 4466 -1656 4500
rect -1366 4466 -1350 4500
rect -1174 4466 -1158 4500
rect -1932 4406 -1898 4422
rect -1115 4456 -1081 4472
rect -1864 4378 -1848 4412
rect -1672 4378 -1656 4412
rect -1366 4378 -1350 4412
rect -1174 4378 -1158 4412
rect -1115 4406 -1081 4422
rect -2020 4320 -1990 4360
rect -2080 4260 -1990 4320
rect -2080 4000 -2060 4260
rect -2020 4208 -1990 4260
rect -2000 4050 -1990 4208
rect -1020 4360 -1012 4518
rect -1020 4320 -990 4360
rect -950 4320 -930 4560
rect -1020 4240 -930 4320
rect -1020 4208 -990 4240
rect -1932 4146 -1898 4162
rect -1864 4156 -1848 4190
rect -1672 4156 -1656 4190
rect -1366 4156 -1350 4190
rect -1174 4156 -1158 4190
rect -1932 4096 -1898 4112
rect -1115 4146 -1081 4162
rect -1864 4068 -1848 4102
rect -1672 4068 -1656 4102
rect -1366 4068 -1350 4102
rect -1174 4068 -1158 4102
rect -1115 4096 -1081 4112
rect -2020 4000 -1990 4050
rect -2080 3880 -1990 4000
rect -1020 4050 -1012 4208
rect -1020 4000 -990 4050
rect -950 4000 -930 4240
rect -1020 3880 -930 4000
rect 82210 4560 82300 4690
rect 82210 4320 82230 4560
rect 82270 4518 82300 4560
rect 82290 4360 82300 4518
rect 83270 4560 83360 4690
rect 83270 4518 83300 4560
rect 82358 4456 82392 4472
rect 82426 4466 82442 4500
rect 82618 4466 82634 4500
rect 82924 4466 82940 4500
rect 83116 4466 83132 4500
rect 82358 4406 82392 4422
rect 83175 4456 83209 4472
rect 82426 4378 82442 4412
rect 82618 4378 82634 4412
rect 82924 4378 82940 4412
rect 83116 4378 83132 4412
rect 83175 4406 83209 4422
rect 82270 4320 82300 4360
rect 82210 4260 82300 4320
rect 82210 4000 82230 4260
rect 82270 4208 82300 4260
rect 82290 4050 82300 4208
rect 83270 4360 83278 4518
rect 83270 4320 83300 4360
rect 83340 4320 83360 4560
rect 83270 4240 83360 4320
rect 83270 4208 83300 4240
rect 82358 4146 82392 4162
rect 82426 4156 82442 4190
rect 82618 4156 82634 4190
rect 82924 4156 82940 4190
rect 83116 4156 83132 4190
rect 82358 4096 82392 4112
rect 83175 4146 83209 4162
rect 82426 4068 82442 4102
rect 82618 4068 82634 4102
rect 82924 4068 82940 4102
rect 83116 4068 83132 4102
rect 83175 4096 83209 4112
rect 82270 4000 82300 4050
rect 82210 3880 82300 4000
rect 83270 4050 83278 4208
rect 83270 4000 83300 4050
rect 83340 4000 83360 4240
rect 83270 3880 83360 4000
rect -2080 2850 -1990 2980
rect -2080 2610 -2060 2850
rect -2020 2808 -1990 2850
rect -2000 2650 -1990 2808
rect -1020 2850 -930 2980
rect -1020 2808 -990 2850
rect -1932 2746 -1898 2762
rect -1864 2756 -1848 2790
rect -1672 2756 -1656 2790
rect -1366 2756 -1350 2790
rect -1174 2756 -1158 2790
rect -1932 2696 -1898 2712
rect -1115 2746 -1081 2762
rect -1864 2668 -1848 2702
rect -1672 2668 -1656 2702
rect -1366 2668 -1350 2702
rect -1174 2668 -1158 2702
rect -1115 2696 -1081 2712
rect -2020 2610 -1990 2650
rect -2080 2550 -1990 2610
rect -2080 2290 -2060 2550
rect -2020 2498 -1990 2550
rect -2000 2340 -1990 2498
rect -1020 2650 -1012 2808
rect -1020 2610 -990 2650
rect -950 2610 -930 2850
rect -1020 2530 -930 2610
rect -1020 2498 -990 2530
rect -1932 2436 -1898 2452
rect -1864 2446 -1848 2480
rect -1672 2446 -1656 2480
rect -1366 2446 -1350 2480
rect -1174 2446 -1158 2480
rect -1932 2386 -1898 2402
rect -1115 2436 -1081 2452
rect -1864 2358 -1848 2392
rect -1672 2358 -1656 2392
rect -1366 2358 -1350 2392
rect -1174 2358 -1158 2392
rect -1115 2386 -1081 2402
rect -2020 2290 -1990 2340
rect -2080 2170 -1990 2290
rect -1020 2340 -1012 2498
rect -1020 2290 -990 2340
rect -950 2290 -930 2530
rect -1020 2170 -930 2290
rect 82210 2850 82300 2980
rect 82210 2610 82230 2850
rect 82270 2808 82300 2850
rect 82290 2650 82300 2808
rect 83270 2850 83360 2980
rect 83270 2808 83300 2850
rect 82358 2746 82392 2762
rect 82426 2756 82442 2790
rect 82618 2756 82634 2790
rect 82924 2756 82940 2790
rect 83116 2756 83132 2790
rect 82358 2696 82392 2712
rect 83175 2746 83209 2762
rect 82426 2668 82442 2702
rect 82618 2668 82634 2702
rect 82924 2668 82940 2702
rect 83116 2668 83132 2702
rect 83175 2696 83209 2712
rect 82270 2610 82300 2650
rect 82210 2550 82300 2610
rect 82210 2290 82230 2550
rect 82270 2498 82300 2550
rect 82290 2340 82300 2498
rect 83270 2650 83278 2808
rect 83270 2610 83300 2650
rect 83340 2610 83360 2850
rect 83270 2530 83360 2610
rect 83270 2498 83300 2530
rect 82358 2436 82392 2452
rect 82426 2446 82442 2480
rect 82618 2446 82634 2480
rect 82924 2446 82940 2480
rect 83116 2446 83132 2480
rect 82358 2386 82392 2402
rect 83175 2436 83209 2452
rect 82426 2358 82442 2392
rect 82618 2358 82634 2392
rect 82924 2358 82940 2392
rect 83116 2358 83132 2392
rect 83175 2386 83209 2402
rect 82270 2290 82300 2340
rect 82210 2170 82300 2290
rect 83270 2340 83278 2498
rect 83270 2290 83300 2340
rect 83340 2290 83360 2530
rect 83270 2170 83360 2290
rect -2080 1140 -1990 1270
rect -2080 900 -2060 1140
rect -2020 1098 -1990 1140
rect -2000 940 -1990 1098
rect -1020 1140 -930 1270
rect -1020 1098 -990 1140
rect -1932 1036 -1898 1052
rect -1864 1046 -1848 1080
rect -1672 1046 -1656 1080
rect -1366 1046 -1350 1080
rect -1174 1046 -1158 1080
rect -1932 986 -1898 1002
rect -1115 1036 -1081 1052
rect -1864 958 -1848 992
rect -1672 958 -1656 992
rect -1366 958 -1350 992
rect -1174 958 -1158 992
rect -1115 986 -1081 1002
rect -2020 900 -1990 940
rect -2080 840 -1990 900
rect -2080 580 -2060 840
rect -2020 788 -1990 840
rect -2000 630 -1990 788
rect -1020 940 -1012 1098
rect -1020 900 -990 940
rect -950 900 -930 1140
rect -1020 820 -930 900
rect -1020 788 -990 820
rect -1932 726 -1898 742
rect -1864 736 -1848 770
rect -1672 736 -1656 770
rect -1366 736 -1350 770
rect -1174 736 -1158 770
rect -1932 676 -1898 692
rect -1115 726 -1081 742
rect -1864 648 -1848 682
rect -1672 648 -1656 682
rect -1366 648 -1350 682
rect -1174 648 -1158 682
rect -1115 676 -1081 692
rect -2020 580 -1990 630
rect -2080 460 -1990 580
rect -1020 630 -1012 788
rect -1020 580 -990 630
rect -950 580 -930 820
rect -1020 460 -930 580
rect 82210 1140 82300 1270
rect 82210 900 82230 1140
rect 82270 1098 82300 1140
rect 82290 940 82300 1098
rect 83270 1140 83360 1270
rect 83270 1098 83300 1140
rect 82358 1036 82392 1052
rect 82426 1046 82442 1080
rect 82618 1046 82634 1080
rect 82924 1046 82940 1080
rect 83116 1046 83132 1080
rect 82358 986 82392 1002
rect 83175 1036 83209 1052
rect 82426 958 82442 992
rect 82618 958 82634 992
rect 82924 958 82940 992
rect 83116 958 83132 992
rect 83175 986 83209 1002
rect 82270 900 82300 940
rect 82210 840 82300 900
rect 82210 580 82230 840
rect 82270 788 82300 840
rect 82290 630 82300 788
rect 83270 940 83278 1098
rect 83270 900 83300 940
rect 83340 900 83360 1140
rect 83270 820 83360 900
rect 83270 788 83300 820
rect 82358 726 82392 742
rect 82426 736 82442 770
rect 82618 736 82634 770
rect 82924 736 82940 770
rect 83116 736 83132 770
rect 82358 676 82392 692
rect 83175 726 83209 742
rect 82426 648 82442 682
rect 82618 648 82634 682
rect 82924 648 82940 682
rect 83116 648 83132 682
rect 83175 676 83209 692
rect 82270 580 82300 630
rect 82210 460 82300 580
rect 83270 630 83278 788
rect 83270 580 83300 630
rect 83340 580 83360 820
rect 83270 460 83360 580
rect -2080 -570 -1990 -440
rect -2080 -810 -2060 -570
rect -2020 -612 -1990 -570
rect -2000 -770 -1990 -612
rect -1020 -570 -930 -440
rect -1020 -612 -990 -570
rect -1932 -674 -1898 -658
rect -1864 -664 -1848 -630
rect -1672 -664 -1656 -630
rect -1366 -664 -1350 -630
rect -1174 -664 -1158 -630
rect -1932 -724 -1898 -708
rect -1115 -674 -1081 -658
rect -1864 -752 -1848 -718
rect -1672 -752 -1656 -718
rect -1366 -752 -1350 -718
rect -1174 -752 -1158 -718
rect -1115 -724 -1081 -708
rect -2020 -810 -1990 -770
rect -2080 -870 -1990 -810
rect -2080 -1130 -2060 -870
rect -2020 -922 -1990 -870
rect -2000 -1080 -1990 -922
rect -1020 -770 -1012 -612
rect -1020 -810 -990 -770
rect -950 -810 -930 -570
rect -1020 -890 -930 -810
rect -1020 -922 -990 -890
rect -1932 -984 -1898 -968
rect -1864 -974 -1848 -940
rect -1672 -974 -1656 -940
rect -1366 -974 -1350 -940
rect -1174 -974 -1158 -940
rect -1932 -1034 -1898 -1018
rect -1115 -984 -1081 -968
rect -1864 -1062 -1848 -1028
rect -1672 -1062 -1656 -1028
rect -1366 -1062 -1350 -1028
rect -1174 -1062 -1158 -1028
rect -1115 -1034 -1081 -1018
rect -2020 -1130 -1990 -1080
rect -2080 -1250 -1990 -1130
rect -1020 -1080 -1012 -922
rect -1020 -1130 -990 -1080
rect -950 -1130 -930 -890
rect -1020 -1250 -930 -1130
rect 2640 -570 2730 -440
rect 2640 -810 2660 -570
rect 2700 -612 2730 -570
rect 2720 -770 2730 -612
rect 3700 -570 3790 -440
rect 3700 -612 3730 -570
rect 2788 -674 2822 -658
rect 2856 -664 2872 -630
rect 3048 -664 3064 -630
rect 3354 -664 3370 -630
rect 3546 -664 3562 -630
rect 2788 -724 2822 -708
rect 3605 -674 3639 -658
rect 2856 -752 2872 -718
rect 3048 -752 3064 -718
rect 3354 -752 3370 -718
rect 3546 -752 3562 -718
rect 3605 -724 3639 -708
rect 2700 -810 2730 -770
rect 2640 -870 2730 -810
rect 2640 -1130 2660 -870
rect 2700 -922 2730 -870
rect 2720 -1080 2730 -922
rect 3700 -770 3708 -612
rect 3700 -810 3730 -770
rect 3770 -810 3790 -570
rect 3700 -890 3790 -810
rect 3700 -922 3730 -890
rect 2788 -984 2822 -968
rect 2856 -974 2872 -940
rect 3048 -974 3064 -940
rect 3354 -974 3370 -940
rect 3546 -974 3562 -940
rect 2788 -1034 2822 -1018
rect 3605 -984 3639 -968
rect 2856 -1062 2872 -1028
rect 3048 -1062 3064 -1028
rect 3354 -1062 3370 -1028
rect 3546 -1062 3562 -1028
rect 3605 -1034 3639 -1018
rect 2700 -1130 2730 -1080
rect 2640 -1250 2730 -1130
rect 3700 -1080 3708 -922
rect 3700 -1130 3730 -1080
rect 3770 -1130 3790 -890
rect 3700 -1250 3790 -1130
rect 7630 -570 7720 -440
rect 7630 -810 7650 -570
rect 7690 -612 7720 -570
rect 7710 -770 7720 -612
rect 8690 -570 8780 -440
rect 8690 -612 8720 -570
rect 7778 -674 7812 -658
rect 7846 -664 7862 -630
rect 8038 -664 8054 -630
rect 8344 -664 8360 -630
rect 8536 -664 8552 -630
rect 7778 -724 7812 -708
rect 8595 -674 8629 -658
rect 7846 -752 7862 -718
rect 8038 -752 8054 -718
rect 8344 -752 8360 -718
rect 8536 -752 8552 -718
rect 8595 -724 8629 -708
rect 7690 -810 7720 -770
rect 7630 -870 7720 -810
rect 7630 -1130 7650 -870
rect 7690 -922 7720 -870
rect 7710 -1080 7720 -922
rect 8690 -770 8698 -612
rect 8690 -810 8720 -770
rect 8760 -810 8780 -570
rect 8690 -890 8780 -810
rect 8690 -922 8720 -890
rect 7778 -984 7812 -968
rect 7846 -974 7862 -940
rect 8038 -974 8054 -940
rect 8344 -974 8360 -940
rect 8536 -974 8552 -940
rect 7778 -1034 7812 -1018
rect 8595 -984 8629 -968
rect 7846 -1062 7862 -1028
rect 8038 -1062 8054 -1028
rect 8344 -1062 8360 -1028
rect 8536 -1062 8552 -1028
rect 8595 -1034 8629 -1018
rect 7690 -1130 7720 -1080
rect 7630 -1250 7720 -1130
rect 8690 -1080 8698 -922
rect 8690 -1130 8720 -1080
rect 8760 -1130 8780 -890
rect 8690 -1250 8780 -1130
rect 12620 -570 12710 -440
rect 12620 -810 12640 -570
rect 12680 -612 12710 -570
rect 12700 -770 12710 -612
rect 13680 -570 13770 -440
rect 13680 -612 13710 -570
rect 12768 -674 12802 -658
rect 12836 -664 12852 -630
rect 13028 -664 13044 -630
rect 13334 -664 13350 -630
rect 13526 -664 13542 -630
rect 12768 -724 12802 -708
rect 13585 -674 13619 -658
rect 12836 -752 12852 -718
rect 13028 -752 13044 -718
rect 13334 -752 13350 -718
rect 13526 -752 13542 -718
rect 13585 -724 13619 -708
rect 12680 -810 12710 -770
rect 12620 -870 12710 -810
rect 12620 -1130 12640 -870
rect 12680 -922 12710 -870
rect 12700 -1080 12710 -922
rect 13680 -770 13688 -612
rect 13680 -810 13710 -770
rect 13750 -810 13770 -570
rect 13680 -890 13770 -810
rect 13680 -922 13710 -890
rect 12768 -984 12802 -968
rect 12836 -974 12852 -940
rect 13028 -974 13044 -940
rect 13334 -974 13350 -940
rect 13526 -974 13542 -940
rect 12768 -1034 12802 -1018
rect 13585 -984 13619 -968
rect 12836 -1062 12852 -1028
rect 13028 -1062 13044 -1028
rect 13334 -1062 13350 -1028
rect 13526 -1062 13542 -1028
rect 13585 -1034 13619 -1018
rect 12680 -1130 12710 -1080
rect 12620 -1250 12710 -1130
rect 13680 -1080 13688 -922
rect 13680 -1130 13710 -1080
rect 13750 -1130 13770 -890
rect 13680 -1250 13770 -1130
rect 17610 -570 17700 -440
rect 17610 -810 17630 -570
rect 17670 -612 17700 -570
rect 17690 -770 17700 -612
rect 18670 -570 18760 -440
rect 18670 -612 18700 -570
rect 17758 -674 17792 -658
rect 17826 -664 17842 -630
rect 18018 -664 18034 -630
rect 18324 -664 18340 -630
rect 18516 -664 18532 -630
rect 17758 -724 17792 -708
rect 18575 -674 18609 -658
rect 17826 -752 17842 -718
rect 18018 -752 18034 -718
rect 18324 -752 18340 -718
rect 18516 -752 18532 -718
rect 18575 -724 18609 -708
rect 17670 -810 17700 -770
rect 17610 -870 17700 -810
rect 17610 -1130 17630 -870
rect 17670 -922 17700 -870
rect 17690 -1080 17700 -922
rect 18670 -770 18678 -612
rect 18670 -810 18700 -770
rect 18740 -810 18760 -570
rect 18670 -890 18760 -810
rect 18670 -922 18700 -890
rect 17758 -984 17792 -968
rect 17826 -974 17842 -940
rect 18018 -974 18034 -940
rect 18324 -974 18340 -940
rect 18516 -974 18532 -940
rect 17758 -1034 17792 -1018
rect 18575 -984 18609 -968
rect 17826 -1062 17842 -1028
rect 18018 -1062 18034 -1028
rect 18324 -1062 18340 -1028
rect 18516 -1062 18532 -1028
rect 18575 -1034 18609 -1018
rect 17670 -1130 17700 -1080
rect 17610 -1250 17700 -1130
rect 18670 -1080 18678 -922
rect 18670 -1130 18700 -1080
rect 18740 -1130 18760 -890
rect 18670 -1250 18760 -1130
rect 22600 -570 22690 -440
rect 22600 -810 22620 -570
rect 22660 -612 22690 -570
rect 22680 -770 22690 -612
rect 23660 -570 23750 -440
rect 23660 -612 23690 -570
rect 22748 -674 22782 -658
rect 22816 -664 22832 -630
rect 23008 -664 23024 -630
rect 23314 -664 23330 -630
rect 23506 -664 23522 -630
rect 22748 -724 22782 -708
rect 23565 -674 23599 -658
rect 22816 -752 22832 -718
rect 23008 -752 23024 -718
rect 23314 -752 23330 -718
rect 23506 -752 23522 -718
rect 23565 -724 23599 -708
rect 22660 -810 22690 -770
rect 22600 -870 22690 -810
rect 22600 -1130 22620 -870
rect 22660 -922 22690 -870
rect 22680 -1080 22690 -922
rect 23660 -770 23668 -612
rect 23660 -810 23690 -770
rect 23730 -810 23750 -570
rect 23660 -890 23750 -810
rect 23660 -922 23690 -890
rect 22748 -984 22782 -968
rect 22816 -974 22832 -940
rect 23008 -974 23024 -940
rect 23314 -974 23330 -940
rect 23506 -974 23522 -940
rect 22748 -1034 22782 -1018
rect 23565 -984 23599 -968
rect 22816 -1062 22832 -1028
rect 23008 -1062 23024 -1028
rect 23314 -1062 23330 -1028
rect 23506 -1062 23522 -1028
rect 23565 -1034 23599 -1018
rect 22660 -1130 22690 -1080
rect 22600 -1250 22690 -1130
rect 23660 -1080 23668 -922
rect 23660 -1130 23690 -1080
rect 23730 -1130 23750 -890
rect 23660 -1250 23750 -1130
rect 27590 -570 27680 -440
rect 27590 -810 27610 -570
rect 27650 -612 27680 -570
rect 27670 -770 27680 -612
rect 28650 -570 28740 -440
rect 28650 -612 28680 -570
rect 27738 -674 27772 -658
rect 27806 -664 27822 -630
rect 27998 -664 28014 -630
rect 28304 -664 28320 -630
rect 28496 -664 28512 -630
rect 27738 -724 27772 -708
rect 28555 -674 28589 -658
rect 27806 -752 27822 -718
rect 27998 -752 28014 -718
rect 28304 -752 28320 -718
rect 28496 -752 28512 -718
rect 28555 -724 28589 -708
rect 27650 -810 27680 -770
rect 27590 -870 27680 -810
rect 27590 -1130 27610 -870
rect 27650 -922 27680 -870
rect 27670 -1080 27680 -922
rect 28650 -770 28658 -612
rect 28650 -810 28680 -770
rect 28720 -810 28740 -570
rect 28650 -890 28740 -810
rect 28650 -922 28680 -890
rect 27738 -984 27772 -968
rect 27806 -974 27822 -940
rect 27998 -974 28014 -940
rect 28304 -974 28320 -940
rect 28496 -974 28512 -940
rect 27738 -1034 27772 -1018
rect 28555 -984 28589 -968
rect 27806 -1062 27822 -1028
rect 27998 -1062 28014 -1028
rect 28304 -1062 28320 -1028
rect 28496 -1062 28512 -1028
rect 28555 -1034 28589 -1018
rect 27650 -1130 27680 -1080
rect 27590 -1250 27680 -1130
rect 28650 -1080 28658 -922
rect 28650 -1130 28680 -1080
rect 28720 -1130 28740 -890
rect 28650 -1250 28740 -1130
rect 32580 -570 32670 -440
rect 32580 -810 32600 -570
rect 32640 -612 32670 -570
rect 32660 -770 32670 -612
rect 33640 -570 33730 -440
rect 33640 -612 33670 -570
rect 32728 -674 32762 -658
rect 32796 -664 32812 -630
rect 32988 -664 33004 -630
rect 33294 -664 33310 -630
rect 33486 -664 33502 -630
rect 32728 -724 32762 -708
rect 33545 -674 33579 -658
rect 32796 -752 32812 -718
rect 32988 -752 33004 -718
rect 33294 -752 33310 -718
rect 33486 -752 33502 -718
rect 33545 -724 33579 -708
rect 32640 -810 32670 -770
rect 32580 -870 32670 -810
rect 32580 -1130 32600 -870
rect 32640 -922 32670 -870
rect 32660 -1080 32670 -922
rect 33640 -770 33648 -612
rect 33640 -810 33670 -770
rect 33710 -810 33730 -570
rect 33640 -890 33730 -810
rect 33640 -922 33670 -890
rect 32728 -984 32762 -968
rect 32796 -974 32812 -940
rect 32988 -974 33004 -940
rect 33294 -974 33310 -940
rect 33486 -974 33502 -940
rect 32728 -1034 32762 -1018
rect 33545 -984 33579 -968
rect 32796 -1062 32812 -1028
rect 32988 -1062 33004 -1028
rect 33294 -1062 33310 -1028
rect 33486 -1062 33502 -1028
rect 33545 -1034 33579 -1018
rect 32640 -1130 32670 -1080
rect 32580 -1250 32670 -1130
rect 33640 -1080 33648 -922
rect 33640 -1130 33670 -1080
rect 33710 -1130 33730 -890
rect 33640 -1250 33730 -1130
rect 37570 -570 37660 -440
rect 37570 -810 37590 -570
rect 37630 -612 37660 -570
rect 37650 -770 37660 -612
rect 38630 -570 38720 -440
rect 38630 -612 38660 -570
rect 37718 -674 37752 -658
rect 37786 -664 37802 -630
rect 37978 -664 37994 -630
rect 38284 -664 38300 -630
rect 38476 -664 38492 -630
rect 37718 -724 37752 -708
rect 38535 -674 38569 -658
rect 37786 -752 37802 -718
rect 37978 -752 37994 -718
rect 38284 -752 38300 -718
rect 38476 -752 38492 -718
rect 38535 -724 38569 -708
rect 37630 -810 37660 -770
rect 37570 -870 37660 -810
rect 37570 -1130 37590 -870
rect 37630 -922 37660 -870
rect 37650 -1080 37660 -922
rect 38630 -770 38638 -612
rect 38630 -810 38660 -770
rect 38700 -810 38720 -570
rect 38630 -890 38720 -810
rect 38630 -922 38660 -890
rect 37718 -984 37752 -968
rect 37786 -974 37802 -940
rect 37978 -974 37994 -940
rect 38284 -974 38300 -940
rect 38476 -974 38492 -940
rect 37718 -1034 37752 -1018
rect 38535 -984 38569 -968
rect 37786 -1062 37802 -1028
rect 37978 -1062 37994 -1028
rect 38284 -1062 38300 -1028
rect 38476 -1062 38492 -1028
rect 38535 -1034 38569 -1018
rect 37630 -1130 37660 -1080
rect 37570 -1250 37660 -1130
rect 38630 -1080 38638 -922
rect 38630 -1130 38660 -1080
rect 38700 -1130 38720 -890
rect 38630 -1250 38720 -1130
rect 42560 -570 42650 -440
rect 42560 -810 42580 -570
rect 42620 -612 42650 -570
rect 42640 -770 42650 -612
rect 43620 -570 43710 -440
rect 43620 -612 43650 -570
rect 42708 -674 42742 -658
rect 42776 -664 42792 -630
rect 42968 -664 42984 -630
rect 43274 -664 43290 -630
rect 43466 -664 43482 -630
rect 42708 -724 42742 -708
rect 43525 -674 43559 -658
rect 42776 -752 42792 -718
rect 42968 -752 42984 -718
rect 43274 -752 43290 -718
rect 43466 -752 43482 -718
rect 43525 -724 43559 -708
rect 42620 -810 42650 -770
rect 42560 -870 42650 -810
rect 42560 -1130 42580 -870
rect 42620 -922 42650 -870
rect 42640 -1080 42650 -922
rect 43620 -770 43628 -612
rect 43620 -810 43650 -770
rect 43690 -810 43710 -570
rect 43620 -890 43710 -810
rect 43620 -922 43650 -890
rect 42708 -984 42742 -968
rect 42776 -974 42792 -940
rect 42968 -974 42984 -940
rect 43274 -974 43290 -940
rect 43466 -974 43482 -940
rect 42708 -1034 42742 -1018
rect 43525 -984 43559 -968
rect 42776 -1062 42792 -1028
rect 42968 -1062 42984 -1028
rect 43274 -1062 43290 -1028
rect 43466 -1062 43482 -1028
rect 43525 -1034 43559 -1018
rect 42620 -1130 42650 -1080
rect 42560 -1250 42650 -1130
rect 43620 -1080 43628 -922
rect 43620 -1130 43650 -1080
rect 43690 -1130 43710 -890
rect 43620 -1250 43710 -1130
rect 47550 -570 47640 -440
rect 47550 -810 47570 -570
rect 47610 -612 47640 -570
rect 47630 -770 47640 -612
rect 48610 -570 48700 -440
rect 48610 -612 48640 -570
rect 47698 -674 47732 -658
rect 47766 -664 47782 -630
rect 47958 -664 47974 -630
rect 48264 -664 48280 -630
rect 48456 -664 48472 -630
rect 47698 -724 47732 -708
rect 48515 -674 48549 -658
rect 47766 -752 47782 -718
rect 47958 -752 47974 -718
rect 48264 -752 48280 -718
rect 48456 -752 48472 -718
rect 48515 -724 48549 -708
rect 47610 -810 47640 -770
rect 47550 -870 47640 -810
rect 47550 -1130 47570 -870
rect 47610 -922 47640 -870
rect 47630 -1080 47640 -922
rect 48610 -770 48618 -612
rect 48610 -810 48640 -770
rect 48680 -810 48700 -570
rect 48610 -890 48700 -810
rect 48610 -922 48640 -890
rect 47698 -984 47732 -968
rect 47766 -974 47782 -940
rect 47958 -974 47974 -940
rect 48264 -974 48280 -940
rect 48456 -974 48472 -940
rect 47698 -1034 47732 -1018
rect 48515 -984 48549 -968
rect 47766 -1062 47782 -1028
rect 47958 -1062 47974 -1028
rect 48264 -1062 48280 -1028
rect 48456 -1062 48472 -1028
rect 48515 -1034 48549 -1018
rect 47610 -1130 47640 -1080
rect 47550 -1250 47640 -1130
rect 48610 -1080 48618 -922
rect 48610 -1130 48640 -1080
rect 48680 -1130 48700 -890
rect 48610 -1250 48700 -1130
rect 52540 -570 52630 -440
rect 52540 -810 52560 -570
rect 52600 -612 52630 -570
rect 52620 -770 52630 -612
rect 53600 -570 53690 -440
rect 53600 -612 53630 -570
rect 52688 -674 52722 -658
rect 52756 -664 52772 -630
rect 52948 -664 52964 -630
rect 53254 -664 53270 -630
rect 53446 -664 53462 -630
rect 52688 -724 52722 -708
rect 53505 -674 53539 -658
rect 52756 -752 52772 -718
rect 52948 -752 52964 -718
rect 53254 -752 53270 -718
rect 53446 -752 53462 -718
rect 53505 -724 53539 -708
rect 52600 -810 52630 -770
rect 52540 -870 52630 -810
rect 52540 -1130 52560 -870
rect 52600 -922 52630 -870
rect 52620 -1080 52630 -922
rect 53600 -770 53608 -612
rect 53600 -810 53630 -770
rect 53670 -810 53690 -570
rect 53600 -890 53690 -810
rect 53600 -922 53630 -890
rect 52688 -984 52722 -968
rect 52756 -974 52772 -940
rect 52948 -974 52964 -940
rect 53254 -974 53270 -940
rect 53446 -974 53462 -940
rect 52688 -1034 52722 -1018
rect 53505 -984 53539 -968
rect 52756 -1062 52772 -1028
rect 52948 -1062 52964 -1028
rect 53254 -1062 53270 -1028
rect 53446 -1062 53462 -1028
rect 53505 -1034 53539 -1018
rect 52600 -1130 52630 -1080
rect 52540 -1250 52630 -1130
rect 53600 -1080 53608 -922
rect 53600 -1130 53630 -1080
rect 53670 -1130 53690 -890
rect 53600 -1250 53690 -1130
rect 57530 -570 57620 -440
rect 57530 -810 57550 -570
rect 57590 -612 57620 -570
rect 57610 -770 57620 -612
rect 58590 -570 58680 -440
rect 58590 -612 58620 -570
rect 57678 -674 57712 -658
rect 57746 -664 57762 -630
rect 57938 -664 57954 -630
rect 58244 -664 58260 -630
rect 58436 -664 58452 -630
rect 57678 -724 57712 -708
rect 58495 -674 58529 -658
rect 57746 -752 57762 -718
rect 57938 -752 57954 -718
rect 58244 -752 58260 -718
rect 58436 -752 58452 -718
rect 58495 -724 58529 -708
rect 57590 -810 57620 -770
rect 57530 -870 57620 -810
rect 57530 -1130 57550 -870
rect 57590 -922 57620 -870
rect 57610 -1080 57620 -922
rect 58590 -770 58598 -612
rect 58590 -810 58620 -770
rect 58660 -810 58680 -570
rect 58590 -890 58680 -810
rect 58590 -922 58620 -890
rect 57678 -984 57712 -968
rect 57746 -974 57762 -940
rect 57938 -974 57954 -940
rect 58244 -974 58260 -940
rect 58436 -974 58452 -940
rect 57678 -1034 57712 -1018
rect 58495 -984 58529 -968
rect 57746 -1062 57762 -1028
rect 57938 -1062 57954 -1028
rect 58244 -1062 58260 -1028
rect 58436 -1062 58452 -1028
rect 58495 -1034 58529 -1018
rect 57590 -1130 57620 -1080
rect 57530 -1250 57620 -1130
rect 58590 -1080 58598 -922
rect 58590 -1130 58620 -1080
rect 58660 -1130 58680 -890
rect 58590 -1250 58680 -1130
rect 62520 -570 62610 -440
rect 62520 -810 62540 -570
rect 62580 -612 62610 -570
rect 62600 -770 62610 -612
rect 63580 -570 63670 -440
rect 63580 -612 63610 -570
rect 62668 -674 62702 -658
rect 62736 -664 62752 -630
rect 62928 -664 62944 -630
rect 63234 -664 63250 -630
rect 63426 -664 63442 -630
rect 62668 -724 62702 -708
rect 63485 -674 63519 -658
rect 62736 -752 62752 -718
rect 62928 -752 62944 -718
rect 63234 -752 63250 -718
rect 63426 -752 63442 -718
rect 63485 -724 63519 -708
rect 62580 -810 62610 -770
rect 62520 -870 62610 -810
rect 62520 -1130 62540 -870
rect 62580 -922 62610 -870
rect 62600 -1080 62610 -922
rect 63580 -770 63588 -612
rect 63580 -810 63610 -770
rect 63650 -810 63670 -570
rect 63580 -890 63670 -810
rect 63580 -922 63610 -890
rect 62668 -984 62702 -968
rect 62736 -974 62752 -940
rect 62928 -974 62944 -940
rect 63234 -974 63250 -940
rect 63426 -974 63442 -940
rect 62668 -1034 62702 -1018
rect 63485 -984 63519 -968
rect 62736 -1062 62752 -1028
rect 62928 -1062 62944 -1028
rect 63234 -1062 63250 -1028
rect 63426 -1062 63442 -1028
rect 63485 -1034 63519 -1018
rect 62580 -1130 62610 -1080
rect 62520 -1250 62610 -1130
rect 63580 -1080 63588 -922
rect 63580 -1130 63610 -1080
rect 63650 -1130 63670 -890
rect 63580 -1250 63670 -1130
rect 67510 -570 67600 -440
rect 67510 -810 67530 -570
rect 67570 -612 67600 -570
rect 67590 -770 67600 -612
rect 68570 -570 68660 -440
rect 68570 -612 68600 -570
rect 67658 -674 67692 -658
rect 67726 -664 67742 -630
rect 67918 -664 67934 -630
rect 68224 -664 68240 -630
rect 68416 -664 68432 -630
rect 67658 -724 67692 -708
rect 68475 -674 68509 -658
rect 67726 -752 67742 -718
rect 67918 -752 67934 -718
rect 68224 -752 68240 -718
rect 68416 -752 68432 -718
rect 68475 -724 68509 -708
rect 67570 -810 67600 -770
rect 67510 -870 67600 -810
rect 67510 -1130 67530 -870
rect 67570 -922 67600 -870
rect 67590 -1080 67600 -922
rect 68570 -770 68578 -612
rect 68570 -810 68600 -770
rect 68640 -810 68660 -570
rect 68570 -890 68660 -810
rect 68570 -922 68600 -890
rect 67658 -984 67692 -968
rect 67726 -974 67742 -940
rect 67918 -974 67934 -940
rect 68224 -974 68240 -940
rect 68416 -974 68432 -940
rect 67658 -1034 67692 -1018
rect 68475 -984 68509 -968
rect 67726 -1062 67742 -1028
rect 67918 -1062 67934 -1028
rect 68224 -1062 68240 -1028
rect 68416 -1062 68432 -1028
rect 68475 -1034 68509 -1018
rect 67570 -1130 67600 -1080
rect 67510 -1250 67600 -1130
rect 68570 -1080 68578 -922
rect 68570 -1130 68600 -1080
rect 68640 -1130 68660 -890
rect 68570 -1250 68660 -1130
rect 72500 -570 72590 -440
rect 72500 -810 72520 -570
rect 72560 -612 72590 -570
rect 72580 -770 72590 -612
rect 73560 -570 73650 -440
rect 73560 -612 73590 -570
rect 72648 -674 72682 -658
rect 72716 -664 72732 -630
rect 72908 -664 72924 -630
rect 73214 -664 73230 -630
rect 73406 -664 73422 -630
rect 72648 -724 72682 -708
rect 73465 -674 73499 -658
rect 72716 -752 72732 -718
rect 72908 -752 72924 -718
rect 73214 -752 73230 -718
rect 73406 -752 73422 -718
rect 73465 -724 73499 -708
rect 72560 -810 72590 -770
rect 72500 -870 72590 -810
rect 72500 -1130 72520 -870
rect 72560 -922 72590 -870
rect 72580 -1080 72590 -922
rect 73560 -770 73568 -612
rect 73560 -810 73590 -770
rect 73630 -810 73650 -570
rect 73560 -890 73650 -810
rect 73560 -922 73590 -890
rect 72648 -984 72682 -968
rect 72716 -974 72732 -940
rect 72908 -974 72924 -940
rect 73214 -974 73230 -940
rect 73406 -974 73422 -940
rect 72648 -1034 72682 -1018
rect 73465 -984 73499 -968
rect 72716 -1062 72732 -1028
rect 72908 -1062 72924 -1028
rect 73214 -1062 73230 -1028
rect 73406 -1062 73422 -1028
rect 73465 -1034 73499 -1018
rect 72560 -1130 72590 -1080
rect 72500 -1250 72590 -1130
rect 73560 -1080 73568 -922
rect 73560 -1130 73590 -1080
rect 73630 -1130 73650 -890
rect 73560 -1250 73650 -1130
rect 77490 -570 77580 -440
rect 77490 -810 77510 -570
rect 77550 -612 77580 -570
rect 77570 -770 77580 -612
rect 78550 -570 78640 -440
rect 78550 -612 78580 -570
rect 77638 -674 77672 -658
rect 77706 -664 77722 -630
rect 77898 -664 77914 -630
rect 78204 -664 78220 -630
rect 78396 -664 78412 -630
rect 77638 -724 77672 -708
rect 78455 -674 78489 -658
rect 77706 -752 77722 -718
rect 77898 -752 77914 -718
rect 78204 -752 78220 -718
rect 78396 -752 78412 -718
rect 78455 -724 78489 -708
rect 77550 -810 77580 -770
rect 77490 -870 77580 -810
rect 77490 -1130 77510 -870
rect 77550 -922 77580 -870
rect 77570 -1080 77580 -922
rect 78550 -770 78558 -612
rect 78550 -810 78580 -770
rect 78620 -810 78640 -570
rect 78550 -890 78640 -810
rect 78550 -922 78580 -890
rect 77638 -984 77672 -968
rect 77706 -974 77722 -940
rect 77898 -974 77914 -940
rect 78204 -974 78220 -940
rect 78396 -974 78412 -940
rect 77638 -1034 77672 -1018
rect 78455 -984 78489 -968
rect 77706 -1062 77722 -1028
rect 77898 -1062 77914 -1028
rect 78204 -1062 78220 -1028
rect 78396 -1062 78412 -1028
rect 78455 -1034 78489 -1018
rect 77550 -1130 77580 -1080
rect 77490 -1250 77580 -1130
rect 78550 -1080 78558 -922
rect 78550 -1130 78580 -1080
rect 78620 -1130 78640 -890
rect 78550 -1250 78640 -1130
rect 82210 -570 82300 -440
rect 82210 -810 82230 -570
rect 82270 -612 82300 -570
rect 82290 -770 82300 -612
rect 83270 -570 83360 -440
rect 83270 -612 83300 -570
rect 82358 -674 82392 -658
rect 82426 -664 82442 -630
rect 82618 -664 82634 -630
rect 82924 -664 82940 -630
rect 83116 -664 83132 -630
rect 82358 -724 82392 -708
rect 83175 -674 83209 -658
rect 82426 -752 82442 -718
rect 82618 -752 82634 -718
rect 82924 -752 82940 -718
rect 83116 -752 83132 -718
rect 83175 -724 83209 -708
rect 82270 -810 82300 -770
rect 82210 -870 82300 -810
rect 82210 -1130 82230 -870
rect 82270 -922 82300 -870
rect 82290 -1080 82300 -922
rect 83270 -770 83278 -612
rect 83270 -810 83300 -770
rect 83340 -810 83360 -570
rect 83270 -890 83360 -810
rect 83270 -922 83300 -890
rect 82358 -984 82392 -968
rect 82426 -974 82442 -940
rect 82618 -974 82634 -940
rect 82924 -974 82940 -940
rect 83116 -974 83132 -940
rect 82358 -1034 82392 -1018
rect 83175 -984 83209 -968
rect 82426 -1062 82442 -1028
rect 82618 -1062 82634 -1028
rect 82924 -1062 82940 -1028
rect 83116 -1062 83132 -1028
rect 83175 -1034 83209 -1018
rect 82270 -1130 82300 -1080
rect 82210 -1250 82300 -1130
rect 83270 -1080 83278 -922
rect 83270 -1130 83300 -1080
rect 83340 -1130 83360 -890
rect 83270 -1250 83360 -1130
<< viali >>
rect 2660 28458 2700 28500
rect 2660 28300 2686 28458
rect 2686 28300 2700 28458
rect 3730 28458 3770 28500
rect 2872 28406 3048 28440
rect 3370 28406 3546 28440
rect 2788 28362 2822 28396
rect 3605 28362 3639 28396
rect 2872 28318 3048 28352
rect 3370 28318 3546 28352
rect 2660 28260 2700 28300
rect 2660 28148 2700 28200
rect 2660 27990 2686 28148
rect 2686 27990 2700 28148
rect 3730 28300 3742 28458
rect 3742 28300 3770 28458
rect 3730 28260 3770 28300
rect 3730 28148 3770 28180
rect 2872 28096 3048 28130
rect 3370 28096 3546 28130
rect 2788 28052 2822 28086
rect 3605 28052 3639 28086
rect 2872 28008 3048 28042
rect 3370 28008 3546 28042
rect 2660 27940 2700 27990
rect 3730 27990 3742 28148
rect 3742 27990 3770 28148
rect 3730 27940 3770 27990
rect 7650 28458 7690 28500
rect 7650 28300 7676 28458
rect 7676 28300 7690 28458
rect 8720 28458 8760 28500
rect 7862 28406 8038 28440
rect 8360 28406 8536 28440
rect 7778 28362 7812 28396
rect 8595 28362 8629 28396
rect 7862 28318 8038 28352
rect 8360 28318 8536 28352
rect 7650 28260 7690 28300
rect 7650 28148 7690 28200
rect 7650 27990 7676 28148
rect 7676 27990 7690 28148
rect 8720 28300 8732 28458
rect 8732 28300 8760 28458
rect 8720 28260 8760 28300
rect 8720 28148 8760 28180
rect 7862 28096 8038 28130
rect 8360 28096 8536 28130
rect 7778 28052 7812 28086
rect 8595 28052 8629 28086
rect 7862 28008 8038 28042
rect 8360 28008 8536 28042
rect 7650 27940 7690 27990
rect 8720 27990 8732 28148
rect 8732 27990 8760 28148
rect 8720 27940 8760 27990
rect 12640 28458 12680 28500
rect 12640 28300 12666 28458
rect 12666 28300 12680 28458
rect 13710 28458 13750 28500
rect 12852 28406 13028 28440
rect 13350 28406 13526 28440
rect 12768 28362 12802 28396
rect 13585 28362 13619 28396
rect 12852 28318 13028 28352
rect 13350 28318 13526 28352
rect 12640 28260 12680 28300
rect 12640 28148 12680 28200
rect 12640 27990 12666 28148
rect 12666 27990 12680 28148
rect 13710 28300 13722 28458
rect 13722 28300 13750 28458
rect 13710 28260 13750 28300
rect 13710 28148 13750 28180
rect 12852 28096 13028 28130
rect 13350 28096 13526 28130
rect 12768 28052 12802 28086
rect 13585 28052 13619 28086
rect 12852 28008 13028 28042
rect 13350 28008 13526 28042
rect 12640 27940 12680 27990
rect 13710 27990 13722 28148
rect 13722 27990 13750 28148
rect 13710 27940 13750 27990
rect 17630 28458 17670 28500
rect 17630 28300 17656 28458
rect 17656 28300 17670 28458
rect 18700 28458 18740 28500
rect 17842 28406 18018 28440
rect 18340 28406 18516 28440
rect 17758 28362 17792 28396
rect 18575 28362 18609 28396
rect 17842 28318 18018 28352
rect 18340 28318 18516 28352
rect 17630 28260 17670 28300
rect 17630 28148 17670 28200
rect 17630 27990 17656 28148
rect 17656 27990 17670 28148
rect 18700 28300 18712 28458
rect 18712 28300 18740 28458
rect 18700 28260 18740 28300
rect 18700 28148 18740 28180
rect 17842 28096 18018 28130
rect 18340 28096 18516 28130
rect 17758 28052 17792 28086
rect 18575 28052 18609 28086
rect 17842 28008 18018 28042
rect 18340 28008 18516 28042
rect 17630 27940 17670 27990
rect 18700 27990 18712 28148
rect 18712 27990 18740 28148
rect 18700 27940 18740 27990
rect 22620 28458 22660 28500
rect 22620 28300 22646 28458
rect 22646 28300 22660 28458
rect 23690 28458 23730 28500
rect 22832 28406 23008 28440
rect 23330 28406 23506 28440
rect 22748 28362 22782 28396
rect 23565 28362 23599 28396
rect 22832 28318 23008 28352
rect 23330 28318 23506 28352
rect 22620 28260 22660 28300
rect 22620 28148 22660 28200
rect 22620 27990 22646 28148
rect 22646 27990 22660 28148
rect 23690 28300 23702 28458
rect 23702 28300 23730 28458
rect 23690 28260 23730 28300
rect 23690 28148 23730 28180
rect 22832 28096 23008 28130
rect 23330 28096 23506 28130
rect 22748 28052 22782 28086
rect 23565 28052 23599 28086
rect 22832 28008 23008 28042
rect 23330 28008 23506 28042
rect 22620 27940 22660 27990
rect 23690 27990 23702 28148
rect 23702 27990 23730 28148
rect 23690 27940 23730 27990
rect 27610 28458 27650 28500
rect 27610 28300 27636 28458
rect 27636 28300 27650 28458
rect 28680 28458 28720 28500
rect 27822 28406 27998 28440
rect 28320 28406 28496 28440
rect 27738 28362 27772 28396
rect 28555 28362 28589 28396
rect 27822 28318 27998 28352
rect 28320 28318 28496 28352
rect 27610 28260 27650 28300
rect 27610 28148 27650 28200
rect 27610 27990 27636 28148
rect 27636 27990 27650 28148
rect 28680 28300 28692 28458
rect 28692 28300 28720 28458
rect 28680 28260 28720 28300
rect 28680 28148 28720 28180
rect 27822 28096 27998 28130
rect 28320 28096 28496 28130
rect 27738 28052 27772 28086
rect 28555 28052 28589 28086
rect 27822 28008 27998 28042
rect 28320 28008 28496 28042
rect 27610 27940 27650 27990
rect 28680 27990 28692 28148
rect 28692 27990 28720 28148
rect 28680 27940 28720 27990
rect 32600 28458 32640 28500
rect 32600 28300 32626 28458
rect 32626 28300 32640 28458
rect 33670 28458 33710 28500
rect 32812 28406 32988 28440
rect 33310 28406 33486 28440
rect 32728 28362 32762 28396
rect 33545 28362 33579 28396
rect 32812 28318 32988 28352
rect 33310 28318 33486 28352
rect 32600 28260 32640 28300
rect 32600 28148 32640 28200
rect 32600 27990 32626 28148
rect 32626 27990 32640 28148
rect 33670 28300 33682 28458
rect 33682 28300 33710 28458
rect 33670 28260 33710 28300
rect 33670 28148 33710 28180
rect 32812 28096 32988 28130
rect 33310 28096 33486 28130
rect 32728 28052 32762 28086
rect 33545 28052 33579 28086
rect 32812 28008 32988 28042
rect 33310 28008 33486 28042
rect 32600 27940 32640 27990
rect 33670 27990 33682 28148
rect 33682 27990 33710 28148
rect 33670 27940 33710 27990
rect 37590 28458 37630 28500
rect 37590 28300 37616 28458
rect 37616 28300 37630 28458
rect 38660 28458 38700 28500
rect 37802 28406 37978 28440
rect 38300 28406 38476 28440
rect 37718 28362 37752 28396
rect 38535 28362 38569 28396
rect 37802 28318 37978 28352
rect 38300 28318 38476 28352
rect 37590 28260 37630 28300
rect 37590 28148 37630 28200
rect 37590 27990 37616 28148
rect 37616 27990 37630 28148
rect 38660 28300 38672 28458
rect 38672 28300 38700 28458
rect 38660 28260 38700 28300
rect 38660 28148 38700 28180
rect 37802 28096 37978 28130
rect 38300 28096 38476 28130
rect 37718 28052 37752 28086
rect 38535 28052 38569 28086
rect 37802 28008 37978 28042
rect 38300 28008 38476 28042
rect 37590 27940 37630 27990
rect 38660 27990 38672 28148
rect 38672 27990 38700 28148
rect 38660 27940 38700 27990
rect 42580 28458 42620 28500
rect 42580 28300 42606 28458
rect 42606 28300 42620 28458
rect 43650 28458 43690 28500
rect 42792 28406 42968 28440
rect 43290 28406 43466 28440
rect 42708 28362 42742 28396
rect 43525 28362 43559 28396
rect 42792 28318 42968 28352
rect 43290 28318 43466 28352
rect 42580 28260 42620 28300
rect 42580 28148 42620 28200
rect 42580 27990 42606 28148
rect 42606 27990 42620 28148
rect 43650 28300 43662 28458
rect 43662 28300 43690 28458
rect 43650 28260 43690 28300
rect 43650 28148 43690 28180
rect 42792 28096 42968 28130
rect 43290 28096 43466 28130
rect 42708 28052 42742 28086
rect 43525 28052 43559 28086
rect 42792 28008 42968 28042
rect 43290 28008 43466 28042
rect 42580 27940 42620 27990
rect 43650 27990 43662 28148
rect 43662 27990 43690 28148
rect 43650 27940 43690 27990
rect 47570 28458 47610 28500
rect 47570 28300 47596 28458
rect 47596 28300 47610 28458
rect 48640 28458 48680 28500
rect 47782 28406 47958 28440
rect 48280 28406 48456 28440
rect 47698 28362 47732 28396
rect 48515 28362 48549 28396
rect 47782 28318 47958 28352
rect 48280 28318 48456 28352
rect 47570 28260 47610 28300
rect 47570 28148 47610 28200
rect 47570 27990 47596 28148
rect 47596 27990 47610 28148
rect 48640 28300 48652 28458
rect 48652 28300 48680 28458
rect 48640 28260 48680 28300
rect 48640 28148 48680 28180
rect 47782 28096 47958 28130
rect 48280 28096 48456 28130
rect 47698 28052 47732 28086
rect 48515 28052 48549 28086
rect 47782 28008 47958 28042
rect 48280 28008 48456 28042
rect 47570 27940 47610 27990
rect 48640 27990 48652 28148
rect 48652 27990 48680 28148
rect 48640 27940 48680 27990
rect 52560 28458 52600 28500
rect 52560 28300 52586 28458
rect 52586 28300 52600 28458
rect 53630 28458 53670 28500
rect 52772 28406 52948 28440
rect 53270 28406 53446 28440
rect 52688 28362 52722 28396
rect 53505 28362 53539 28396
rect 52772 28318 52948 28352
rect 53270 28318 53446 28352
rect 52560 28260 52600 28300
rect 52560 28148 52600 28200
rect 52560 27990 52586 28148
rect 52586 27990 52600 28148
rect 53630 28300 53642 28458
rect 53642 28300 53670 28458
rect 53630 28260 53670 28300
rect 53630 28148 53670 28180
rect 52772 28096 52948 28130
rect 53270 28096 53446 28130
rect 52688 28052 52722 28086
rect 53505 28052 53539 28086
rect 52772 28008 52948 28042
rect 53270 28008 53446 28042
rect 52560 27940 52600 27990
rect 53630 27990 53642 28148
rect 53642 27990 53670 28148
rect 53630 27940 53670 27990
rect 57550 28458 57590 28500
rect 57550 28300 57576 28458
rect 57576 28300 57590 28458
rect 58620 28458 58660 28500
rect 57762 28406 57938 28440
rect 58260 28406 58436 28440
rect 57678 28362 57712 28396
rect 58495 28362 58529 28396
rect 57762 28318 57938 28352
rect 58260 28318 58436 28352
rect 57550 28260 57590 28300
rect 57550 28148 57590 28200
rect 57550 27990 57576 28148
rect 57576 27990 57590 28148
rect 58620 28300 58632 28458
rect 58632 28300 58660 28458
rect 58620 28260 58660 28300
rect 58620 28148 58660 28180
rect 57762 28096 57938 28130
rect 58260 28096 58436 28130
rect 57678 28052 57712 28086
rect 58495 28052 58529 28086
rect 57762 28008 57938 28042
rect 58260 28008 58436 28042
rect 57550 27940 57590 27990
rect 58620 27990 58632 28148
rect 58632 27990 58660 28148
rect 58620 27940 58660 27990
rect 62540 28458 62580 28500
rect 62540 28300 62566 28458
rect 62566 28300 62580 28458
rect 63610 28458 63650 28500
rect 62752 28406 62928 28440
rect 63250 28406 63426 28440
rect 62668 28362 62702 28396
rect 63485 28362 63519 28396
rect 62752 28318 62928 28352
rect 63250 28318 63426 28352
rect 62540 28260 62580 28300
rect 62540 28148 62580 28200
rect 62540 27990 62566 28148
rect 62566 27990 62580 28148
rect 63610 28300 63622 28458
rect 63622 28300 63650 28458
rect 63610 28260 63650 28300
rect 63610 28148 63650 28180
rect 62752 28096 62928 28130
rect 63250 28096 63426 28130
rect 62668 28052 62702 28086
rect 63485 28052 63519 28086
rect 62752 28008 62928 28042
rect 63250 28008 63426 28042
rect 62540 27940 62580 27990
rect 63610 27990 63622 28148
rect 63622 27990 63650 28148
rect 63610 27940 63650 27990
rect 67530 28458 67570 28500
rect 67530 28300 67556 28458
rect 67556 28300 67570 28458
rect 68600 28458 68640 28500
rect 67742 28406 67918 28440
rect 68240 28406 68416 28440
rect 67658 28362 67692 28396
rect 68475 28362 68509 28396
rect 67742 28318 67918 28352
rect 68240 28318 68416 28352
rect 67530 28260 67570 28300
rect 67530 28148 67570 28200
rect 67530 27990 67556 28148
rect 67556 27990 67570 28148
rect 68600 28300 68612 28458
rect 68612 28300 68640 28458
rect 68600 28260 68640 28300
rect 68600 28148 68640 28180
rect 67742 28096 67918 28130
rect 68240 28096 68416 28130
rect 67658 28052 67692 28086
rect 68475 28052 68509 28086
rect 67742 28008 67918 28042
rect 68240 28008 68416 28042
rect 67530 27940 67570 27990
rect 68600 27990 68612 28148
rect 68612 27990 68640 28148
rect 68600 27940 68640 27990
rect 72520 28458 72560 28500
rect 72520 28300 72546 28458
rect 72546 28300 72560 28458
rect 73590 28458 73630 28500
rect 72732 28406 72908 28440
rect 73230 28406 73406 28440
rect 72648 28362 72682 28396
rect 73465 28362 73499 28396
rect 72732 28318 72908 28352
rect 73230 28318 73406 28352
rect 72520 28260 72560 28300
rect 72520 28148 72560 28200
rect 72520 27990 72546 28148
rect 72546 27990 72560 28148
rect 73590 28300 73602 28458
rect 73602 28300 73630 28458
rect 73590 28260 73630 28300
rect 73590 28148 73630 28180
rect 72732 28096 72908 28130
rect 73230 28096 73406 28130
rect 72648 28052 72682 28086
rect 73465 28052 73499 28086
rect 72732 28008 72908 28042
rect 73230 28008 73406 28042
rect 72520 27940 72560 27990
rect 73590 27990 73602 28148
rect 73602 27990 73630 28148
rect 73590 27940 73630 27990
rect 77510 28458 77550 28500
rect 77510 28300 77536 28458
rect 77536 28300 77550 28458
rect 78580 28458 78620 28500
rect 77722 28406 77898 28440
rect 78220 28406 78396 28440
rect 77638 28362 77672 28396
rect 78455 28362 78489 28396
rect 77722 28318 77898 28352
rect 78220 28318 78396 28352
rect 77510 28260 77550 28300
rect 77510 28148 77550 28200
rect 77510 27990 77536 28148
rect 77536 27990 77550 28148
rect 78580 28300 78592 28458
rect 78592 28300 78620 28458
rect 78580 28260 78620 28300
rect 78580 28148 78620 28180
rect 77722 28096 77898 28130
rect 78220 28096 78396 28130
rect 77638 28052 77672 28086
rect 78455 28052 78489 28086
rect 77722 28008 77898 28042
rect 78220 28008 78396 28042
rect 77510 27940 77550 27990
rect 78580 27990 78592 28148
rect 78592 27990 78620 28148
rect 78580 27940 78620 27990
rect 82230 28458 82270 28500
rect 82230 28300 82256 28458
rect 82256 28300 82270 28458
rect 83300 28458 83340 28500
rect 82442 28406 82618 28440
rect 82940 28406 83116 28440
rect 82358 28362 82392 28396
rect 83175 28362 83209 28396
rect 82442 28318 82618 28352
rect 82940 28318 83116 28352
rect 82230 28260 82270 28300
rect 82230 28148 82270 28200
rect 82230 27990 82256 28148
rect 82256 27990 82270 28148
rect 83300 28300 83312 28458
rect 83312 28300 83340 28458
rect 83300 28260 83340 28300
rect 83300 28148 83340 28180
rect 82442 28096 82618 28130
rect 82940 28096 83116 28130
rect 82358 28052 82392 28086
rect 83175 28052 83209 28086
rect 82442 28008 82618 28042
rect 82940 28008 83116 28042
rect 82230 27940 82270 27990
rect 83300 27990 83312 28148
rect 83312 27990 83340 28148
rect 83300 27940 83340 27990
rect 82230 26748 82270 26790
rect 82230 26590 82256 26748
rect 82256 26590 82270 26748
rect 83300 26748 83340 26790
rect 82442 26696 82618 26730
rect 82940 26696 83116 26730
rect 82358 26652 82392 26686
rect 83175 26652 83209 26686
rect 82442 26608 82618 26642
rect 82940 26608 83116 26642
rect 82230 26550 82270 26590
rect 82230 26438 82270 26490
rect 82230 26280 82256 26438
rect 82256 26280 82270 26438
rect 83300 26590 83312 26748
rect 83312 26590 83340 26748
rect 83300 26550 83340 26590
rect 83300 26438 83340 26470
rect 82442 26386 82618 26420
rect 82940 26386 83116 26420
rect 82358 26342 82392 26376
rect 83175 26342 83209 26376
rect 82442 26298 82618 26332
rect 82940 26298 83116 26332
rect 82230 26230 82270 26280
rect 83300 26280 83312 26438
rect 83312 26280 83340 26438
rect 83300 26230 83340 26280
rect 82230 25038 82270 25080
rect 82230 24880 82256 25038
rect 82256 24880 82270 25038
rect 83300 25038 83340 25080
rect 82442 24986 82618 25020
rect 82940 24986 83116 25020
rect 82358 24942 82392 24976
rect 83175 24942 83209 24976
rect 82442 24898 82618 24932
rect 82940 24898 83116 24932
rect 82230 24840 82270 24880
rect 82230 24728 82270 24780
rect 82230 24570 82256 24728
rect 82256 24570 82270 24728
rect 83300 24880 83312 25038
rect 83312 24880 83340 25038
rect 83300 24840 83340 24880
rect 83300 24728 83340 24760
rect 82442 24676 82618 24710
rect 82940 24676 83116 24710
rect 82358 24632 82392 24666
rect 83175 24632 83209 24666
rect 82442 24588 82618 24622
rect 82940 24588 83116 24622
rect 82230 24520 82270 24570
rect 83300 24570 83312 24728
rect 83312 24570 83340 24728
rect 83300 24520 83340 24570
rect -2060 23328 -2020 23370
rect -2060 23170 -2034 23328
rect -2034 23170 -2020 23328
rect -990 23328 -950 23370
rect -1848 23276 -1672 23310
rect -1350 23276 -1174 23310
rect -1932 23232 -1898 23266
rect -1115 23232 -1081 23266
rect -1848 23188 -1672 23222
rect -1350 23188 -1174 23222
rect -2060 23130 -2020 23170
rect -2060 23018 -2020 23070
rect -2060 22860 -2034 23018
rect -2034 22860 -2020 23018
rect -990 23170 -978 23328
rect -978 23170 -950 23328
rect -990 23130 -950 23170
rect -990 23018 -950 23050
rect -1848 22966 -1672 23000
rect -1350 22966 -1174 23000
rect -1932 22922 -1898 22956
rect -1115 22922 -1081 22956
rect -1848 22878 -1672 22912
rect -1350 22878 -1174 22912
rect -2060 22810 -2020 22860
rect -990 22860 -978 23018
rect -978 22860 -950 23018
rect -990 22810 -950 22860
rect 82230 23328 82270 23370
rect 82230 23170 82256 23328
rect 82256 23170 82270 23328
rect 83300 23328 83340 23370
rect 82442 23276 82618 23310
rect 82940 23276 83116 23310
rect 82358 23232 82392 23266
rect 83175 23232 83209 23266
rect 82442 23188 82618 23222
rect 82940 23188 83116 23222
rect 82230 23130 82270 23170
rect 82230 23018 82270 23070
rect 82230 22860 82256 23018
rect 82256 22860 82270 23018
rect 83300 23170 83312 23328
rect 83312 23170 83340 23328
rect 83300 23130 83340 23170
rect 83300 23018 83340 23050
rect 82442 22966 82618 23000
rect 82940 22966 83116 23000
rect 82358 22922 82392 22956
rect 83175 22922 83209 22956
rect 82442 22878 82618 22912
rect 82940 22878 83116 22912
rect 82230 22810 82270 22860
rect 83300 22860 83312 23018
rect 83312 22860 83340 23018
rect 83300 22810 83340 22860
rect -2060 21618 -2020 21660
rect -2060 21460 -2034 21618
rect -2034 21460 -2020 21618
rect -990 21618 -950 21660
rect -1848 21566 -1672 21600
rect -1350 21566 -1174 21600
rect -1932 21522 -1898 21556
rect -1115 21522 -1081 21556
rect -1848 21478 -1672 21512
rect -1350 21478 -1174 21512
rect -2060 21420 -2020 21460
rect -2060 21308 -2020 21360
rect -2060 21150 -2034 21308
rect -2034 21150 -2020 21308
rect -990 21460 -978 21618
rect -978 21460 -950 21618
rect -990 21420 -950 21460
rect -990 21308 -950 21340
rect -1848 21256 -1672 21290
rect -1350 21256 -1174 21290
rect -1932 21212 -1898 21246
rect -1115 21212 -1081 21246
rect -1848 21168 -1672 21202
rect -1350 21168 -1174 21202
rect -2060 21100 -2020 21150
rect -990 21150 -978 21308
rect -978 21150 -950 21308
rect -990 21100 -950 21150
rect 82230 21618 82270 21660
rect 82230 21460 82256 21618
rect 82256 21460 82270 21618
rect 83300 21618 83340 21660
rect 82442 21566 82618 21600
rect 82940 21566 83116 21600
rect 82358 21522 82392 21556
rect 83175 21522 83209 21556
rect 82442 21478 82618 21512
rect 82940 21478 83116 21512
rect 82230 21420 82270 21460
rect 82230 21308 82270 21360
rect 82230 21150 82256 21308
rect 82256 21150 82270 21308
rect 83300 21460 83312 21618
rect 83312 21460 83340 21618
rect 83300 21420 83340 21460
rect 83300 21308 83340 21340
rect 82442 21256 82618 21290
rect 82940 21256 83116 21290
rect 82358 21212 82392 21246
rect 83175 21212 83209 21246
rect 82442 21168 82618 21202
rect 82940 21168 83116 21202
rect 82230 21100 82270 21150
rect 83300 21150 83312 21308
rect 83312 21150 83340 21308
rect 83300 21100 83340 21150
rect -2060 19908 -2020 19950
rect -2060 19750 -2034 19908
rect -2034 19750 -2020 19908
rect -990 19908 -950 19950
rect -1848 19856 -1672 19890
rect -1350 19856 -1174 19890
rect -1932 19812 -1898 19846
rect -1115 19812 -1081 19846
rect -1848 19768 -1672 19802
rect -1350 19768 -1174 19802
rect -2060 19710 -2020 19750
rect -2060 19598 -2020 19650
rect -2060 19440 -2034 19598
rect -2034 19440 -2020 19598
rect -990 19750 -978 19908
rect -978 19750 -950 19908
rect -990 19710 -950 19750
rect -990 19598 -950 19630
rect -1848 19546 -1672 19580
rect -1350 19546 -1174 19580
rect -1932 19502 -1898 19536
rect -1115 19502 -1081 19536
rect -1848 19458 -1672 19492
rect -1350 19458 -1174 19492
rect -2060 19390 -2020 19440
rect -990 19440 -978 19598
rect -978 19440 -950 19598
rect -990 19390 -950 19440
rect 82230 19908 82270 19950
rect 82230 19750 82256 19908
rect 82256 19750 82270 19908
rect 83300 19908 83340 19950
rect 82442 19856 82618 19890
rect 82940 19856 83116 19890
rect 82358 19812 82392 19846
rect 83175 19812 83209 19846
rect 82442 19768 82618 19802
rect 82940 19768 83116 19802
rect 82230 19710 82270 19750
rect 82230 19598 82270 19650
rect 82230 19440 82256 19598
rect 82256 19440 82270 19598
rect 83300 19750 83312 19908
rect 83312 19750 83340 19908
rect 83300 19710 83340 19750
rect 83300 19598 83340 19630
rect 82442 19546 82618 19580
rect 82940 19546 83116 19580
rect 82358 19502 82392 19536
rect 83175 19502 83209 19536
rect 82442 19458 82618 19492
rect 82940 19458 83116 19492
rect 82230 19390 82270 19440
rect 83300 19440 83312 19598
rect 83312 19440 83340 19598
rect 83300 19390 83340 19440
rect -2060 18198 -2020 18240
rect -2060 18040 -2034 18198
rect -2034 18040 -2020 18198
rect -990 18198 -950 18240
rect -1848 18146 -1672 18180
rect -1350 18146 -1174 18180
rect -1932 18102 -1898 18136
rect -1115 18102 -1081 18136
rect -1848 18058 -1672 18092
rect -1350 18058 -1174 18092
rect -2060 18000 -2020 18040
rect -2060 17888 -2020 17940
rect -2060 17730 -2034 17888
rect -2034 17730 -2020 17888
rect -990 18040 -978 18198
rect -978 18040 -950 18198
rect -990 18000 -950 18040
rect -990 17888 -950 17920
rect -1848 17836 -1672 17870
rect -1350 17836 -1174 17870
rect -1932 17792 -1898 17826
rect -1115 17792 -1081 17826
rect -1848 17748 -1672 17782
rect -1350 17748 -1174 17782
rect -2060 17680 -2020 17730
rect -990 17730 -978 17888
rect -978 17730 -950 17888
rect -990 17680 -950 17730
rect 82230 18198 82270 18240
rect 82230 18040 82256 18198
rect 82256 18040 82270 18198
rect 83300 18198 83340 18240
rect 82442 18146 82618 18180
rect 82940 18146 83116 18180
rect 82358 18102 82392 18136
rect 83175 18102 83209 18136
rect 82442 18058 82618 18092
rect 82940 18058 83116 18092
rect 82230 18000 82270 18040
rect 82230 17888 82270 17940
rect 82230 17730 82256 17888
rect 82256 17730 82270 17888
rect 83300 18040 83312 18198
rect 83312 18040 83340 18198
rect 83300 18000 83340 18040
rect 83300 17888 83340 17920
rect 82442 17836 82618 17870
rect 82940 17836 83116 17870
rect 82358 17792 82392 17826
rect 83175 17792 83209 17826
rect 82442 17748 82618 17782
rect 82940 17748 83116 17782
rect 82230 17680 82270 17730
rect 83300 17730 83312 17888
rect 83312 17730 83340 17888
rect 83300 17680 83340 17730
rect -2060 16488 -2020 16530
rect -2060 16330 -2034 16488
rect -2034 16330 -2020 16488
rect -990 16488 -950 16530
rect -1848 16436 -1672 16470
rect -1350 16436 -1174 16470
rect -1932 16392 -1898 16426
rect -1115 16392 -1081 16426
rect -1848 16348 -1672 16382
rect -1350 16348 -1174 16382
rect -2060 16290 -2020 16330
rect -2060 16178 -2020 16230
rect -2060 16020 -2034 16178
rect -2034 16020 -2020 16178
rect -990 16330 -978 16488
rect -978 16330 -950 16488
rect -990 16290 -950 16330
rect -990 16178 -950 16210
rect -1848 16126 -1672 16160
rect -1350 16126 -1174 16160
rect -1932 16082 -1898 16116
rect -1115 16082 -1081 16116
rect -1848 16038 -1672 16072
rect -1350 16038 -1174 16072
rect -2060 15970 -2020 16020
rect -990 16020 -978 16178
rect -978 16020 -950 16178
rect -990 15970 -950 16020
rect 82230 16488 82270 16530
rect 82230 16330 82256 16488
rect 82256 16330 82270 16488
rect 83300 16488 83340 16530
rect 82442 16436 82618 16470
rect 82940 16436 83116 16470
rect 82358 16392 82392 16426
rect 83175 16392 83209 16426
rect 82442 16348 82618 16382
rect 82940 16348 83116 16382
rect 82230 16290 82270 16330
rect 82230 16178 82270 16230
rect 82230 16020 82256 16178
rect 82256 16020 82270 16178
rect 83300 16330 83312 16488
rect 83312 16330 83340 16488
rect 83300 16290 83340 16330
rect 83300 16178 83340 16210
rect 82442 16126 82618 16160
rect 82940 16126 83116 16160
rect 82358 16082 82392 16116
rect 83175 16082 83209 16116
rect 82442 16038 82618 16072
rect 82940 16038 83116 16072
rect 82230 15970 82270 16020
rect 83300 16020 83312 16178
rect 83312 16020 83340 16178
rect 83300 15970 83340 16020
rect -2060 14778 -2020 14820
rect -2060 14620 -2034 14778
rect -2034 14620 -2020 14778
rect -990 14778 -950 14820
rect -1848 14726 -1672 14760
rect -1350 14726 -1174 14760
rect -1932 14682 -1898 14716
rect -1115 14682 -1081 14716
rect -1848 14638 -1672 14672
rect -1350 14638 -1174 14672
rect -2060 14580 -2020 14620
rect -2060 14468 -2020 14520
rect -2060 14310 -2034 14468
rect -2034 14310 -2020 14468
rect -990 14620 -978 14778
rect -978 14620 -950 14778
rect -990 14580 -950 14620
rect -990 14468 -950 14500
rect -1848 14416 -1672 14450
rect -1350 14416 -1174 14450
rect -1932 14372 -1898 14406
rect -1115 14372 -1081 14406
rect -1848 14328 -1672 14362
rect -1350 14328 -1174 14362
rect -2060 14260 -2020 14310
rect -990 14310 -978 14468
rect -978 14310 -950 14468
rect -990 14260 -950 14310
rect 82230 14778 82270 14820
rect 82230 14620 82256 14778
rect 82256 14620 82270 14778
rect 83300 14778 83340 14820
rect 82442 14726 82618 14760
rect 82940 14726 83116 14760
rect 82358 14682 82392 14716
rect 83175 14682 83209 14716
rect 82442 14638 82618 14672
rect 82940 14638 83116 14672
rect 82230 14580 82270 14620
rect 82230 14468 82270 14520
rect 82230 14310 82256 14468
rect 82256 14310 82270 14468
rect 83300 14620 83312 14778
rect 83312 14620 83340 14778
rect 83300 14580 83340 14620
rect 83300 14468 83340 14500
rect 82442 14416 82618 14450
rect 82940 14416 83116 14450
rect 82358 14372 82392 14406
rect 83175 14372 83209 14406
rect 82442 14328 82618 14362
rect 82940 14328 83116 14362
rect 82230 14260 82270 14310
rect 83300 14310 83312 14468
rect 83312 14310 83340 14468
rect 83300 14260 83340 14310
rect -2060 13068 -2020 13110
rect -2060 12910 -2034 13068
rect -2034 12910 -2020 13068
rect -990 13068 -950 13110
rect -1848 13016 -1672 13050
rect -1350 13016 -1174 13050
rect -1932 12972 -1898 13006
rect -1115 12972 -1081 13006
rect -1848 12928 -1672 12962
rect -1350 12928 -1174 12962
rect -2060 12870 -2020 12910
rect -2060 12758 -2020 12810
rect -2060 12600 -2034 12758
rect -2034 12600 -2020 12758
rect -990 12910 -978 13068
rect -978 12910 -950 13068
rect -990 12870 -950 12910
rect -990 12758 -950 12790
rect -1848 12706 -1672 12740
rect -1350 12706 -1174 12740
rect -1932 12662 -1898 12696
rect -1115 12662 -1081 12696
rect -1848 12618 -1672 12652
rect -1350 12618 -1174 12652
rect -2060 12550 -2020 12600
rect -990 12600 -978 12758
rect -978 12600 -950 12758
rect -990 12550 -950 12600
rect 82230 13068 82270 13110
rect 82230 12910 82256 13068
rect 82256 12910 82270 13068
rect 83300 13068 83340 13110
rect 82442 13016 82618 13050
rect 82940 13016 83116 13050
rect 82358 12972 82392 13006
rect 83175 12972 83209 13006
rect 82442 12928 82618 12962
rect 82940 12928 83116 12962
rect 82230 12870 82270 12910
rect 82230 12758 82270 12810
rect 82230 12600 82256 12758
rect 82256 12600 82270 12758
rect 83300 12910 83312 13068
rect 83312 12910 83340 13068
rect 83300 12870 83340 12910
rect 83300 12758 83340 12790
rect 82442 12706 82618 12740
rect 82940 12706 83116 12740
rect 82358 12662 82392 12696
rect 83175 12662 83209 12696
rect 82442 12618 82618 12652
rect 82940 12618 83116 12652
rect 82230 12550 82270 12600
rect 83300 12600 83312 12758
rect 83312 12600 83340 12758
rect 83300 12550 83340 12600
rect -2060 11358 -2020 11400
rect -2060 11200 -2034 11358
rect -2034 11200 -2020 11358
rect -990 11358 -950 11400
rect -1848 11306 -1672 11340
rect -1350 11306 -1174 11340
rect -1932 11262 -1898 11296
rect -1115 11262 -1081 11296
rect -1848 11218 -1672 11252
rect -1350 11218 -1174 11252
rect -2060 11160 -2020 11200
rect -2060 11048 -2020 11100
rect -2060 10890 -2034 11048
rect -2034 10890 -2020 11048
rect -990 11200 -978 11358
rect -978 11200 -950 11358
rect -990 11160 -950 11200
rect -990 11048 -950 11080
rect -1848 10996 -1672 11030
rect -1350 10996 -1174 11030
rect -1932 10952 -1898 10986
rect -1115 10952 -1081 10986
rect -1848 10908 -1672 10942
rect -1350 10908 -1174 10942
rect -2060 10840 -2020 10890
rect -990 10890 -978 11048
rect -978 10890 -950 11048
rect -990 10840 -950 10890
rect 82230 11358 82270 11400
rect 82230 11200 82256 11358
rect 82256 11200 82270 11358
rect 83300 11358 83340 11400
rect 82442 11306 82618 11340
rect 82940 11306 83116 11340
rect 82358 11262 82392 11296
rect 83175 11262 83209 11296
rect 82442 11218 82618 11252
rect 82940 11218 83116 11252
rect 82230 11160 82270 11200
rect 82230 11048 82270 11100
rect 82230 10890 82256 11048
rect 82256 10890 82270 11048
rect 83300 11200 83312 11358
rect 83312 11200 83340 11358
rect 83300 11160 83340 11200
rect 83300 11048 83340 11080
rect 82442 10996 82618 11030
rect 82940 10996 83116 11030
rect 82358 10952 82392 10986
rect 83175 10952 83209 10986
rect 82442 10908 82618 10942
rect 82940 10908 83116 10942
rect 82230 10840 82270 10890
rect 83300 10890 83312 11048
rect 83312 10890 83340 11048
rect 83300 10840 83340 10890
rect -2060 9648 -2020 9690
rect -2060 9490 -2034 9648
rect -2034 9490 -2020 9648
rect -990 9648 -950 9690
rect -1848 9596 -1672 9630
rect -1350 9596 -1174 9630
rect -1932 9552 -1898 9586
rect -1115 9552 -1081 9586
rect -1848 9508 -1672 9542
rect -1350 9508 -1174 9542
rect -2060 9450 -2020 9490
rect -2060 9338 -2020 9390
rect -2060 9180 -2034 9338
rect -2034 9180 -2020 9338
rect -990 9490 -978 9648
rect -978 9490 -950 9648
rect -990 9450 -950 9490
rect -990 9338 -950 9370
rect -1848 9286 -1672 9320
rect -1350 9286 -1174 9320
rect -1932 9242 -1898 9276
rect -1115 9242 -1081 9276
rect -1848 9198 -1672 9232
rect -1350 9198 -1174 9232
rect -2060 9130 -2020 9180
rect -990 9180 -978 9338
rect -978 9180 -950 9338
rect -990 9130 -950 9180
rect 82230 9648 82270 9690
rect 82230 9490 82256 9648
rect 82256 9490 82270 9648
rect 83300 9648 83340 9690
rect 82442 9596 82618 9630
rect 82940 9596 83116 9630
rect 82358 9552 82392 9586
rect 83175 9552 83209 9586
rect 82442 9508 82618 9542
rect 82940 9508 83116 9542
rect 82230 9450 82270 9490
rect 82230 9338 82270 9390
rect 82230 9180 82256 9338
rect 82256 9180 82270 9338
rect 83300 9490 83312 9648
rect 83312 9490 83340 9648
rect 83300 9450 83340 9490
rect 83300 9338 83340 9370
rect 82442 9286 82618 9320
rect 82940 9286 83116 9320
rect 82358 9242 82392 9276
rect 83175 9242 83209 9276
rect 82442 9198 82618 9232
rect 82940 9198 83116 9232
rect 82230 9130 82270 9180
rect 83300 9180 83312 9338
rect 83312 9180 83340 9338
rect 83300 9130 83340 9180
rect -2060 7938 -2020 7980
rect -2060 7780 -2034 7938
rect -2034 7780 -2020 7938
rect -990 7938 -950 7980
rect -1848 7886 -1672 7920
rect -1350 7886 -1174 7920
rect -1932 7842 -1898 7876
rect -1115 7842 -1081 7876
rect -1848 7798 -1672 7832
rect -1350 7798 -1174 7832
rect -2060 7740 -2020 7780
rect -2060 7628 -2020 7680
rect -2060 7470 -2034 7628
rect -2034 7470 -2020 7628
rect -990 7780 -978 7938
rect -978 7780 -950 7938
rect -990 7740 -950 7780
rect -990 7628 -950 7660
rect -1848 7576 -1672 7610
rect -1350 7576 -1174 7610
rect -1932 7532 -1898 7566
rect -1115 7532 -1081 7566
rect -1848 7488 -1672 7522
rect -1350 7488 -1174 7522
rect -2060 7420 -2020 7470
rect -990 7470 -978 7628
rect -978 7470 -950 7628
rect -990 7420 -950 7470
rect 82230 7938 82270 7980
rect 82230 7780 82256 7938
rect 82256 7780 82270 7938
rect 83300 7938 83340 7980
rect 82442 7886 82618 7920
rect 82940 7886 83116 7920
rect 82358 7842 82392 7876
rect 83175 7842 83209 7876
rect 82442 7798 82618 7832
rect 82940 7798 83116 7832
rect 82230 7740 82270 7780
rect 82230 7628 82270 7680
rect 82230 7470 82256 7628
rect 82256 7470 82270 7628
rect 83300 7780 83312 7938
rect 83312 7780 83340 7938
rect 83300 7740 83340 7780
rect 83300 7628 83340 7660
rect 82442 7576 82618 7610
rect 82940 7576 83116 7610
rect 82358 7532 82392 7566
rect 83175 7532 83209 7566
rect 82442 7488 82618 7522
rect 82940 7488 83116 7522
rect 82230 7420 82270 7470
rect 83300 7470 83312 7628
rect 83312 7470 83340 7628
rect 83300 7420 83340 7470
rect -2060 6228 -2020 6270
rect -2060 6070 -2034 6228
rect -2034 6070 -2020 6228
rect -990 6228 -950 6270
rect -1848 6176 -1672 6210
rect -1350 6176 -1174 6210
rect -1932 6132 -1898 6166
rect -1115 6132 -1081 6166
rect -1848 6088 -1672 6122
rect -1350 6088 -1174 6122
rect -2060 6030 -2020 6070
rect -2060 5918 -2020 5970
rect -2060 5760 -2034 5918
rect -2034 5760 -2020 5918
rect -990 6070 -978 6228
rect -978 6070 -950 6228
rect -990 6030 -950 6070
rect -990 5918 -950 5950
rect -1848 5866 -1672 5900
rect -1350 5866 -1174 5900
rect -1932 5822 -1898 5856
rect -1115 5822 -1081 5856
rect -1848 5778 -1672 5812
rect -1350 5778 -1174 5812
rect -2060 5710 -2020 5760
rect -990 5760 -978 5918
rect -978 5760 -950 5918
rect -990 5710 -950 5760
rect 82230 6228 82270 6270
rect 82230 6070 82256 6228
rect 82256 6070 82270 6228
rect 83300 6228 83340 6270
rect 82442 6176 82618 6210
rect 82940 6176 83116 6210
rect 82358 6132 82392 6166
rect 83175 6132 83209 6166
rect 82442 6088 82618 6122
rect 82940 6088 83116 6122
rect 82230 6030 82270 6070
rect 82230 5918 82270 5970
rect 82230 5760 82256 5918
rect 82256 5760 82270 5918
rect 83300 6070 83312 6228
rect 83312 6070 83340 6228
rect 83300 6030 83340 6070
rect 83300 5918 83340 5950
rect 82442 5866 82618 5900
rect 82940 5866 83116 5900
rect 82358 5822 82392 5856
rect 83175 5822 83209 5856
rect 82442 5778 82618 5812
rect 82940 5778 83116 5812
rect 82230 5710 82270 5760
rect 83300 5760 83312 5918
rect 83312 5760 83340 5918
rect 83300 5710 83340 5760
rect -2060 4518 -2020 4560
rect -2060 4360 -2034 4518
rect -2034 4360 -2020 4518
rect -990 4518 -950 4560
rect -1848 4466 -1672 4500
rect -1350 4466 -1174 4500
rect -1932 4422 -1898 4456
rect -1115 4422 -1081 4456
rect -1848 4378 -1672 4412
rect -1350 4378 -1174 4412
rect -2060 4320 -2020 4360
rect -2060 4208 -2020 4260
rect -2060 4050 -2034 4208
rect -2034 4050 -2020 4208
rect -990 4360 -978 4518
rect -978 4360 -950 4518
rect -990 4320 -950 4360
rect -990 4208 -950 4240
rect -1848 4156 -1672 4190
rect -1350 4156 -1174 4190
rect -1932 4112 -1898 4146
rect -1115 4112 -1081 4146
rect -1848 4068 -1672 4102
rect -1350 4068 -1174 4102
rect -2060 4000 -2020 4050
rect -990 4050 -978 4208
rect -978 4050 -950 4208
rect -990 4000 -950 4050
rect 82230 4518 82270 4560
rect 82230 4360 82256 4518
rect 82256 4360 82270 4518
rect 83300 4518 83340 4560
rect 82442 4466 82618 4500
rect 82940 4466 83116 4500
rect 82358 4422 82392 4456
rect 83175 4422 83209 4456
rect 82442 4378 82618 4412
rect 82940 4378 83116 4412
rect 82230 4320 82270 4360
rect 82230 4208 82270 4260
rect 82230 4050 82256 4208
rect 82256 4050 82270 4208
rect 83300 4360 83312 4518
rect 83312 4360 83340 4518
rect 83300 4320 83340 4360
rect 83300 4208 83340 4240
rect 82442 4156 82618 4190
rect 82940 4156 83116 4190
rect 82358 4112 82392 4146
rect 83175 4112 83209 4146
rect 82442 4068 82618 4102
rect 82940 4068 83116 4102
rect 82230 4000 82270 4050
rect 83300 4050 83312 4208
rect 83312 4050 83340 4208
rect 83300 4000 83340 4050
rect -2060 2808 -2020 2850
rect -2060 2650 -2034 2808
rect -2034 2650 -2020 2808
rect -990 2808 -950 2850
rect -1848 2756 -1672 2790
rect -1350 2756 -1174 2790
rect -1932 2712 -1898 2746
rect -1115 2712 -1081 2746
rect -1848 2668 -1672 2702
rect -1350 2668 -1174 2702
rect -2060 2610 -2020 2650
rect -2060 2498 -2020 2550
rect -2060 2340 -2034 2498
rect -2034 2340 -2020 2498
rect -990 2650 -978 2808
rect -978 2650 -950 2808
rect -990 2610 -950 2650
rect -990 2498 -950 2530
rect -1848 2446 -1672 2480
rect -1350 2446 -1174 2480
rect -1932 2402 -1898 2436
rect -1115 2402 -1081 2436
rect -1848 2358 -1672 2392
rect -1350 2358 -1174 2392
rect -2060 2290 -2020 2340
rect -990 2340 -978 2498
rect -978 2340 -950 2498
rect -990 2290 -950 2340
rect 82230 2808 82270 2850
rect 82230 2650 82256 2808
rect 82256 2650 82270 2808
rect 83300 2808 83340 2850
rect 82442 2756 82618 2790
rect 82940 2756 83116 2790
rect 82358 2712 82392 2746
rect 83175 2712 83209 2746
rect 82442 2668 82618 2702
rect 82940 2668 83116 2702
rect 82230 2610 82270 2650
rect 82230 2498 82270 2550
rect 82230 2340 82256 2498
rect 82256 2340 82270 2498
rect 83300 2650 83312 2808
rect 83312 2650 83340 2808
rect 83300 2610 83340 2650
rect 83300 2498 83340 2530
rect 82442 2446 82618 2480
rect 82940 2446 83116 2480
rect 82358 2402 82392 2436
rect 83175 2402 83209 2436
rect 82442 2358 82618 2392
rect 82940 2358 83116 2392
rect 82230 2290 82270 2340
rect 83300 2340 83312 2498
rect 83312 2340 83340 2498
rect 83300 2290 83340 2340
rect -2060 1098 -2020 1140
rect -2060 940 -2034 1098
rect -2034 940 -2020 1098
rect -990 1098 -950 1140
rect -1848 1046 -1672 1080
rect -1350 1046 -1174 1080
rect -1932 1002 -1898 1036
rect -1115 1002 -1081 1036
rect -1848 958 -1672 992
rect -1350 958 -1174 992
rect -2060 900 -2020 940
rect -2060 788 -2020 840
rect -2060 630 -2034 788
rect -2034 630 -2020 788
rect -990 940 -978 1098
rect -978 940 -950 1098
rect -990 900 -950 940
rect -990 788 -950 820
rect -1848 736 -1672 770
rect -1350 736 -1174 770
rect -1932 692 -1898 726
rect -1115 692 -1081 726
rect -1848 648 -1672 682
rect -1350 648 -1174 682
rect -2060 580 -2020 630
rect -990 630 -978 788
rect -978 630 -950 788
rect -990 580 -950 630
rect 82230 1098 82270 1140
rect 82230 940 82256 1098
rect 82256 940 82270 1098
rect 83300 1098 83340 1140
rect 82442 1046 82618 1080
rect 82940 1046 83116 1080
rect 82358 1002 82392 1036
rect 83175 1002 83209 1036
rect 82442 958 82618 992
rect 82940 958 83116 992
rect 82230 900 82270 940
rect 82230 788 82270 840
rect 82230 630 82256 788
rect 82256 630 82270 788
rect 83300 940 83312 1098
rect 83312 940 83340 1098
rect 83300 900 83340 940
rect 83300 788 83340 820
rect 82442 736 82618 770
rect 82940 736 83116 770
rect 82358 692 82392 726
rect 83175 692 83209 726
rect 82442 648 82618 682
rect 82940 648 83116 682
rect 82230 580 82270 630
rect 83300 630 83312 788
rect 83312 630 83340 788
rect 83300 580 83340 630
rect -2060 -612 -2020 -570
rect -2060 -770 -2034 -612
rect -2034 -770 -2020 -612
rect -990 -612 -950 -570
rect -1848 -664 -1672 -630
rect -1350 -664 -1174 -630
rect -1932 -708 -1898 -674
rect -1115 -708 -1081 -674
rect -1848 -752 -1672 -718
rect -1350 -752 -1174 -718
rect -2060 -810 -2020 -770
rect -2060 -922 -2020 -870
rect -2060 -1080 -2034 -922
rect -2034 -1080 -2020 -922
rect -990 -770 -978 -612
rect -978 -770 -950 -612
rect -990 -810 -950 -770
rect -990 -922 -950 -890
rect -1848 -974 -1672 -940
rect -1350 -974 -1174 -940
rect -1932 -1018 -1898 -984
rect -1115 -1018 -1081 -984
rect -1848 -1062 -1672 -1028
rect -1350 -1062 -1174 -1028
rect -2060 -1130 -2020 -1080
rect -990 -1080 -978 -922
rect -978 -1080 -950 -922
rect -990 -1130 -950 -1080
rect 2660 -612 2700 -570
rect 2660 -770 2686 -612
rect 2686 -770 2700 -612
rect 3730 -612 3770 -570
rect 2872 -664 3048 -630
rect 3370 -664 3546 -630
rect 2788 -708 2822 -674
rect 3605 -708 3639 -674
rect 2872 -752 3048 -718
rect 3370 -752 3546 -718
rect 2660 -810 2700 -770
rect 2660 -922 2700 -870
rect 2660 -1080 2686 -922
rect 2686 -1080 2700 -922
rect 3730 -770 3742 -612
rect 3742 -770 3770 -612
rect 3730 -810 3770 -770
rect 3730 -922 3770 -890
rect 2872 -974 3048 -940
rect 3370 -974 3546 -940
rect 2788 -1018 2822 -984
rect 3605 -1018 3639 -984
rect 2872 -1062 3048 -1028
rect 3370 -1062 3546 -1028
rect 2660 -1130 2700 -1080
rect 3730 -1080 3742 -922
rect 3742 -1080 3770 -922
rect 3730 -1130 3770 -1080
rect 7650 -612 7690 -570
rect 7650 -770 7676 -612
rect 7676 -770 7690 -612
rect 8720 -612 8760 -570
rect 7862 -664 8038 -630
rect 8360 -664 8536 -630
rect 7778 -708 7812 -674
rect 8595 -708 8629 -674
rect 7862 -752 8038 -718
rect 8360 -752 8536 -718
rect 7650 -810 7690 -770
rect 7650 -922 7690 -870
rect 7650 -1080 7676 -922
rect 7676 -1080 7690 -922
rect 8720 -770 8732 -612
rect 8732 -770 8760 -612
rect 8720 -810 8760 -770
rect 8720 -922 8760 -890
rect 7862 -974 8038 -940
rect 8360 -974 8536 -940
rect 7778 -1018 7812 -984
rect 8595 -1018 8629 -984
rect 7862 -1062 8038 -1028
rect 8360 -1062 8536 -1028
rect 7650 -1130 7690 -1080
rect 8720 -1080 8732 -922
rect 8732 -1080 8760 -922
rect 8720 -1130 8760 -1080
rect 12640 -612 12680 -570
rect 12640 -770 12666 -612
rect 12666 -770 12680 -612
rect 13710 -612 13750 -570
rect 12852 -664 13028 -630
rect 13350 -664 13526 -630
rect 12768 -708 12802 -674
rect 13585 -708 13619 -674
rect 12852 -752 13028 -718
rect 13350 -752 13526 -718
rect 12640 -810 12680 -770
rect 12640 -922 12680 -870
rect 12640 -1080 12666 -922
rect 12666 -1080 12680 -922
rect 13710 -770 13722 -612
rect 13722 -770 13750 -612
rect 13710 -810 13750 -770
rect 13710 -922 13750 -890
rect 12852 -974 13028 -940
rect 13350 -974 13526 -940
rect 12768 -1018 12802 -984
rect 13585 -1018 13619 -984
rect 12852 -1062 13028 -1028
rect 13350 -1062 13526 -1028
rect 12640 -1130 12680 -1080
rect 13710 -1080 13722 -922
rect 13722 -1080 13750 -922
rect 13710 -1130 13750 -1080
rect 17630 -612 17670 -570
rect 17630 -770 17656 -612
rect 17656 -770 17670 -612
rect 18700 -612 18740 -570
rect 17842 -664 18018 -630
rect 18340 -664 18516 -630
rect 17758 -708 17792 -674
rect 18575 -708 18609 -674
rect 17842 -752 18018 -718
rect 18340 -752 18516 -718
rect 17630 -810 17670 -770
rect 17630 -922 17670 -870
rect 17630 -1080 17656 -922
rect 17656 -1080 17670 -922
rect 18700 -770 18712 -612
rect 18712 -770 18740 -612
rect 18700 -810 18740 -770
rect 18700 -922 18740 -890
rect 17842 -974 18018 -940
rect 18340 -974 18516 -940
rect 17758 -1018 17792 -984
rect 18575 -1018 18609 -984
rect 17842 -1062 18018 -1028
rect 18340 -1062 18516 -1028
rect 17630 -1130 17670 -1080
rect 18700 -1080 18712 -922
rect 18712 -1080 18740 -922
rect 18700 -1130 18740 -1080
rect 22620 -612 22660 -570
rect 22620 -770 22646 -612
rect 22646 -770 22660 -612
rect 23690 -612 23730 -570
rect 22832 -664 23008 -630
rect 23330 -664 23506 -630
rect 22748 -708 22782 -674
rect 23565 -708 23599 -674
rect 22832 -752 23008 -718
rect 23330 -752 23506 -718
rect 22620 -810 22660 -770
rect 22620 -922 22660 -870
rect 22620 -1080 22646 -922
rect 22646 -1080 22660 -922
rect 23690 -770 23702 -612
rect 23702 -770 23730 -612
rect 23690 -810 23730 -770
rect 23690 -922 23730 -890
rect 22832 -974 23008 -940
rect 23330 -974 23506 -940
rect 22748 -1018 22782 -984
rect 23565 -1018 23599 -984
rect 22832 -1062 23008 -1028
rect 23330 -1062 23506 -1028
rect 22620 -1130 22660 -1080
rect 23690 -1080 23702 -922
rect 23702 -1080 23730 -922
rect 23690 -1130 23730 -1080
rect 27610 -612 27650 -570
rect 27610 -770 27636 -612
rect 27636 -770 27650 -612
rect 28680 -612 28720 -570
rect 27822 -664 27998 -630
rect 28320 -664 28496 -630
rect 27738 -708 27772 -674
rect 28555 -708 28589 -674
rect 27822 -752 27998 -718
rect 28320 -752 28496 -718
rect 27610 -810 27650 -770
rect 27610 -922 27650 -870
rect 27610 -1080 27636 -922
rect 27636 -1080 27650 -922
rect 28680 -770 28692 -612
rect 28692 -770 28720 -612
rect 28680 -810 28720 -770
rect 28680 -922 28720 -890
rect 27822 -974 27998 -940
rect 28320 -974 28496 -940
rect 27738 -1018 27772 -984
rect 28555 -1018 28589 -984
rect 27822 -1062 27998 -1028
rect 28320 -1062 28496 -1028
rect 27610 -1130 27650 -1080
rect 28680 -1080 28692 -922
rect 28692 -1080 28720 -922
rect 28680 -1130 28720 -1080
rect 32600 -612 32640 -570
rect 32600 -770 32626 -612
rect 32626 -770 32640 -612
rect 33670 -612 33710 -570
rect 32812 -664 32988 -630
rect 33310 -664 33486 -630
rect 32728 -708 32762 -674
rect 33545 -708 33579 -674
rect 32812 -752 32988 -718
rect 33310 -752 33486 -718
rect 32600 -810 32640 -770
rect 32600 -922 32640 -870
rect 32600 -1080 32626 -922
rect 32626 -1080 32640 -922
rect 33670 -770 33682 -612
rect 33682 -770 33710 -612
rect 33670 -810 33710 -770
rect 33670 -922 33710 -890
rect 32812 -974 32988 -940
rect 33310 -974 33486 -940
rect 32728 -1018 32762 -984
rect 33545 -1018 33579 -984
rect 32812 -1062 32988 -1028
rect 33310 -1062 33486 -1028
rect 32600 -1130 32640 -1080
rect 33670 -1080 33682 -922
rect 33682 -1080 33710 -922
rect 33670 -1130 33710 -1080
rect 37590 -612 37630 -570
rect 37590 -770 37616 -612
rect 37616 -770 37630 -612
rect 38660 -612 38700 -570
rect 37802 -664 37978 -630
rect 38300 -664 38476 -630
rect 37718 -708 37752 -674
rect 38535 -708 38569 -674
rect 37802 -752 37978 -718
rect 38300 -752 38476 -718
rect 37590 -810 37630 -770
rect 37590 -922 37630 -870
rect 37590 -1080 37616 -922
rect 37616 -1080 37630 -922
rect 38660 -770 38672 -612
rect 38672 -770 38700 -612
rect 38660 -810 38700 -770
rect 38660 -922 38700 -890
rect 37802 -974 37978 -940
rect 38300 -974 38476 -940
rect 37718 -1018 37752 -984
rect 38535 -1018 38569 -984
rect 37802 -1062 37978 -1028
rect 38300 -1062 38476 -1028
rect 37590 -1130 37630 -1080
rect 38660 -1080 38672 -922
rect 38672 -1080 38700 -922
rect 38660 -1130 38700 -1080
rect 42580 -612 42620 -570
rect 42580 -770 42606 -612
rect 42606 -770 42620 -612
rect 43650 -612 43690 -570
rect 42792 -664 42968 -630
rect 43290 -664 43466 -630
rect 42708 -708 42742 -674
rect 43525 -708 43559 -674
rect 42792 -752 42968 -718
rect 43290 -752 43466 -718
rect 42580 -810 42620 -770
rect 42580 -922 42620 -870
rect 42580 -1080 42606 -922
rect 42606 -1080 42620 -922
rect 43650 -770 43662 -612
rect 43662 -770 43690 -612
rect 43650 -810 43690 -770
rect 43650 -922 43690 -890
rect 42792 -974 42968 -940
rect 43290 -974 43466 -940
rect 42708 -1018 42742 -984
rect 43525 -1018 43559 -984
rect 42792 -1062 42968 -1028
rect 43290 -1062 43466 -1028
rect 42580 -1130 42620 -1080
rect 43650 -1080 43662 -922
rect 43662 -1080 43690 -922
rect 43650 -1130 43690 -1080
rect 47570 -612 47610 -570
rect 47570 -770 47596 -612
rect 47596 -770 47610 -612
rect 48640 -612 48680 -570
rect 47782 -664 47958 -630
rect 48280 -664 48456 -630
rect 47698 -708 47732 -674
rect 48515 -708 48549 -674
rect 47782 -752 47958 -718
rect 48280 -752 48456 -718
rect 47570 -810 47610 -770
rect 47570 -922 47610 -870
rect 47570 -1080 47596 -922
rect 47596 -1080 47610 -922
rect 48640 -770 48652 -612
rect 48652 -770 48680 -612
rect 48640 -810 48680 -770
rect 48640 -922 48680 -890
rect 47782 -974 47958 -940
rect 48280 -974 48456 -940
rect 47698 -1018 47732 -984
rect 48515 -1018 48549 -984
rect 47782 -1062 47958 -1028
rect 48280 -1062 48456 -1028
rect 47570 -1130 47610 -1080
rect 48640 -1080 48652 -922
rect 48652 -1080 48680 -922
rect 48640 -1130 48680 -1080
rect 52560 -612 52600 -570
rect 52560 -770 52586 -612
rect 52586 -770 52600 -612
rect 53630 -612 53670 -570
rect 52772 -664 52948 -630
rect 53270 -664 53446 -630
rect 52688 -708 52722 -674
rect 53505 -708 53539 -674
rect 52772 -752 52948 -718
rect 53270 -752 53446 -718
rect 52560 -810 52600 -770
rect 52560 -922 52600 -870
rect 52560 -1080 52586 -922
rect 52586 -1080 52600 -922
rect 53630 -770 53642 -612
rect 53642 -770 53670 -612
rect 53630 -810 53670 -770
rect 53630 -922 53670 -890
rect 52772 -974 52948 -940
rect 53270 -974 53446 -940
rect 52688 -1018 52722 -984
rect 53505 -1018 53539 -984
rect 52772 -1062 52948 -1028
rect 53270 -1062 53446 -1028
rect 52560 -1130 52600 -1080
rect 53630 -1080 53642 -922
rect 53642 -1080 53670 -922
rect 53630 -1130 53670 -1080
rect 57550 -612 57590 -570
rect 57550 -770 57576 -612
rect 57576 -770 57590 -612
rect 58620 -612 58660 -570
rect 57762 -664 57938 -630
rect 58260 -664 58436 -630
rect 57678 -708 57712 -674
rect 58495 -708 58529 -674
rect 57762 -752 57938 -718
rect 58260 -752 58436 -718
rect 57550 -810 57590 -770
rect 57550 -922 57590 -870
rect 57550 -1080 57576 -922
rect 57576 -1080 57590 -922
rect 58620 -770 58632 -612
rect 58632 -770 58660 -612
rect 58620 -810 58660 -770
rect 58620 -922 58660 -890
rect 57762 -974 57938 -940
rect 58260 -974 58436 -940
rect 57678 -1018 57712 -984
rect 58495 -1018 58529 -984
rect 57762 -1062 57938 -1028
rect 58260 -1062 58436 -1028
rect 57550 -1130 57590 -1080
rect 58620 -1080 58632 -922
rect 58632 -1080 58660 -922
rect 58620 -1130 58660 -1080
rect 62540 -612 62580 -570
rect 62540 -770 62566 -612
rect 62566 -770 62580 -612
rect 63610 -612 63650 -570
rect 62752 -664 62928 -630
rect 63250 -664 63426 -630
rect 62668 -708 62702 -674
rect 63485 -708 63519 -674
rect 62752 -752 62928 -718
rect 63250 -752 63426 -718
rect 62540 -810 62580 -770
rect 62540 -922 62580 -870
rect 62540 -1080 62566 -922
rect 62566 -1080 62580 -922
rect 63610 -770 63622 -612
rect 63622 -770 63650 -612
rect 63610 -810 63650 -770
rect 63610 -922 63650 -890
rect 62752 -974 62928 -940
rect 63250 -974 63426 -940
rect 62668 -1018 62702 -984
rect 63485 -1018 63519 -984
rect 62752 -1062 62928 -1028
rect 63250 -1062 63426 -1028
rect 62540 -1130 62580 -1080
rect 63610 -1080 63622 -922
rect 63622 -1080 63650 -922
rect 63610 -1130 63650 -1080
rect 67530 -612 67570 -570
rect 67530 -770 67556 -612
rect 67556 -770 67570 -612
rect 68600 -612 68640 -570
rect 67742 -664 67918 -630
rect 68240 -664 68416 -630
rect 67658 -708 67692 -674
rect 68475 -708 68509 -674
rect 67742 -752 67918 -718
rect 68240 -752 68416 -718
rect 67530 -810 67570 -770
rect 67530 -922 67570 -870
rect 67530 -1080 67556 -922
rect 67556 -1080 67570 -922
rect 68600 -770 68612 -612
rect 68612 -770 68640 -612
rect 68600 -810 68640 -770
rect 68600 -922 68640 -890
rect 67742 -974 67918 -940
rect 68240 -974 68416 -940
rect 67658 -1018 67692 -984
rect 68475 -1018 68509 -984
rect 67742 -1062 67918 -1028
rect 68240 -1062 68416 -1028
rect 67530 -1130 67570 -1080
rect 68600 -1080 68612 -922
rect 68612 -1080 68640 -922
rect 68600 -1130 68640 -1080
rect 72520 -612 72560 -570
rect 72520 -770 72546 -612
rect 72546 -770 72560 -612
rect 73590 -612 73630 -570
rect 72732 -664 72908 -630
rect 73230 -664 73406 -630
rect 72648 -708 72682 -674
rect 73465 -708 73499 -674
rect 72732 -752 72908 -718
rect 73230 -752 73406 -718
rect 72520 -810 72560 -770
rect 72520 -922 72560 -870
rect 72520 -1080 72546 -922
rect 72546 -1080 72560 -922
rect 73590 -770 73602 -612
rect 73602 -770 73630 -612
rect 73590 -810 73630 -770
rect 73590 -922 73630 -890
rect 72732 -974 72908 -940
rect 73230 -974 73406 -940
rect 72648 -1018 72682 -984
rect 73465 -1018 73499 -984
rect 72732 -1062 72908 -1028
rect 73230 -1062 73406 -1028
rect 72520 -1130 72560 -1080
rect 73590 -1080 73602 -922
rect 73602 -1080 73630 -922
rect 73590 -1130 73630 -1080
rect 77510 -612 77550 -570
rect 77510 -770 77536 -612
rect 77536 -770 77550 -612
rect 78580 -612 78620 -570
rect 77722 -664 77898 -630
rect 78220 -664 78396 -630
rect 77638 -708 77672 -674
rect 78455 -708 78489 -674
rect 77722 -752 77898 -718
rect 78220 -752 78396 -718
rect 77510 -810 77550 -770
rect 77510 -922 77550 -870
rect 77510 -1080 77536 -922
rect 77536 -1080 77550 -922
rect 78580 -770 78592 -612
rect 78592 -770 78620 -612
rect 78580 -810 78620 -770
rect 78580 -922 78620 -890
rect 77722 -974 77898 -940
rect 78220 -974 78396 -940
rect 77638 -1018 77672 -984
rect 78455 -1018 78489 -984
rect 77722 -1062 77898 -1028
rect 78220 -1062 78396 -1028
rect 77510 -1130 77550 -1080
rect 78580 -1080 78592 -922
rect 78592 -1080 78620 -922
rect 78580 -1130 78620 -1080
rect 82230 -612 82270 -570
rect 82230 -770 82256 -612
rect 82256 -770 82270 -612
rect 83300 -612 83340 -570
rect 82442 -664 82618 -630
rect 82940 -664 83116 -630
rect 82358 -708 82392 -674
rect 83175 -708 83209 -674
rect 82442 -752 82618 -718
rect 82940 -752 83116 -718
rect 82230 -810 82270 -770
rect 82230 -922 82270 -870
rect 82230 -1080 82256 -922
rect 82256 -1080 82270 -922
rect 83300 -770 83312 -612
rect 83312 -770 83340 -612
rect 83300 -810 83340 -770
rect 83300 -922 83340 -890
rect 82442 -974 82618 -940
rect 82940 -974 83116 -940
rect 82358 -1018 82392 -984
rect 83175 -1018 83209 -984
rect 82442 -1062 82618 -1028
rect 82940 -1062 83116 -1028
rect 82230 -1130 82270 -1080
rect 83300 -1080 83312 -922
rect 83312 -1080 83340 -922
rect 83300 -1130 83340 -1080
<< metal1 >>
rect 4150 32620 4160 32650
rect -5140 32590 4160 32620
rect 4220 32620 4230 32650
rect 9140 32620 9150 32650
rect 4220 32590 9150 32620
rect 9210 32620 9220 32650
rect 14130 32620 14140 32650
rect 9210 32590 14140 32620
rect 14200 32620 14210 32650
rect 19120 32620 19130 32650
rect 14200 32590 19130 32620
rect 19190 32620 19200 32650
rect 24110 32620 24120 32650
rect 19190 32590 24120 32620
rect 24180 32620 24190 32650
rect 29100 32620 29110 32650
rect 24180 32590 29110 32620
rect 29170 32620 29180 32650
rect 34090 32620 34100 32650
rect 29170 32590 34100 32620
rect 34160 32620 34170 32650
rect 39080 32620 39090 32650
rect 34160 32590 39090 32620
rect 39150 32620 39160 32650
rect 44070 32620 44080 32650
rect 39150 32590 44080 32620
rect 44140 32620 44150 32650
rect 49060 32620 49070 32650
rect 44140 32590 49070 32620
rect 49130 32620 49140 32650
rect 54050 32620 54060 32650
rect 49130 32590 54060 32620
rect 54120 32620 54130 32650
rect 59040 32620 59050 32650
rect 54120 32590 59050 32620
rect 59110 32620 59120 32650
rect 64030 32620 64040 32650
rect 59110 32590 64040 32620
rect 64100 32620 64110 32650
rect 69020 32620 69030 32650
rect 64100 32590 69030 32620
rect 69090 32620 69100 32650
rect 74010 32620 74020 32650
rect 69090 32590 74020 32620
rect 74080 32620 74090 32650
rect 79000 32620 79010 32650
rect 74080 32590 79010 32620
rect 79070 32620 79080 32650
rect 79070 32590 84650 32620
rect 2420 32480 2480 32520
rect 4090 32480 4100 32510
rect -5140 32450 4100 32480
rect 4160 32480 4170 32510
rect 7410 32480 7470 32520
rect 9080 32480 9090 32510
rect 4160 32450 9090 32480
rect 9150 32480 9160 32510
rect 12400 32480 12460 32520
rect 14070 32480 14080 32510
rect 9150 32450 14080 32480
rect 14140 32480 14150 32510
rect 17390 32480 17450 32520
rect 19060 32480 19070 32510
rect 14140 32450 19070 32480
rect 19130 32480 19140 32510
rect 22380 32480 22440 32520
rect 24050 32480 24060 32510
rect 19130 32450 24060 32480
rect 24120 32480 24130 32510
rect 27370 32480 27430 32520
rect 29040 32480 29050 32510
rect 24120 32450 29050 32480
rect 29110 32480 29120 32510
rect 32360 32480 32420 32520
rect 34030 32480 34040 32510
rect 29110 32450 34040 32480
rect 34100 32480 34110 32510
rect 37350 32480 37410 32520
rect 39020 32480 39030 32510
rect 34100 32450 39030 32480
rect 39090 32480 39100 32510
rect 42340 32480 42400 32520
rect 44010 32480 44020 32510
rect 39090 32450 44020 32480
rect 44080 32480 44090 32510
rect 47330 32480 47390 32520
rect 49000 32480 49010 32510
rect 44080 32450 49010 32480
rect 49070 32480 49080 32510
rect 52320 32480 52380 32520
rect 53990 32480 54000 32510
rect 49070 32450 54000 32480
rect 54060 32480 54070 32510
rect 57310 32480 57370 32520
rect 58980 32480 58990 32510
rect 54060 32450 58990 32480
rect 59050 32480 59060 32510
rect 62300 32480 62360 32520
rect 63970 32480 63980 32510
rect 59050 32450 63980 32480
rect 64040 32480 64050 32510
rect 67290 32480 67350 32520
rect 68960 32480 68970 32510
rect 64040 32450 68970 32480
rect 69030 32480 69040 32510
rect 72280 32480 72340 32520
rect 73950 32480 73960 32510
rect 69030 32450 73960 32480
rect 74020 32480 74030 32510
rect 77270 32480 77330 32520
rect 78940 32480 78950 32510
rect 74020 32450 78950 32480
rect 79010 32480 79020 32510
rect 79010 32450 84650 32480
rect 14310 32340 14320 32370
rect -5140 32310 14320 32340
rect 14380 32340 14390 32370
rect 19300 32340 19310 32370
rect 14380 32310 19310 32340
rect 19370 32340 19380 32370
rect 24290 32340 24300 32370
rect 19370 32310 24300 32340
rect 24360 32340 24370 32370
rect 29280 32340 29290 32370
rect 24360 32310 29290 32340
rect 29350 32340 29360 32370
rect 34270 32340 34280 32370
rect 29350 32310 34280 32340
rect 34340 32340 34350 32370
rect 39260 32340 39270 32370
rect 34340 32310 39270 32340
rect 39330 32340 39340 32370
rect 44250 32340 44260 32370
rect 39330 32310 44260 32340
rect 44320 32340 44330 32370
rect 49240 32340 49250 32370
rect 44320 32310 49250 32340
rect 49310 32340 49320 32370
rect 54230 32340 54240 32370
rect 49310 32310 54240 32340
rect 54300 32340 54310 32370
rect 59220 32340 59230 32370
rect 54300 32310 59230 32340
rect 59290 32340 59300 32370
rect 64210 32340 64220 32370
rect 59290 32310 64220 32340
rect 64280 32340 64290 32370
rect 69200 32340 69210 32370
rect 64280 32310 69210 32340
rect 69270 32340 69280 32370
rect 69270 32310 84650 32340
rect 12220 32200 12280 32240
rect 14250 32200 14260 32230
rect -5140 32170 14260 32200
rect 14320 32200 14330 32230
rect 17210 32200 17270 32240
rect 19240 32200 19250 32230
rect 14320 32170 19250 32200
rect 19310 32200 19320 32230
rect 22200 32200 22260 32240
rect 24230 32200 24240 32230
rect 19310 32170 24240 32200
rect 24300 32200 24310 32230
rect 27190 32200 27250 32240
rect 29220 32200 29230 32230
rect 24300 32170 29230 32200
rect 29290 32200 29300 32230
rect 32180 32200 32240 32240
rect 34210 32200 34220 32230
rect 29290 32170 34220 32200
rect 34280 32200 34290 32230
rect 37170 32200 37230 32240
rect 39200 32200 39210 32230
rect 34280 32170 39210 32200
rect 39270 32200 39280 32230
rect 42160 32200 42220 32240
rect 44190 32200 44200 32230
rect 39270 32170 44200 32200
rect 44260 32200 44270 32230
rect 47150 32200 47210 32240
rect 49180 32200 49190 32230
rect 44260 32170 49190 32200
rect 49250 32200 49260 32230
rect 52140 32200 52200 32240
rect 54170 32200 54180 32230
rect 49250 32170 54180 32200
rect 54240 32200 54250 32230
rect 57130 32200 57190 32240
rect 59160 32200 59170 32230
rect 54240 32170 59170 32200
rect 59230 32200 59240 32230
rect 62120 32200 62180 32240
rect 64150 32200 64160 32230
rect 59230 32170 64160 32200
rect 64220 32200 64230 32230
rect 67110 32200 67170 32240
rect 69140 32200 69150 32230
rect 64220 32170 69150 32200
rect 69210 32200 69220 32230
rect 69210 32170 84650 32200
rect 24650 32060 24660 32090
rect -5140 32030 24660 32060
rect 24720 32060 24730 32090
rect 29640 32060 29650 32090
rect 24720 32030 29650 32060
rect 29710 32060 29720 32090
rect 34450 32060 34460 32090
rect 29710 32030 34460 32060
rect 34520 32060 34530 32090
rect 39440 32060 39450 32090
rect 34520 32030 39450 32060
rect 39510 32060 39520 32090
rect 44430 32060 44440 32090
rect 39510 32030 44440 32060
rect 44500 32060 44510 32090
rect 49420 32060 49430 32090
rect 44500 32030 49430 32060
rect 49490 32060 49500 32090
rect 54590 32060 54600 32090
rect 49490 32030 54600 32060
rect 54660 32060 54670 32090
rect 59580 32060 59590 32090
rect 54660 32030 59590 32060
rect 59650 32060 59660 32090
rect 59650 32030 84650 32060
rect 21840 31920 21900 31960
rect 24590 31920 24600 31950
rect -5140 31890 24600 31920
rect 24660 31920 24670 31950
rect 26830 31920 26890 31960
rect 29580 31920 29590 31950
rect 24660 31890 29590 31920
rect 29650 31920 29660 31950
rect 32000 31920 32060 31960
rect 34390 31920 34400 31950
rect 29650 31890 34400 31920
rect 34460 31920 34470 31950
rect 36990 31920 37050 31960
rect 39380 31920 39390 31950
rect 34460 31890 39390 31920
rect 39450 31920 39460 31950
rect 41980 31920 42040 31960
rect 44370 31920 44380 31950
rect 39450 31890 44380 31920
rect 44440 31920 44450 31950
rect 46970 31920 47030 31960
rect 49360 31920 49370 31950
rect 44440 31890 49370 31920
rect 49430 31920 49440 31950
rect 51780 31920 51840 31960
rect 54530 31920 54540 31950
rect 49430 31890 54540 31920
rect 54600 31920 54610 31950
rect 56770 31920 56830 31960
rect 59520 31920 59530 31950
rect 54600 31890 59530 31920
rect 59590 31920 59600 31950
rect 59590 31890 84650 31920
rect 24470 31780 24480 31810
rect -5140 31750 24480 31780
rect 24540 31780 24550 31810
rect 29460 31780 29470 31810
rect 24540 31750 29470 31780
rect 29530 31780 29540 31810
rect 34630 31780 34640 31810
rect 29530 31750 34640 31780
rect 34700 31780 34710 31810
rect 39620 31780 39630 31810
rect 34700 31750 39630 31780
rect 39690 31780 39700 31810
rect 44610 31780 44620 31810
rect 39690 31750 44620 31780
rect 44680 31780 44690 31810
rect 49600 31780 49610 31810
rect 44680 31750 49610 31780
rect 49670 31780 49680 31810
rect 54410 31780 54420 31810
rect 49670 31750 54420 31780
rect 54480 31780 54490 31810
rect 59400 31780 59410 31810
rect 54480 31750 59410 31780
rect 59470 31780 59480 31810
rect 59470 31750 84650 31780
rect 22020 31640 22080 31680
rect 24410 31640 24420 31670
rect -5140 31610 24420 31640
rect 24480 31640 24490 31670
rect 27010 31640 27070 31680
rect 29400 31640 29410 31670
rect 24480 31610 29410 31640
rect 29470 31640 29480 31670
rect 31820 31640 31880 31680
rect 34570 31640 34580 31670
rect 29470 31610 34580 31640
rect 34640 31640 34650 31670
rect 36810 31640 36870 31680
rect 39560 31640 39570 31670
rect 34640 31610 39570 31640
rect 39630 31640 39640 31670
rect 41800 31640 41860 31680
rect 44550 31640 44560 31670
rect 39630 31610 44560 31640
rect 44620 31640 44630 31670
rect 46790 31640 46850 31680
rect 49540 31640 49550 31670
rect 44620 31610 49550 31640
rect 49610 31640 49620 31670
rect 51960 31640 52020 31680
rect 54350 31640 54360 31670
rect 49610 31610 54360 31640
rect 54420 31640 54430 31670
rect 56950 31640 57010 31680
rect 59340 31640 59350 31670
rect 54420 31610 59350 31640
rect 59410 31640 59420 31670
rect 59410 31610 84650 31640
rect 34990 31500 35000 31530
rect -5140 31470 35000 31500
rect 35060 31500 35070 31530
rect 39800 31500 39810 31530
rect 35060 31470 39810 31500
rect 39870 31500 39880 31530
rect 44790 31500 44800 31530
rect 39870 31470 44800 31500
rect 44860 31500 44870 31530
rect 49960 31500 49970 31530
rect 44860 31470 49970 31500
rect 50030 31500 50040 31530
rect 50030 31470 84650 31500
rect 31460 31360 31520 31400
rect 34930 31360 34940 31390
rect -5140 31330 34940 31360
rect 35000 31360 35010 31390
rect 36630 31360 36690 31400
rect 39740 31360 39750 31390
rect 35000 31330 39750 31360
rect 39810 31360 39820 31390
rect 41620 31360 41680 31400
rect 44730 31360 44740 31390
rect 39810 31330 44740 31360
rect 44800 31360 44810 31390
rect 46430 31360 46490 31400
rect 49900 31360 49910 31390
rect 44800 31330 49910 31360
rect 49970 31360 49980 31390
rect 49970 31330 84650 31360
rect 34810 31220 34820 31250
rect -5140 31190 34820 31220
rect 34880 31220 34890 31250
rect 49780 31220 49790 31250
rect 34880 31190 49790 31220
rect 49850 31220 49860 31250
rect 49850 31190 84650 31220
rect 31640 31080 31700 31120
rect 34750 31080 34760 31110
rect -5140 31050 34760 31080
rect 34820 31080 34830 31110
rect 46610 31080 46670 31120
rect 49720 31080 49730 31110
rect 34820 31050 49730 31080
rect 49790 31080 49800 31110
rect 49790 31050 84650 31080
rect 39980 30940 39990 30970
rect -5140 30910 39990 30940
rect 40050 30940 40060 30970
rect 45150 30940 45160 30970
rect 40050 30910 45160 30940
rect 45220 30940 45230 30970
rect 45220 30910 84650 30940
rect 36450 30800 36510 30840
rect 39920 30800 39930 30830
rect -5140 30770 39930 30800
rect 39990 30800 40000 30830
rect 45090 30800 45100 30830
rect 39990 30770 45100 30800
rect 45160 30800 45170 30830
rect 45160 30770 84650 30800
rect 45000 30660 45010 30690
rect -5140 30630 45010 30660
rect 45070 30660 45080 30690
rect 45070 30630 84650 30660
rect 44910 30520 44920 30550
rect -5140 30490 44920 30520
rect 44980 30520 44990 30550
rect 44980 30490 84650 30520
rect 36210 30380 36270 30420
rect 40160 30380 40170 30410
rect -5180 30370 40170 30380
rect -5580 30350 40170 30370
rect 40230 30380 40240 30410
rect 40230 30350 84650 30380
rect -5580 30340 -5140 30350
rect 36270 30240 36330 30280
rect 40090 30240 40100 30270
rect -5170 30230 40100 30240
rect -5580 30210 40100 30230
rect 40160 30240 40170 30270
rect 40160 30210 84650 30240
rect -5580 30200 -5140 30210
rect -5590 29950 -5560 30140
rect -5530 30120 -5430 30140
rect -5110 30120 -5100 30180
rect -5040 30150 84650 30180
rect -5040 30120 -5030 30150
rect -5530 30060 -5510 30120
rect -5450 30090 -5430 30120
rect 3860 30090 3870 30120
rect -5450 30060 3870 30090
rect 3930 30090 3940 30120
rect 8850 30090 8860 30120
rect 3930 30060 8860 30090
rect 8920 30090 8930 30120
rect 13840 30090 13850 30120
rect 8920 30060 13850 30090
rect 13910 30090 13920 30120
rect 18830 30090 18840 30120
rect 13910 30060 18840 30090
rect 18900 30090 18910 30120
rect 23820 30090 23830 30120
rect 18900 30060 23830 30090
rect 23890 30090 23900 30120
rect 28810 30090 28820 30120
rect 23890 30060 28820 30090
rect 28880 30090 28890 30120
rect 33800 30090 33810 30120
rect 28880 30060 33810 30090
rect 33870 30090 33880 30120
rect 38790 30090 38800 30120
rect 33870 30060 38800 30090
rect 38860 30090 38870 30120
rect 43780 30090 43790 30120
rect 38860 30060 43790 30090
rect 43850 30090 43860 30120
rect 48770 30090 48780 30120
rect 43850 30060 48780 30090
rect 48840 30090 48850 30120
rect 53760 30090 53770 30120
rect 48840 30060 53770 30090
rect 53830 30090 53840 30120
rect 58750 30090 58760 30120
rect 53830 30060 58760 30090
rect 58820 30090 58830 30120
rect 63740 30090 63750 30120
rect 58820 30060 63750 30090
rect 63810 30090 63820 30120
rect 68730 30090 68740 30120
rect 63810 30060 68740 30090
rect 68800 30090 68810 30120
rect 73720 30090 73730 30120
rect 68800 30060 73730 30090
rect 73790 30090 73800 30120
rect 78710 30090 78720 30120
rect 73790 30060 78720 30090
rect 78780 30090 78790 30120
rect 78780 30060 84650 30090
rect -5530 30040 -5430 30060
rect -5250 29990 -5170 30000
rect -5250 29950 -5240 29990
rect -5590 29930 -5240 29950
rect -5180 29930 -5170 29990
rect -5590 29920 -5170 29930
rect -5140 29920 84650 29950
rect -5370 29850 -5290 29860
rect -5370 29790 -5360 29850
rect -5300 29790 -5290 29850
rect -5370 29780 -5290 29790
rect -5370 29050 -5310 29780
rect 2350 29590 2410 29600
rect 2410 29530 2610 29550
rect 2350 29520 2610 29530
rect -2080 29080 -2070 29140
rect -2010 29080 -2000 29140
rect -2080 29070 -2000 29080
rect -5590 28990 -5310 29050
rect -940 27400 -930 27420
rect 1860 27360 1890 29070
rect 1980 27360 2010 29070
rect 2100 27360 2130 29070
rect 2220 27360 2250 29070
rect 2340 27360 2370 29070
rect 2460 27360 2490 29070
rect 2580 27360 2610 29520
rect 3710 29140 3790 29150
rect 2640 29080 2650 29140
rect 2710 29080 2720 29140
rect 2640 29070 2720 29080
rect 3710 29080 3720 29140
rect 3780 29080 3790 29140
rect 3710 29070 3790 29080
rect 2640 28960 2710 29070
rect 2640 28950 3790 28960
rect 2640 28890 2650 28950
rect 2710 28900 3790 28950
rect 2710 28890 2720 28900
rect 2640 28880 2720 28890
rect 2640 28500 2710 28880
rect 2640 28260 2660 28500
rect 2700 28260 2710 28500
rect 3720 28500 3790 28900
rect 3170 28480 3250 28490
rect 2860 28440 3060 28446
rect 3170 28440 3180 28480
rect 2750 28410 2830 28430
rect 2750 28350 2760 28410
rect 2820 28396 2830 28410
rect 2860 28406 2872 28440
rect 3048 28420 3180 28440
rect 3240 28440 3250 28480
rect 3358 28440 3558 28446
rect 3240 28420 3370 28440
rect 3048 28410 3370 28420
rect 3048 28406 3060 28410
rect 2860 28400 3060 28406
rect 3358 28406 3370 28410
rect 3546 28406 3558 28440
rect 3358 28400 3558 28406
rect 3590 28410 3670 28430
rect 2822 28362 2830 28396
rect 2820 28350 2830 28362
rect 2750 28330 2830 28350
rect 2860 28352 3060 28358
rect 2860 28318 2872 28352
rect 3048 28350 3060 28352
rect 3358 28352 3558 28358
rect 3358 28350 3370 28352
rect 3048 28320 3370 28350
rect 3048 28318 3060 28320
rect 2860 28312 3060 28318
rect 2640 28200 2710 28260
rect 2640 27940 2660 28200
rect 2700 27940 2710 28200
rect 3170 28310 3250 28320
rect 3358 28318 3370 28320
rect 3546 28318 3558 28352
rect 3590 28350 3600 28410
rect 3660 28350 3670 28410
rect 3590 28330 3670 28350
rect 3358 28312 3558 28318
rect 3170 28250 3180 28310
rect 3240 28250 3250 28310
rect 3170 28200 3250 28250
rect 3170 28140 3180 28200
rect 3240 28140 3250 28200
rect 2860 28130 3060 28136
rect 3170 28130 3250 28140
rect 3720 28260 3730 28500
rect 3770 28260 3790 28500
rect 3720 28180 3790 28260
rect 3358 28130 3558 28136
rect 2750 28100 2830 28120
rect 2750 28040 2760 28100
rect 2820 28086 2830 28100
rect 2860 28096 2872 28130
rect 3048 28100 3370 28130
rect 3048 28096 3060 28100
rect 2860 28090 3060 28096
rect 3358 28096 3370 28100
rect 3546 28096 3558 28130
rect 3358 28090 3558 28096
rect 3590 28100 3670 28120
rect 2822 28052 2830 28086
rect 2820 28040 2830 28052
rect 2750 28020 2830 28040
rect 2860 28042 3060 28048
rect 2860 28008 2872 28042
rect 3048 28040 3060 28042
rect 3358 28042 3558 28048
rect 3358 28040 3370 28042
rect 3048 28030 3370 28040
rect 3048 28010 3180 28030
rect 3048 28008 3060 28010
rect 2860 28002 3060 28008
rect 3170 27970 3180 28010
rect 3240 28010 3370 28030
rect 3240 27970 3250 28010
rect 3358 28008 3370 28010
rect 3546 28008 3558 28042
rect 3590 28040 3600 28100
rect 3660 28040 3670 28100
rect 3590 28020 3670 28040
rect 3358 28002 3558 28008
rect 3170 27960 3250 27970
rect 2640 27360 2710 27940
rect 3720 27940 3730 28180
rect 3770 27940 3790 28180
rect 3720 27530 3790 27940
rect 3780 27400 3790 27440
rect 3720 27360 3790 27390
rect 3820 27360 3850 29920
rect 4170 29590 4230 29600
rect 3970 29530 4170 29550
rect 3970 29520 4230 29530
rect 7340 29590 7400 29600
rect 7400 29530 7600 29550
rect 7340 29520 7600 29530
rect 3880 29140 3940 29150
rect 3880 29070 3940 29080
rect 3910 27360 3940 29070
rect 3970 27360 4000 29520
rect 4090 27360 4120 29070
rect 4210 27360 4240 29070
rect 4330 27360 4360 29070
rect 4450 27360 4480 29070
rect 4570 27360 4600 29070
rect 4690 27360 4720 29070
rect 6850 27360 6880 29070
rect 6970 27360 7000 29070
rect 7090 27360 7120 29070
rect 7210 27360 7240 29070
rect 7330 27360 7360 29070
rect 7450 27360 7480 29070
rect 7570 27360 7600 29520
rect 8700 29140 8780 29150
rect 7630 29080 7640 29140
rect 7700 29080 7710 29140
rect 7630 29070 7710 29080
rect 8700 29080 8710 29140
rect 8770 29080 8780 29140
rect 8700 29070 8780 29080
rect 7630 28960 7700 29070
rect 7630 28950 8780 28960
rect 7630 28890 7640 28950
rect 7700 28900 8780 28950
rect 7700 28890 7710 28900
rect 7630 28880 7710 28890
rect 7630 28500 7700 28880
rect 7630 28260 7650 28500
rect 7690 28260 7700 28500
rect 8710 28500 8780 28900
rect 8160 28480 8240 28490
rect 7850 28440 8050 28446
rect 8160 28440 8170 28480
rect 7740 28410 7820 28430
rect 7740 28350 7750 28410
rect 7810 28396 7820 28410
rect 7850 28406 7862 28440
rect 8038 28420 8170 28440
rect 8230 28440 8240 28480
rect 8348 28440 8548 28446
rect 8230 28420 8360 28440
rect 8038 28410 8360 28420
rect 8038 28406 8050 28410
rect 7850 28400 8050 28406
rect 8348 28406 8360 28410
rect 8536 28406 8548 28440
rect 8348 28400 8548 28406
rect 8580 28410 8660 28430
rect 7812 28362 7820 28396
rect 7810 28350 7820 28362
rect 7740 28330 7820 28350
rect 7850 28352 8050 28358
rect 7850 28318 7862 28352
rect 8038 28350 8050 28352
rect 8348 28352 8548 28358
rect 8348 28350 8360 28352
rect 8038 28320 8360 28350
rect 8038 28318 8050 28320
rect 7850 28312 8050 28318
rect 7630 28200 7700 28260
rect 7630 27940 7650 28200
rect 7690 27940 7700 28200
rect 8160 28310 8240 28320
rect 8348 28318 8360 28320
rect 8536 28318 8548 28352
rect 8580 28350 8590 28410
rect 8650 28350 8660 28410
rect 8580 28330 8660 28350
rect 8348 28312 8548 28318
rect 8160 28250 8170 28310
rect 8230 28250 8240 28310
rect 8160 28200 8240 28250
rect 8160 28140 8170 28200
rect 8230 28140 8240 28200
rect 7850 28130 8050 28136
rect 8160 28130 8240 28140
rect 8710 28260 8720 28500
rect 8760 28260 8780 28500
rect 8710 28180 8780 28260
rect 8348 28130 8548 28136
rect 7740 28100 7820 28120
rect 7740 28040 7750 28100
rect 7810 28086 7820 28100
rect 7850 28096 7862 28130
rect 8038 28100 8360 28130
rect 8038 28096 8050 28100
rect 7850 28090 8050 28096
rect 8348 28096 8360 28100
rect 8536 28096 8548 28130
rect 8348 28090 8548 28096
rect 8580 28100 8660 28120
rect 7812 28052 7820 28086
rect 7810 28040 7820 28052
rect 7740 28020 7820 28040
rect 7850 28042 8050 28048
rect 7850 28008 7862 28042
rect 8038 28040 8050 28042
rect 8348 28042 8548 28048
rect 8348 28040 8360 28042
rect 8038 28030 8360 28040
rect 8038 28010 8170 28030
rect 8038 28008 8050 28010
rect 7850 28002 8050 28008
rect 8160 27970 8170 28010
rect 8230 28010 8360 28030
rect 8230 27970 8240 28010
rect 8348 28008 8360 28010
rect 8536 28008 8548 28042
rect 8580 28040 8590 28100
rect 8650 28040 8660 28100
rect 8580 28020 8660 28040
rect 8348 28002 8548 28008
rect 8160 27960 8240 27970
rect 7630 27360 7700 27940
rect 8710 27940 8720 28180
rect 8760 27940 8780 28180
rect 8710 27530 8780 27940
rect 8770 27400 8780 27440
rect 8710 27360 8780 27390
rect 8810 27360 8840 29920
rect 9160 29590 9220 29600
rect 8960 29530 9160 29550
rect 12330 29590 12390 29600
rect 8960 29520 9220 29530
rect 12150 29530 12210 29540
rect 8870 29140 8930 29150
rect 8870 29070 8930 29080
rect 8900 27360 8930 29070
rect 8960 27360 8990 29520
rect 12390 29530 12590 29550
rect 12330 29520 12590 29530
rect 12210 29470 12470 29490
rect 12150 29460 12470 29470
rect 9080 27360 9110 29070
rect 9200 27360 9230 29070
rect 9320 27360 9350 29070
rect 9440 27360 9470 29070
rect 9560 27360 9590 29070
rect 9680 27360 9710 29070
rect 11840 27360 11870 29070
rect 11960 27360 11990 29070
rect 12080 27360 12110 29070
rect 12200 27360 12230 29070
rect 12320 27360 12350 29070
rect 12440 27360 12470 29460
rect 12560 27360 12590 29520
rect 13690 29140 13770 29150
rect 12620 29080 12630 29140
rect 12690 29080 12700 29140
rect 12620 29070 12700 29080
rect 13690 29080 13700 29140
rect 13760 29080 13770 29140
rect 13690 29070 13770 29080
rect 12620 28960 12690 29070
rect 12620 28950 13770 28960
rect 12620 28890 12630 28950
rect 12690 28900 13770 28950
rect 12690 28890 12700 28900
rect 12620 28880 12700 28890
rect 12620 28500 12690 28880
rect 12620 28260 12640 28500
rect 12680 28260 12690 28500
rect 13700 28500 13770 28900
rect 13150 28480 13230 28490
rect 12840 28440 13040 28446
rect 13150 28440 13160 28480
rect 12730 28410 12810 28430
rect 12730 28350 12740 28410
rect 12800 28396 12810 28410
rect 12840 28406 12852 28440
rect 13028 28420 13160 28440
rect 13220 28440 13230 28480
rect 13338 28440 13538 28446
rect 13220 28420 13350 28440
rect 13028 28410 13350 28420
rect 13028 28406 13040 28410
rect 12840 28400 13040 28406
rect 13338 28406 13350 28410
rect 13526 28406 13538 28440
rect 13338 28400 13538 28406
rect 13570 28410 13650 28430
rect 12802 28362 12810 28396
rect 12800 28350 12810 28362
rect 12730 28330 12810 28350
rect 12840 28352 13040 28358
rect 12840 28318 12852 28352
rect 13028 28350 13040 28352
rect 13338 28352 13538 28358
rect 13338 28350 13350 28352
rect 13028 28320 13350 28350
rect 13028 28318 13040 28320
rect 12840 28312 13040 28318
rect 12620 28200 12690 28260
rect 12620 27940 12640 28200
rect 12680 27940 12690 28200
rect 13150 28310 13230 28320
rect 13338 28318 13350 28320
rect 13526 28318 13538 28352
rect 13570 28350 13580 28410
rect 13640 28350 13650 28410
rect 13570 28330 13650 28350
rect 13338 28312 13538 28318
rect 13150 28250 13160 28310
rect 13220 28250 13230 28310
rect 13150 28200 13230 28250
rect 13150 28140 13160 28200
rect 13220 28140 13230 28200
rect 12840 28130 13040 28136
rect 13150 28130 13230 28140
rect 13700 28260 13710 28500
rect 13750 28260 13770 28500
rect 13700 28180 13770 28260
rect 13338 28130 13538 28136
rect 12730 28100 12810 28120
rect 12730 28040 12740 28100
rect 12800 28086 12810 28100
rect 12840 28096 12852 28130
rect 13028 28100 13350 28130
rect 13028 28096 13040 28100
rect 12840 28090 13040 28096
rect 13338 28096 13350 28100
rect 13526 28096 13538 28130
rect 13338 28090 13538 28096
rect 13570 28100 13650 28120
rect 12802 28052 12810 28086
rect 12800 28040 12810 28052
rect 12730 28020 12810 28040
rect 12840 28042 13040 28048
rect 12840 28008 12852 28042
rect 13028 28040 13040 28042
rect 13338 28042 13538 28048
rect 13338 28040 13350 28042
rect 13028 28030 13350 28040
rect 13028 28010 13160 28030
rect 13028 28008 13040 28010
rect 12840 28002 13040 28008
rect 13150 27970 13160 28010
rect 13220 28010 13350 28030
rect 13220 27970 13230 28010
rect 13338 28008 13350 28010
rect 13526 28008 13538 28042
rect 13570 28040 13580 28100
rect 13640 28040 13650 28100
rect 13570 28020 13650 28040
rect 13338 28002 13538 28008
rect 13150 27960 13230 27970
rect 12620 27360 12690 27940
rect 13700 27940 13710 28180
rect 13750 27940 13770 28180
rect 13700 27530 13770 27940
rect 13760 27400 13770 27440
rect 13700 27360 13770 27390
rect 13800 27360 13830 29920
rect 14150 29590 14210 29600
rect 13950 29530 14150 29550
rect 17320 29590 17380 29600
rect 13950 29520 14210 29530
rect 14330 29530 14390 29540
rect 13860 29140 13920 29150
rect 13860 29070 13920 29080
rect 13890 27360 13920 29070
rect 13950 27360 13980 29520
rect 14070 29470 14330 29490
rect 14070 29460 14390 29470
rect 17140 29530 17200 29540
rect 17380 29530 17580 29550
rect 17320 29520 17580 29530
rect 17200 29470 17460 29490
rect 17140 29460 17460 29470
rect 14070 27360 14100 29460
rect 14190 27360 14220 29070
rect 14310 27360 14340 29070
rect 14430 27360 14460 29070
rect 14550 27360 14580 29070
rect 14670 27360 14700 29070
rect 16830 27360 16860 29070
rect 16950 27360 16980 29070
rect 17070 27360 17100 29070
rect 17190 27360 17220 29070
rect 17310 27360 17340 29070
rect 17430 27360 17460 29460
rect 17550 27360 17580 29520
rect 18680 29140 18760 29150
rect 17610 29080 17620 29140
rect 17680 29080 17690 29140
rect 17610 29070 17690 29080
rect 18680 29080 18690 29140
rect 18750 29080 18760 29140
rect 18680 29070 18760 29080
rect 17610 28960 17680 29070
rect 17610 28950 18760 28960
rect 17610 28890 17620 28950
rect 17680 28900 18760 28950
rect 17680 28890 17690 28900
rect 17610 28880 17690 28890
rect 17610 28500 17680 28880
rect 17610 28260 17630 28500
rect 17670 28260 17680 28500
rect 18690 28500 18760 28900
rect 18140 28480 18220 28490
rect 17830 28440 18030 28446
rect 18140 28440 18150 28480
rect 17720 28410 17800 28430
rect 17720 28350 17730 28410
rect 17790 28396 17800 28410
rect 17830 28406 17842 28440
rect 18018 28420 18150 28440
rect 18210 28440 18220 28480
rect 18328 28440 18528 28446
rect 18210 28420 18340 28440
rect 18018 28410 18340 28420
rect 18018 28406 18030 28410
rect 17830 28400 18030 28406
rect 18328 28406 18340 28410
rect 18516 28406 18528 28440
rect 18328 28400 18528 28406
rect 18560 28410 18640 28430
rect 17792 28362 17800 28396
rect 17790 28350 17800 28362
rect 17720 28330 17800 28350
rect 17830 28352 18030 28358
rect 17830 28318 17842 28352
rect 18018 28350 18030 28352
rect 18328 28352 18528 28358
rect 18328 28350 18340 28352
rect 18018 28320 18340 28350
rect 18018 28318 18030 28320
rect 17830 28312 18030 28318
rect 17610 28200 17680 28260
rect 17610 27940 17630 28200
rect 17670 27940 17680 28200
rect 18140 28310 18220 28320
rect 18328 28318 18340 28320
rect 18516 28318 18528 28352
rect 18560 28350 18570 28410
rect 18630 28350 18640 28410
rect 18560 28330 18640 28350
rect 18328 28312 18528 28318
rect 18140 28250 18150 28310
rect 18210 28250 18220 28310
rect 18140 28200 18220 28250
rect 18140 28140 18150 28200
rect 18210 28140 18220 28200
rect 17830 28130 18030 28136
rect 18140 28130 18220 28140
rect 18690 28260 18700 28500
rect 18740 28260 18760 28500
rect 18690 28180 18760 28260
rect 18328 28130 18528 28136
rect 17720 28100 17800 28120
rect 17720 28040 17730 28100
rect 17790 28086 17800 28100
rect 17830 28096 17842 28130
rect 18018 28100 18340 28130
rect 18018 28096 18030 28100
rect 17830 28090 18030 28096
rect 18328 28096 18340 28100
rect 18516 28096 18528 28130
rect 18328 28090 18528 28096
rect 18560 28100 18640 28120
rect 17792 28052 17800 28086
rect 17790 28040 17800 28052
rect 17720 28020 17800 28040
rect 17830 28042 18030 28048
rect 17830 28008 17842 28042
rect 18018 28040 18030 28042
rect 18328 28042 18528 28048
rect 18328 28040 18340 28042
rect 18018 28030 18340 28040
rect 18018 28010 18150 28030
rect 18018 28008 18030 28010
rect 17830 28002 18030 28008
rect 18140 27970 18150 28010
rect 18210 28010 18340 28030
rect 18210 27970 18220 28010
rect 18328 28008 18340 28010
rect 18516 28008 18528 28042
rect 18560 28040 18570 28100
rect 18630 28040 18640 28100
rect 18560 28020 18640 28040
rect 18328 28002 18528 28008
rect 18140 27960 18220 27970
rect 17610 27360 17680 27940
rect 18690 27940 18700 28180
rect 18740 27940 18760 28180
rect 18690 27530 18760 27940
rect 18750 27400 18760 27440
rect 18690 27360 18760 27390
rect 18790 27360 18820 29920
rect 19140 29590 19200 29600
rect 18940 29530 19140 29550
rect 22310 29590 22370 29600
rect 18940 29520 19200 29530
rect 19320 29530 19380 29540
rect 18850 29140 18910 29150
rect 18850 29070 18910 29080
rect 18880 27360 18910 29070
rect 18940 27360 18970 29520
rect 19060 29470 19320 29490
rect 22130 29530 22190 29540
rect 19060 29460 19380 29470
rect 21950 29470 22010 29480
rect 19060 27360 19090 29460
rect 21770 29410 21830 29420
rect 22370 29530 22570 29550
rect 22310 29520 22570 29530
rect 22190 29470 22450 29490
rect 22130 29460 22450 29470
rect 22010 29410 22330 29430
rect 21950 29400 22330 29410
rect 21830 29350 22210 29370
rect 21770 29340 22210 29350
rect 19180 27360 19210 29070
rect 19300 27360 19330 29070
rect 19420 27360 19450 29070
rect 19540 27360 19570 29070
rect 19660 27360 19690 29070
rect 21820 27360 21850 29070
rect 21940 27360 21970 29070
rect 22060 27360 22090 29070
rect 22180 27360 22210 29340
rect 22300 27360 22330 29400
rect 22420 27360 22450 29460
rect 22540 27360 22570 29520
rect 23670 29140 23750 29150
rect 22600 29080 22610 29140
rect 22670 29080 22680 29140
rect 22600 29070 22680 29080
rect 23670 29080 23680 29140
rect 23740 29080 23750 29140
rect 23670 29070 23750 29080
rect 22600 28960 22670 29070
rect 22600 28950 23750 28960
rect 22600 28890 22610 28950
rect 22670 28900 23750 28950
rect 22670 28890 22680 28900
rect 22600 28880 22680 28890
rect 22600 28500 22670 28880
rect 22600 28260 22620 28500
rect 22660 28260 22670 28500
rect 23680 28500 23750 28900
rect 23130 28480 23210 28490
rect 22820 28440 23020 28446
rect 23130 28440 23140 28480
rect 22710 28410 22790 28430
rect 22710 28350 22720 28410
rect 22780 28396 22790 28410
rect 22820 28406 22832 28440
rect 23008 28420 23140 28440
rect 23200 28440 23210 28480
rect 23318 28440 23518 28446
rect 23200 28420 23330 28440
rect 23008 28410 23330 28420
rect 23008 28406 23020 28410
rect 22820 28400 23020 28406
rect 23318 28406 23330 28410
rect 23506 28406 23518 28440
rect 23318 28400 23518 28406
rect 23550 28410 23630 28430
rect 22782 28362 22790 28396
rect 22780 28350 22790 28362
rect 22710 28330 22790 28350
rect 22820 28352 23020 28358
rect 22820 28318 22832 28352
rect 23008 28350 23020 28352
rect 23318 28352 23518 28358
rect 23318 28350 23330 28352
rect 23008 28320 23330 28350
rect 23008 28318 23020 28320
rect 22820 28312 23020 28318
rect 22600 28200 22670 28260
rect 22600 27940 22620 28200
rect 22660 27940 22670 28200
rect 23130 28310 23210 28320
rect 23318 28318 23330 28320
rect 23506 28318 23518 28352
rect 23550 28350 23560 28410
rect 23620 28350 23630 28410
rect 23550 28330 23630 28350
rect 23318 28312 23518 28318
rect 23130 28250 23140 28310
rect 23200 28250 23210 28310
rect 23130 28200 23210 28250
rect 23130 28140 23140 28200
rect 23200 28140 23210 28200
rect 22820 28130 23020 28136
rect 23130 28130 23210 28140
rect 23680 28260 23690 28500
rect 23730 28260 23750 28500
rect 23680 28180 23750 28260
rect 23318 28130 23518 28136
rect 22710 28100 22790 28120
rect 22710 28040 22720 28100
rect 22780 28086 22790 28100
rect 22820 28096 22832 28130
rect 23008 28100 23330 28130
rect 23008 28096 23020 28100
rect 22820 28090 23020 28096
rect 23318 28096 23330 28100
rect 23506 28096 23518 28130
rect 23318 28090 23518 28096
rect 23550 28100 23630 28120
rect 22782 28052 22790 28086
rect 22780 28040 22790 28052
rect 22710 28020 22790 28040
rect 22820 28042 23020 28048
rect 22820 28008 22832 28042
rect 23008 28040 23020 28042
rect 23318 28042 23518 28048
rect 23318 28040 23330 28042
rect 23008 28030 23330 28040
rect 23008 28010 23140 28030
rect 23008 28008 23020 28010
rect 22820 28002 23020 28008
rect 23130 27970 23140 28010
rect 23200 28010 23330 28030
rect 23200 27970 23210 28010
rect 23318 28008 23330 28010
rect 23506 28008 23518 28042
rect 23550 28040 23560 28100
rect 23620 28040 23630 28100
rect 23550 28020 23630 28040
rect 23318 28002 23518 28008
rect 23130 27960 23210 27970
rect 22600 27360 22670 27940
rect 23680 27940 23690 28180
rect 23730 27940 23750 28180
rect 23680 27530 23750 27940
rect 23740 27400 23750 27440
rect 23680 27360 23750 27390
rect 23780 27360 23810 29920
rect 24130 29590 24190 29600
rect 23930 29530 24130 29550
rect 27300 29590 27360 29600
rect 23930 29520 24190 29530
rect 24310 29530 24370 29540
rect 23840 29140 23900 29150
rect 23840 29070 23900 29080
rect 23870 27360 23900 29070
rect 23930 27360 23960 29520
rect 24050 29470 24310 29490
rect 27120 29530 27180 29540
rect 24050 29460 24370 29470
rect 24490 29470 24550 29480
rect 24050 27360 24080 29460
rect 24170 29410 24490 29430
rect 26940 29470 27000 29480
rect 24170 29400 24550 29410
rect 24670 29410 24730 29420
rect 24170 27360 24200 29400
rect 24290 29350 24670 29370
rect 24290 29340 24730 29350
rect 26760 29410 26820 29420
rect 27360 29530 27560 29550
rect 27300 29520 27560 29530
rect 27180 29470 27440 29490
rect 27120 29460 27440 29470
rect 27000 29410 27320 29430
rect 26940 29400 27320 29410
rect 26820 29350 27200 29370
rect 26760 29340 27200 29350
rect 24290 27360 24320 29340
rect 24410 27360 24440 29070
rect 24530 27360 24560 29070
rect 24650 27360 24680 29070
rect 26810 27360 26840 29070
rect 26930 27360 26960 29070
rect 27050 27360 27080 29070
rect 27170 27360 27200 29340
rect 27290 27360 27320 29400
rect 27410 27360 27440 29460
rect 27530 27360 27560 29520
rect 28660 29140 28740 29150
rect 27590 29080 27600 29140
rect 27660 29080 27670 29140
rect 27590 29070 27670 29080
rect 28660 29080 28670 29140
rect 28730 29080 28740 29140
rect 28660 29070 28740 29080
rect 27590 28960 27660 29070
rect 27590 28950 28740 28960
rect 27590 28890 27600 28950
rect 27660 28900 28740 28950
rect 27660 28890 27670 28900
rect 27590 28880 27670 28890
rect 27590 28500 27660 28880
rect 27590 28260 27610 28500
rect 27650 28260 27660 28500
rect 28670 28500 28740 28900
rect 28120 28480 28200 28490
rect 27810 28440 28010 28446
rect 28120 28440 28130 28480
rect 27700 28410 27780 28430
rect 27700 28350 27710 28410
rect 27770 28396 27780 28410
rect 27810 28406 27822 28440
rect 27998 28420 28130 28440
rect 28190 28440 28200 28480
rect 28308 28440 28508 28446
rect 28190 28420 28320 28440
rect 27998 28410 28320 28420
rect 27998 28406 28010 28410
rect 27810 28400 28010 28406
rect 28308 28406 28320 28410
rect 28496 28406 28508 28440
rect 28308 28400 28508 28406
rect 28540 28410 28620 28430
rect 27772 28362 27780 28396
rect 27770 28350 27780 28362
rect 27700 28330 27780 28350
rect 27810 28352 28010 28358
rect 27810 28318 27822 28352
rect 27998 28350 28010 28352
rect 28308 28352 28508 28358
rect 28308 28350 28320 28352
rect 27998 28320 28320 28350
rect 27998 28318 28010 28320
rect 27810 28312 28010 28318
rect 27590 28200 27660 28260
rect 27590 27940 27610 28200
rect 27650 27940 27660 28200
rect 28120 28310 28200 28320
rect 28308 28318 28320 28320
rect 28496 28318 28508 28352
rect 28540 28350 28550 28410
rect 28610 28350 28620 28410
rect 28540 28330 28620 28350
rect 28308 28312 28508 28318
rect 28120 28250 28130 28310
rect 28190 28250 28200 28310
rect 28120 28200 28200 28250
rect 28120 28140 28130 28200
rect 28190 28140 28200 28200
rect 27810 28130 28010 28136
rect 28120 28130 28200 28140
rect 28670 28260 28680 28500
rect 28720 28260 28740 28500
rect 28670 28180 28740 28260
rect 28308 28130 28508 28136
rect 27700 28100 27780 28120
rect 27700 28040 27710 28100
rect 27770 28086 27780 28100
rect 27810 28096 27822 28130
rect 27998 28100 28320 28130
rect 27998 28096 28010 28100
rect 27810 28090 28010 28096
rect 28308 28096 28320 28100
rect 28496 28096 28508 28130
rect 28308 28090 28508 28096
rect 28540 28100 28620 28120
rect 27772 28052 27780 28086
rect 27770 28040 27780 28052
rect 27700 28020 27780 28040
rect 27810 28042 28010 28048
rect 27810 28008 27822 28042
rect 27998 28040 28010 28042
rect 28308 28042 28508 28048
rect 28308 28040 28320 28042
rect 27998 28030 28320 28040
rect 27998 28010 28130 28030
rect 27998 28008 28010 28010
rect 27810 28002 28010 28008
rect 28120 27970 28130 28010
rect 28190 28010 28320 28030
rect 28190 27970 28200 28010
rect 28308 28008 28320 28010
rect 28496 28008 28508 28042
rect 28540 28040 28550 28100
rect 28610 28040 28620 28100
rect 28540 28020 28620 28040
rect 28308 28002 28508 28008
rect 28120 27960 28200 27970
rect 27590 27360 27660 27940
rect 28670 27940 28680 28180
rect 28720 27940 28740 28180
rect 28670 27530 28740 27940
rect 28730 27400 28740 27440
rect 28670 27360 28740 27390
rect 28770 27360 28800 29920
rect 29120 29590 29180 29600
rect 28920 29530 29120 29550
rect 32290 29590 32350 29600
rect 28920 29520 29180 29530
rect 29300 29530 29360 29540
rect 28830 29140 28890 29150
rect 28830 29070 28890 29080
rect 28860 27360 28890 29070
rect 28920 27360 28950 29520
rect 29040 29470 29300 29490
rect 32110 29530 32170 29540
rect 29040 29460 29360 29470
rect 29480 29470 29540 29480
rect 29040 27360 29070 29460
rect 29160 29410 29480 29430
rect 31930 29470 31990 29480
rect 29160 29400 29540 29410
rect 29660 29410 29720 29420
rect 29160 27360 29190 29400
rect 29280 29350 29660 29370
rect 31750 29410 31810 29420
rect 29280 29340 29720 29350
rect 31570 29350 31630 29360
rect 29280 27360 29310 29340
rect 31390 29290 31450 29300
rect 32350 29530 32550 29550
rect 32290 29520 32550 29530
rect 32170 29470 32430 29490
rect 32110 29460 32430 29470
rect 31990 29410 32310 29430
rect 31930 29400 32310 29410
rect 31810 29350 32190 29370
rect 31750 29340 32190 29350
rect 31630 29290 32070 29310
rect 31570 29280 32070 29290
rect 31450 29230 31950 29250
rect 31390 29220 31950 29230
rect 29400 27360 29430 29070
rect 29520 27360 29550 29070
rect 29640 27360 29670 29070
rect 31800 27360 31830 29070
rect 31920 27360 31950 29220
rect 32040 27360 32070 29280
rect 32160 27360 32190 29340
rect 32280 27360 32310 29400
rect 32400 27360 32430 29460
rect 32520 27360 32550 29520
rect 33650 29140 33730 29150
rect 32580 29080 32590 29140
rect 32650 29080 32660 29140
rect 32580 29070 32660 29080
rect 33650 29080 33660 29140
rect 33720 29080 33730 29140
rect 33650 29070 33730 29080
rect 32580 28960 32650 29070
rect 32580 28950 33730 28960
rect 32580 28890 32590 28950
rect 32650 28900 33730 28950
rect 32650 28890 32660 28900
rect 32580 28880 32660 28890
rect 32580 28500 32650 28880
rect 32580 28260 32600 28500
rect 32640 28260 32650 28500
rect 33660 28500 33730 28900
rect 33110 28480 33190 28490
rect 32800 28440 33000 28446
rect 33110 28440 33120 28480
rect 32690 28410 32770 28430
rect 32690 28350 32700 28410
rect 32760 28396 32770 28410
rect 32800 28406 32812 28440
rect 32988 28420 33120 28440
rect 33180 28440 33190 28480
rect 33298 28440 33498 28446
rect 33180 28420 33310 28440
rect 32988 28410 33310 28420
rect 32988 28406 33000 28410
rect 32800 28400 33000 28406
rect 33298 28406 33310 28410
rect 33486 28406 33498 28440
rect 33298 28400 33498 28406
rect 33530 28410 33610 28430
rect 32762 28362 32770 28396
rect 32760 28350 32770 28362
rect 32690 28330 32770 28350
rect 32800 28352 33000 28358
rect 32800 28318 32812 28352
rect 32988 28350 33000 28352
rect 33298 28352 33498 28358
rect 33298 28350 33310 28352
rect 32988 28320 33310 28350
rect 32988 28318 33000 28320
rect 32800 28312 33000 28318
rect 32580 28200 32650 28260
rect 32580 27940 32600 28200
rect 32640 27940 32650 28200
rect 33110 28310 33190 28320
rect 33298 28318 33310 28320
rect 33486 28318 33498 28352
rect 33530 28350 33540 28410
rect 33600 28350 33610 28410
rect 33530 28330 33610 28350
rect 33298 28312 33498 28318
rect 33110 28250 33120 28310
rect 33180 28250 33190 28310
rect 33110 28200 33190 28250
rect 33110 28140 33120 28200
rect 33180 28140 33190 28200
rect 32800 28130 33000 28136
rect 33110 28130 33190 28140
rect 33660 28260 33670 28500
rect 33710 28260 33730 28500
rect 33660 28180 33730 28260
rect 33298 28130 33498 28136
rect 32690 28100 32770 28120
rect 32690 28040 32700 28100
rect 32760 28086 32770 28100
rect 32800 28096 32812 28130
rect 32988 28100 33310 28130
rect 32988 28096 33000 28100
rect 32800 28090 33000 28096
rect 33298 28096 33310 28100
rect 33486 28096 33498 28130
rect 33298 28090 33498 28096
rect 33530 28100 33610 28120
rect 32762 28052 32770 28086
rect 32760 28040 32770 28052
rect 32690 28020 32770 28040
rect 32800 28042 33000 28048
rect 32800 28008 32812 28042
rect 32988 28040 33000 28042
rect 33298 28042 33498 28048
rect 33298 28040 33310 28042
rect 32988 28030 33310 28040
rect 32988 28010 33120 28030
rect 32988 28008 33000 28010
rect 32800 28002 33000 28008
rect 33110 27970 33120 28010
rect 33180 28010 33310 28030
rect 33180 27970 33190 28010
rect 33298 28008 33310 28010
rect 33486 28008 33498 28042
rect 33530 28040 33540 28100
rect 33600 28040 33610 28100
rect 33530 28020 33610 28040
rect 33298 28002 33498 28008
rect 33110 27960 33190 27970
rect 32580 27360 32650 27940
rect 33660 27940 33670 28180
rect 33710 27940 33730 28180
rect 33660 27530 33730 27940
rect 33720 27400 33730 27440
rect 33660 27360 33730 27390
rect 33760 27360 33790 29920
rect 34110 29590 34170 29600
rect 33910 29530 34110 29550
rect 37280 29590 37340 29600
rect 33910 29520 34170 29530
rect 34290 29530 34350 29540
rect 33820 29140 33880 29150
rect 33820 29070 33880 29080
rect 33850 27360 33880 29070
rect 33910 27360 33940 29520
rect 34030 29470 34290 29490
rect 37100 29530 37160 29540
rect 34030 29460 34350 29470
rect 34470 29470 34530 29480
rect 34030 27360 34060 29460
rect 34150 29410 34470 29430
rect 36920 29470 36980 29480
rect 34150 29400 34530 29410
rect 34650 29410 34710 29420
rect 34150 27360 34180 29400
rect 34270 29350 34650 29370
rect 36740 29410 36800 29420
rect 34270 29340 34710 29350
rect 34830 29350 34890 29360
rect 34270 27360 34300 29340
rect 34390 29290 34830 29310
rect 36560 29350 36620 29360
rect 34390 29280 34890 29290
rect 35010 29290 35070 29300
rect 34390 27360 34420 29280
rect 34510 29230 35010 29250
rect 36380 29290 36440 29300
rect 34510 29220 35070 29230
rect 36200 29230 36260 29240
rect 34510 27360 34540 29220
rect 37340 29530 37540 29550
rect 37280 29520 37540 29530
rect 37160 29470 37420 29490
rect 37100 29460 37420 29470
rect 36980 29410 37300 29430
rect 36920 29400 37300 29410
rect 36800 29350 37180 29370
rect 36740 29340 37180 29350
rect 36620 29290 37060 29310
rect 36560 29280 37060 29290
rect 36440 29230 36940 29250
rect 36380 29220 36940 29230
rect 36260 29170 36820 29190
rect 36200 29160 36820 29170
rect 34630 27360 34660 29070
rect 36790 27360 36820 29160
rect 36910 27360 36940 29220
rect 37030 27360 37060 29280
rect 37150 27360 37180 29340
rect 37270 27360 37300 29400
rect 37390 27360 37420 29460
rect 37510 27360 37540 29520
rect 38640 29140 38720 29150
rect 37570 29080 37580 29140
rect 37640 29080 37650 29140
rect 37570 29070 37650 29080
rect 38640 29080 38650 29140
rect 38710 29080 38720 29140
rect 38640 29070 38720 29080
rect 37570 28960 37640 29070
rect 37570 28950 38720 28960
rect 37570 28890 37580 28950
rect 37640 28900 38720 28950
rect 37640 28890 37650 28900
rect 37570 28880 37650 28890
rect 37570 28500 37640 28880
rect 37570 28260 37590 28500
rect 37630 28260 37640 28500
rect 38650 28500 38720 28900
rect 38100 28480 38180 28490
rect 37790 28440 37990 28446
rect 38100 28440 38110 28480
rect 37680 28410 37760 28430
rect 37680 28350 37690 28410
rect 37750 28396 37760 28410
rect 37790 28406 37802 28440
rect 37978 28420 38110 28440
rect 38170 28440 38180 28480
rect 38288 28440 38488 28446
rect 38170 28420 38300 28440
rect 37978 28410 38300 28420
rect 37978 28406 37990 28410
rect 37790 28400 37990 28406
rect 38288 28406 38300 28410
rect 38476 28406 38488 28440
rect 38288 28400 38488 28406
rect 38520 28410 38600 28430
rect 37752 28362 37760 28396
rect 37750 28350 37760 28362
rect 37680 28330 37760 28350
rect 37790 28352 37990 28358
rect 37790 28318 37802 28352
rect 37978 28350 37990 28352
rect 38288 28352 38488 28358
rect 38288 28350 38300 28352
rect 37978 28320 38300 28350
rect 37978 28318 37990 28320
rect 37790 28312 37990 28318
rect 37570 28200 37640 28260
rect 37570 27940 37590 28200
rect 37630 27940 37640 28200
rect 38100 28310 38180 28320
rect 38288 28318 38300 28320
rect 38476 28318 38488 28352
rect 38520 28350 38530 28410
rect 38590 28350 38600 28410
rect 38520 28330 38600 28350
rect 38288 28312 38488 28318
rect 38100 28250 38110 28310
rect 38170 28250 38180 28310
rect 38100 28200 38180 28250
rect 38100 28140 38110 28200
rect 38170 28140 38180 28200
rect 37790 28130 37990 28136
rect 38100 28130 38180 28140
rect 38650 28260 38660 28500
rect 38700 28260 38720 28500
rect 38650 28180 38720 28260
rect 38288 28130 38488 28136
rect 37680 28100 37760 28120
rect 37680 28040 37690 28100
rect 37750 28086 37760 28100
rect 37790 28096 37802 28130
rect 37978 28100 38300 28130
rect 37978 28096 37990 28100
rect 37790 28090 37990 28096
rect 38288 28096 38300 28100
rect 38476 28096 38488 28130
rect 38288 28090 38488 28096
rect 38520 28100 38600 28120
rect 37752 28052 37760 28086
rect 37750 28040 37760 28052
rect 37680 28020 37760 28040
rect 37790 28042 37990 28048
rect 37790 28008 37802 28042
rect 37978 28040 37990 28042
rect 38288 28042 38488 28048
rect 38288 28040 38300 28042
rect 37978 28030 38300 28040
rect 37978 28010 38110 28030
rect 37978 28008 37990 28010
rect 37790 28002 37990 28008
rect 38100 27970 38110 28010
rect 38170 28010 38300 28030
rect 38170 27970 38180 28010
rect 38288 28008 38300 28010
rect 38476 28008 38488 28042
rect 38520 28040 38530 28100
rect 38590 28040 38600 28100
rect 38520 28020 38600 28040
rect 38288 28002 38488 28008
rect 38100 27960 38180 27970
rect 37570 27360 37640 27940
rect 38650 27940 38660 28180
rect 38700 27940 38720 28180
rect 38650 27530 38720 27940
rect 38710 27400 38720 27440
rect 38650 27360 38720 27390
rect 38750 27360 38780 29920
rect 39100 29590 39160 29600
rect 38900 29530 39100 29550
rect 42270 29590 42330 29600
rect 38900 29520 39160 29530
rect 39280 29530 39340 29540
rect 38810 29140 38870 29150
rect 38810 29070 38870 29080
rect 38840 27360 38870 29070
rect 38900 27360 38930 29520
rect 39020 29470 39280 29490
rect 42090 29530 42150 29540
rect 39020 29460 39340 29470
rect 39460 29470 39520 29480
rect 39020 27360 39050 29460
rect 39140 29410 39460 29430
rect 41910 29470 41970 29480
rect 39140 29400 39520 29410
rect 39640 29410 39700 29420
rect 39140 27360 39170 29400
rect 39260 29350 39640 29370
rect 41730 29410 41790 29420
rect 39260 29340 39700 29350
rect 39820 29350 39880 29360
rect 39260 27360 39290 29340
rect 39380 29290 39820 29310
rect 41550 29350 41610 29360
rect 39380 29280 39880 29290
rect 40000 29290 40060 29300
rect 39380 27360 39410 29280
rect 39500 29230 40000 29250
rect 41370 29290 41430 29300
rect 39500 29220 40060 29230
rect 40180 29230 40240 29240
rect 39500 27360 39530 29220
rect 39620 29170 40180 29190
rect 39620 29160 40240 29170
rect 41190 29230 41250 29240
rect 42330 29530 42530 29550
rect 42270 29520 42530 29530
rect 42150 29470 42410 29490
rect 42090 29460 42410 29470
rect 41970 29410 42290 29430
rect 41910 29400 42290 29410
rect 41790 29350 42170 29370
rect 41730 29340 42170 29350
rect 41610 29290 42050 29310
rect 41550 29280 42050 29290
rect 41430 29230 41930 29250
rect 41370 29220 41930 29230
rect 41250 29170 41810 29190
rect 41190 29160 41810 29170
rect 39620 27360 39650 29160
rect 41780 27360 41810 29160
rect 41900 27360 41930 29220
rect 42020 27360 42050 29280
rect 42140 27360 42170 29340
rect 42260 27360 42290 29400
rect 42380 27360 42410 29460
rect 42500 27360 42530 29520
rect 43630 29140 43710 29150
rect 42560 29080 42570 29140
rect 42630 29080 42640 29140
rect 42560 29070 42640 29080
rect 43630 29080 43640 29140
rect 43700 29080 43710 29140
rect 43630 29070 43710 29080
rect 42560 28960 42630 29070
rect 42560 28950 43710 28960
rect 42560 28890 42570 28950
rect 42630 28900 43710 28950
rect 42630 28890 42640 28900
rect 42560 28880 42640 28890
rect 42560 28500 42630 28880
rect 42560 28260 42580 28500
rect 42620 28260 42630 28500
rect 43640 28500 43710 28900
rect 43090 28480 43170 28490
rect 42780 28440 42980 28446
rect 43090 28440 43100 28480
rect 42670 28410 42750 28430
rect 42670 28350 42680 28410
rect 42740 28396 42750 28410
rect 42780 28406 42792 28440
rect 42968 28420 43100 28440
rect 43160 28440 43170 28480
rect 43278 28440 43478 28446
rect 43160 28420 43290 28440
rect 42968 28410 43290 28420
rect 42968 28406 42980 28410
rect 42780 28400 42980 28406
rect 43278 28406 43290 28410
rect 43466 28406 43478 28440
rect 43278 28400 43478 28406
rect 43510 28410 43590 28430
rect 42742 28362 42750 28396
rect 42740 28350 42750 28362
rect 42670 28330 42750 28350
rect 42780 28352 42980 28358
rect 42780 28318 42792 28352
rect 42968 28350 42980 28352
rect 43278 28352 43478 28358
rect 43278 28350 43290 28352
rect 42968 28320 43290 28350
rect 42968 28318 42980 28320
rect 42780 28312 42980 28318
rect 42560 28200 42630 28260
rect 42560 27940 42580 28200
rect 42620 27940 42630 28200
rect 43090 28310 43170 28320
rect 43278 28318 43290 28320
rect 43466 28318 43478 28352
rect 43510 28350 43520 28410
rect 43580 28350 43590 28410
rect 43510 28330 43590 28350
rect 43278 28312 43478 28318
rect 43090 28250 43100 28310
rect 43160 28250 43170 28310
rect 43090 28200 43170 28250
rect 43090 28140 43100 28200
rect 43160 28140 43170 28200
rect 42780 28130 42980 28136
rect 43090 28130 43170 28140
rect 43640 28260 43650 28500
rect 43690 28260 43710 28500
rect 43640 28180 43710 28260
rect 43278 28130 43478 28136
rect 42670 28100 42750 28120
rect 42670 28040 42680 28100
rect 42740 28086 42750 28100
rect 42780 28096 42792 28130
rect 42968 28100 43290 28130
rect 42968 28096 42980 28100
rect 42780 28090 42980 28096
rect 43278 28096 43290 28100
rect 43466 28096 43478 28130
rect 43278 28090 43478 28096
rect 43510 28100 43590 28120
rect 42742 28052 42750 28086
rect 42740 28040 42750 28052
rect 42670 28020 42750 28040
rect 42780 28042 42980 28048
rect 42780 28008 42792 28042
rect 42968 28040 42980 28042
rect 43278 28042 43478 28048
rect 43278 28040 43290 28042
rect 42968 28030 43290 28040
rect 42968 28010 43100 28030
rect 42968 28008 42980 28010
rect 42780 28002 42980 28008
rect 43090 27970 43100 28010
rect 43160 28010 43290 28030
rect 43160 27970 43170 28010
rect 43278 28008 43290 28010
rect 43466 28008 43478 28042
rect 43510 28040 43520 28100
rect 43580 28040 43590 28100
rect 43510 28020 43590 28040
rect 43278 28002 43478 28008
rect 43090 27960 43170 27970
rect 42560 27360 42630 27940
rect 43640 27940 43650 28180
rect 43690 27940 43710 28180
rect 43640 27530 43710 27940
rect 43700 27400 43710 27440
rect 43640 27360 43710 27390
rect 43740 27360 43770 29920
rect 44090 29590 44150 29600
rect 43890 29530 44090 29550
rect 47260 29590 47320 29600
rect 43890 29520 44150 29530
rect 44270 29530 44330 29540
rect 43800 29140 43860 29150
rect 43800 29070 43860 29080
rect 43830 27360 43860 29070
rect 43890 27360 43920 29520
rect 44010 29470 44270 29490
rect 47080 29530 47140 29540
rect 44010 29460 44330 29470
rect 44450 29470 44510 29480
rect 44010 27360 44040 29460
rect 44130 29410 44450 29430
rect 46900 29470 46960 29480
rect 44130 29400 44510 29410
rect 44630 29410 44690 29420
rect 44130 27360 44160 29400
rect 44250 29350 44630 29370
rect 46720 29410 46780 29420
rect 44250 29340 44690 29350
rect 44810 29350 44870 29360
rect 44250 27360 44280 29340
rect 44370 29290 44810 29310
rect 46540 29350 46600 29360
rect 44370 29280 44870 29290
rect 44990 29290 45050 29300
rect 44370 27330 44400 29280
rect 44490 29230 44990 29250
rect 46360 29290 46420 29300
rect 44490 29220 45050 29230
rect 45170 29230 45230 29240
rect 44490 27360 44520 29220
rect 44610 29170 45170 29190
rect 47320 29530 47520 29550
rect 47260 29520 47520 29530
rect 47140 29470 47400 29490
rect 47080 29460 47400 29470
rect 46960 29410 47280 29430
rect 46900 29400 47280 29410
rect 46780 29350 47160 29370
rect 46720 29340 47160 29350
rect 46600 29290 47040 29310
rect 46540 29280 47040 29290
rect 46420 29230 46920 29250
rect 46360 29220 46920 29230
rect 44610 29160 45230 29170
rect 44610 27360 44640 29160
rect 46770 27360 46800 29070
rect 46890 27360 46920 29220
rect 47010 27360 47040 29280
rect 47130 27360 47160 29340
rect 47250 27360 47280 29400
rect 47370 27360 47400 29460
rect 47490 27360 47520 29520
rect 48620 29140 48700 29150
rect 47550 29080 47560 29140
rect 47620 29080 47630 29140
rect 47550 29070 47630 29080
rect 48620 29080 48630 29140
rect 48690 29080 48700 29140
rect 48620 29070 48700 29080
rect 47550 28960 47620 29070
rect 47550 28950 48700 28960
rect 47550 28890 47560 28950
rect 47620 28900 48700 28950
rect 47620 28890 47630 28900
rect 47550 28880 47630 28890
rect 47550 28500 47620 28880
rect 47550 28260 47570 28500
rect 47610 28260 47620 28500
rect 48630 28500 48700 28900
rect 48080 28480 48160 28490
rect 47770 28440 47970 28446
rect 48080 28440 48090 28480
rect 47660 28410 47740 28430
rect 47660 28350 47670 28410
rect 47730 28396 47740 28410
rect 47770 28406 47782 28440
rect 47958 28420 48090 28440
rect 48150 28440 48160 28480
rect 48268 28440 48468 28446
rect 48150 28420 48280 28440
rect 47958 28410 48280 28420
rect 47958 28406 47970 28410
rect 47770 28400 47970 28406
rect 48268 28406 48280 28410
rect 48456 28406 48468 28440
rect 48268 28400 48468 28406
rect 48500 28410 48580 28430
rect 47732 28362 47740 28396
rect 47730 28350 47740 28362
rect 47660 28330 47740 28350
rect 47770 28352 47970 28358
rect 47770 28318 47782 28352
rect 47958 28350 47970 28352
rect 48268 28352 48468 28358
rect 48268 28350 48280 28352
rect 47958 28320 48280 28350
rect 47958 28318 47970 28320
rect 47770 28312 47970 28318
rect 47550 28200 47620 28260
rect 47550 27940 47570 28200
rect 47610 27940 47620 28200
rect 48080 28310 48160 28320
rect 48268 28318 48280 28320
rect 48456 28318 48468 28352
rect 48500 28350 48510 28410
rect 48570 28350 48580 28410
rect 48500 28330 48580 28350
rect 48268 28312 48468 28318
rect 48080 28250 48090 28310
rect 48150 28250 48160 28310
rect 48080 28200 48160 28250
rect 48080 28140 48090 28200
rect 48150 28140 48160 28200
rect 47770 28130 47970 28136
rect 48080 28130 48160 28140
rect 48630 28260 48640 28500
rect 48680 28260 48700 28500
rect 48630 28180 48700 28260
rect 48268 28130 48468 28136
rect 47660 28100 47740 28120
rect 47660 28040 47670 28100
rect 47730 28086 47740 28100
rect 47770 28096 47782 28130
rect 47958 28100 48280 28130
rect 47958 28096 47970 28100
rect 47770 28090 47970 28096
rect 48268 28096 48280 28100
rect 48456 28096 48468 28130
rect 48268 28090 48468 28096
rect 48500 28100 48580 28120
rect 47732 28052 47740 28086
rect 47730 28040 47740 28052
rect 47660 28020 47740 28040
rect 47770 28042 47970 28048
rect 47770 28008 47782 28042
rect 47958 28040 47970 28042
rect 48268 28042 48468 28048
rect 48268 28040 48280 28042
rect 47958 28030 48280 28040
rect 47958 28010 48090 28030
rect 47958 28008 47970 28010
rect 47770 28002 47970 28008
rect 48080 27970 48090 28010
rect 48150 28010 48280 28030
rect 48150 27970 48160 28010
rect 48268 28008 48280 28010
rect 48456 28008 48468 28042
rect 48500 28040 48510 28100
rect 48570 28040 48580 28100
rect 48500 28020 48580 28040
rect 48268 28002 48468 28008
rect 48080 27960 48160 27970
rect 47550 27360 47620 27940
rect 48630 27940 48640 28180
rect 48680 27940 48700 28180
rect 48630 27530 48700 27940
rect 48690 27400 48700 27440
rect 48630 27360 48700 27390
rect 48730 27360 48760 29920
rect 49080 29590 49140 29600
rect 48880 29530 49080 29550
rect 52250 29590 52310 29600
rect 48880 29520 49140 29530
rect 49260 29530 49320 29540
rect 48790 29140 48850 29150
rect 48790 29070 48850 29080
rect 48820 27360 48850 29070
rect 48880 27360 48910 29520
rect 49000 29470 49260 29490
rect 52070 29530 52130 29540
rect 49000 29460 49320 29470
rect 49440 29470 49500 29480
rect 49000 27360 49030 29460
rect 49120 29410 49440 29430
rect 51890 29470 51950 29480
rect 49120 29400 49500 29410
rect 49620 29410 49680 29420
rect 49120 27360 49150 29400
rect 49240 29350 49620 29370
rect 51710 29410 51770 29420
rect 49240 29340 49680 29350
rect 49800 29350 49860 29360
rect 49240 27360 49270 29340
rect 49360 29290 49800 29310
rect 52310 29530 52510 29550
rect 52250 29520 52510 29530
rect 52130 29470 52390 29490
rect 52070 29460 52390 29470
rect 51950 29410 52270 29430
rect 51890 29400 52270 29410
rect 51770 29350 52150 29370
rect 51710 29340 52150 29350
rect 49360 29280 49860 29290
rect 49980 29290 50040 29300
rect 49360 27360 49390 29280
rect 49480 29230 49980 29250
rect 49480 29220 50040 29230
rect 49480 27360 49510 29220
rect 49600 27360 49630 29070
rect 51760 27360 51790 29070
rect 51880 27360 51910 29070
rect 52000 27360 52030 29070
rect 52120 27360 52150 29340
rect 52240 27360 52270 29400
rect 52360 27360 52390 29460
rect 52480 27360 52510 29520
rect 53610 29140 53690 29150
rect 52540 29080 52550 29140
rect 52610 29080 52620 29140
rect 52540 29070 52620 29080
rect 53610 29080 53620 29140
rect 53680 29080 53690 29140
rect 53610 29070 53690 29080
rect 52540 28960 52610 29070
rect 52540 28950 53690 28960
rect 52540 28890 52550 28950
rect 52610 28900 53690 28950
rect 52610 28890 52620 28900
rect 52540 28880 52620 28890
rect 52540 28500 52610 28880
rect 52540 28260 52560 28500
rect 52600 28260 52610 28500
rect 53620 28500 53690 28900
rect 53070 28480 53150 28490
rect 52760 28440 52960 28446
rect 53070 28440 53080 28480
rect 52650 28410 52730 28430
rect 52650 28350 52660 28410
rect 52720 28396 52730 28410
rect 52760 28406 52772 28440
rect 52948 28420 53080 28440
rect 53140 28440 53150 28480
rect 53258 28440 53458 28446
rect 53140 28420 53270 28440
rect 52948 28410 53270 28420
rect 52948 28406 52960 28410
rect 52760 28400 52960 28406
rect 53258 28406 53270 28410
rect 53446 28406 53458 28440
rect 53258 28400 53458 28406
rect 53490 28410 53570 28430
rect 52722 28362 52730 28396
rect 52720 28350 52730 28362
rect 52650 28330 52730 28350
rect 52760 28352 52960 28358
rect 52760 28318 52772 28352
rect 52948 28350 52960 28352
rect 53258 28352 53458 28358
rect 53258 28350 53270 28352
rect 52948 28320 53270 28350
rect 52948 28318 52960 28320
rect 52760 28312 52960 28318
rect 52540 28200 52610 28260
rect 52540 27940 52560 28200
rect 52600 27940 52610 28200
rect 53070 28310 53150 28320
rect 53258 28318 53270 28320
rect 53446 28318 53458 28352
rect 53490 28350 53500 28410
rect 53560 28350 53570 28410
rect 53490 28330 53570 28350
rect 53258 28312 53458 28318
rect 53070 28250 53080 28310
rect 53140 28250 53150 28310
rect 53070 28200 53150 28250
rect 53070 28140 53080 28200
rect 53140 28140 53150 28200
rect 52760 28130 52960 28136
rect 53070 28130 53150 28140
rect 53620 28260 53630 28500
rect 53670 28260 53690 28500
rect 53620 28180 53690 28260
rect 53258 28130 53458 28136
rect 52650 28100 52730 28120
rect 52650 28040 52660 28100
rect 52720 28086 52730 28100
rect 52760 28096 52772 28130
rect 52948 28100 53270 28130
rect 52948 28096 52960 28100
rect 52760 28090 52960 28096
rect 53258 28096 53270 28100
rect 53446 28096 53458 28130
rect 53258 28090 53458 28096
rect 53490 28100 53570 28120
rect 52722 28052 52730 28086
rect 52720 28040 52730 28052
rect 52650 28020 52730 28040
rect 52760 28042 52960 28048
rect 52760 28008 52772 28042
rect 52948 28040 52960 28042
rect 53258 28042 53458 28048
rect 53258 28040 53270 28042
rect 52948 28030 53270 28040
rect 52948 28010 53080 28030
rect 52948 28008 52960 28010
rect 52760 28002 52960 28008
rect 53070 27970 53080 28010
rect 53140 28010 53270 28030
rect 53140 27970 53150 28010
rect 53258 28008 53270 28010
rect 53446 28008 53458 28042
rect 53490 28040 53500 28100
rect 53560 28040 53570 28100
rect 53490 28020 53570 28040
rect 53258 28002 53458 28008
rect 53070 27960 53150 27970
rect 52540 27360 52610 27940
rect 53620 27940 53630 28180
rect 53670 27940 53690 28180
rect 53620 27530 53690 27940
rect 53680 27400 53690 27440
rect 53620 27360 53690 27390
rect 53720 27360 53750 29920
rect 54070 29590 54130 29600
rect 53870 29530 54070 29550
rect 57240 29590 57300 29600
rect 53870 29520 54130 29530
rect 54250 29530 54310 29540
rect 53780 29140 53840 29150
rect 53780 29070 53840 29080
rect 53810 27360 53840 29070
rect 53870 27360 53900 29520
rect 53990 29470 54250 29490
rect 57060 29530 57120 29540
rect 53990 29460 54310 29470
rect 54430 29470 54490 29480
rect 53990 27360 54020 29460
rect 54110 29410 54430 29430
rect 56880 29470 56940 29480
rect 54110 29400 54490 29410
rect 54610 29410 54670 29420
rect 54110 27360 54140 29400
rect 54230 29350 54610 29370
rect 54230 29340 54670 29350
rect 56700 29410 56760 29420
rect 57300 29530 57500 29550
rect 57240 29520 57500 29530
rect 57120 29470 57380 29490
rect 57060 29460 57380 29470
rect 56940 29410 57260 29430
rect 56880 29400 57260 29410
rect 56760 29350 57140 29370
rect 56700 29340 57140 29350
rect 54230 27360 54260 29340
rect 54350 27360 54380 29070
rect 54470 27360 54500 29070
rect 54590 27360 54620 29070
rect 56750 27360 56780 29070
rect 56870 27360 56900 29070
rect 56990 27360 57020 29070
rect 57110 27360 57140 29340
rect 57230 27360 57260 29400
rect 57350 27360 57380 29460
rect 57470 27360 57500 29520
rect 58600 29140 58680 29150
rect 57530 29080 57540 29140
rect 57600 29080 57610 29140
rect 57530 29070 57610 29080
rect 58600 29080 58610 29140
rect 58670 29080 58680 29140
rect 58600 29070 58680 29080
rect 57530 28960 57600 29070
rect 57530 28950 58680 28960
rect 57530 28890 57540 28950
rect 57600 28900 58680 28950
rect 57600 28890 57610 28900
rect 57530 28880 57610 28890
rect 57530 28500 57600 28880
rect 57530 28260 57550 28500
rect 57590 28260 57600 28500
rect 58610 28500 58680 28900
rect 58060 28480 58140 28490
rect 57750 28440 57950 28446
rect 58060 28440 58070 28480
rect 57640 28410 57720 28430
rect 57640 28350 57650 28410
rect 57710 28396 57720 28410
rect 57750 28406 57762 28440
rect 57938 28420 58070 28440
rect 58130 28440 58140 28480
rect 58248 28440 58448 28446
rect 58130 28420 58260 28440
rect 57938 28410 58260 28420
rect 57938 28406 57950 28410
rect 57750 28400 57950 28406
rect 58248 28406 58260 28410
rect 58436 28406 58448 28440
rect 58248 28400 58448 28406
rect 58480 28410 58560 28430
rect 57712 28362 57720 28396
rect 57710 28350 57720 28362
rect 57640 28330 57720 28350
rect 57750 28352 57950 28358
rect 57750 28318 57762 28352
rect 57938 28350 57950 28352
rect 58248 28352 58448 28358
rect 58248 28350 58260 28352
rect 57938 28320 58260 28350
rect 57938 28318 57950 28320
rect 57750 28312 57950 28318
rect 57530 28200 57600 28260
rect 57530 27940 57550 28200
rect 57590 27940 57600 28200
rect 58060 28310 58140 28320
rect 58248 28318 58260 28320
rect 58436 28318 58448 28352
rect 58480 28350 58490 28410
rect 58550 28350 58560 28410
rect 58480 28330 58560 28350
rect 58248 28312 58448 28318
rect 58060 28250 58070 28310
rect 58130 28250 58140 28310
rect 58060 28200 58140 28250
rect 58060 28140 58070 28200
rect 58130 28140 58140 28200
rect 57750 28130 57950 28136
rect 58060 28130 58140 28140
rect 58610 28260 58620 28500
rect 58660 28260 58680 28500
rect 58610 28180 58680 28260
rect 58248 28130 58448 28136
rect 57640 28100 57720 28120
rect 57640 28040 57650 28100
rect 57710 28086 57720 28100
rect 57750 28096 57762 28130
rect 57938 28100 58260 28130
rect 57938 28096 57950 28100
rect 57750 28090 57950 28096
rect 58248 28096 58260 28100
rect 58436 28096 58448 28130
rect 58248 28090 58448 28096
rect 58480 28100 58560 28120
rect 57712 28052 57720 28086
rect 57710 28040 57720 28052
rect 57640 28020 57720 28040
rect 57750 28042 57950 28048
rect 57750 28008 57762 28042
rect 57938 28040 57950 28042
rect 58248 28042 58448 28048
rect 58248 28040 58260 28042
rect 57938 28030 58260 28040
rect 57938 28010 58070 28030
rect 57938 28008 57950 28010
rect 57750 28002 57950 28008
rect 58060 27970 58070 28010
rect 58130 28010 58260 28030
rect 58130 27970 58140 28010
rect 58248 28008 58260 28010
rect 58436 28008 58448 28042
rect 58480 28040 58490 28100
rect 58550 28040 58560 28100
rect 58480 28020 58560 28040
rect 58248 28002 58448 28008
rect 58060 27960 58140 27970
rect 57530 27360 57600 27940
rect 58610 27940 58620 28180
rect 58660 27940 58680 28180
rect 58610 27530 58680 27940
rect 58670 27400 58680 27440
rect 58610 27360 58680 27390
rect 58710 27360 58740 29920
rect 59060 29590 59120 29600
rect 58860 29530 59060 29550
rect 62230 29590 62290 29600
rect 58860 29520 59120 29530
rect 59240 29530 59300 29540
rect 58770 29140 58830 29150
rect 58770 29070 58830 29080
rect 58800 27360 58830 29070
rect 58860 27360 58890 29520
rect 58980 29470 59240 29490
rect 62050 29530 62110 29540
rect 58980 29460 59300 29470
rect 59420 29470 59480 29480
rect 58980 27360 59010 29460
rect 59100 29410 59420 29430
rect 62290 29530 62490 29550
rect 62230 29520 62490 29530
rect 62110 29470 62370 29490
rect 62050 29460 62370 29470
rect 59100 29400 59480 29410
rect 59600 29410 59660 29420
rect 59100 27360 59130 29400
rect 59220 29350 59600 29370
rect 59220 29340 59660 29350
rect 59220 27360 59250 29340
rect 59340 27360 59370 29070
rect 59460 27360 59490 29070
rect 59580 27360 59610 29070
rect 61740 27360 61770 29070
rect 61860 27360 61890 29070
rect 61980 27360 62010 29070
rect 62100 27360 62130 29070
rect 62220 27360 62250 29070
rect 62340 27360 62370 29460
rect 62460 27360 62490 29520
rect 63590 29140 63670 29150
rect 62520 29080 62530 29140
rect 62590 29080 62600 29140
rect 62520 29070 62600 29080
rect 63590 29080 63600 29140
rect 63660 29080 63670 29140
rect 63590 29070 63670 29080
rect 62520 28960 62590 29070
rect 62520 28950 63670 28960
rect 62520 28890 62530 28950
rect 62590 28900 63670 28950
rect 62590 28890 62600 28900
rect 62520 28880 62600 28890
rect 62520 28500 62590 28880
rect 62520 28260 62540 28500
rect 62580 28260 62590 28500
rect 63600 28500 63670 28900
rect 63050 28480 63130 28490
rect 62740 28440 62940 28446
rect 63050 28440 63060 28480
rect 62630 28410 62710 28430
rect 62630 28350 62640 28410
rect 62700 28396 62710 28410
rect 62740 28406 62752 28440
rect 62928 28420 63060 28440
rect 63120 28440 63130 28480
rect 63238 28440 63438 28446
rect 63120 28420 63250 28440
rect 62928 28410 63250 28420
rect 62928 28406 62940 28410
rect 62740 28400 62940 28406
rect 63238 28406 63250 28410
rect 63426 28406 63438 28440
rect 63238 28400 63438 28406
rect 63470 28410 63550 28430
rect 62702 28362 62710 28396
rect 62700 28350 62710 28362
rect 62630 28330 62710 28350
rect 62740 28352 62940 28358
rect 62740 28318 62752 28352
rect 62928 28350 62940 28352
rect 63238 28352 63438 28358
rect 63238 28350 63250 28352
rect 62928 28320 63250 28350
rect 62928 28318 62940 28320
rect 62740 28312 62940 28318
rect 62520 28200 62590 28260
rect 62520 27940 62540 28200
rect 62580 27940 62590 28200
rect 63050 28310 63130 28320
rect 63238 28318 63250 28320
rect 63426 28318 63438 28352
rect 63470 28350 63480 28410
rect 63540 28350 63550 28410
rect 63470 28330 63550 28350
rect 63238 28312 63438 28318
rect 63050 28250 63060 28310
rect 63120 28250 63130 28310
rect 63050 28200 63130 28250
rect 63050 28140 63060 28200
rect 63120 28140 63130 28200
rect 62740 28130 62940 28136
rect 63050 28130 63130 28140
rect 63600 28260 63610 28500
rect 63650 28260 63670 28500
rect 63600 28180 63670 28260
rect 63238 28130 63438 28136
rect 62630 28100 62710 28120
rect 62630 28040 62640 28100
rect 62700 28086 62710 28100
rect 62740 28096 62752 28130
rect 62928 28100 63250 28130
rect 62928 28096 62940 28100
rect 62740 28090 62940 28096
rect 63238 28096 63250 28100
rect 63426 28096 63438 28130
rect 63238 28090 63438 28096
rect 63470 28100 63550 28120
rect 62702 28052 62710 28086
rect 62700 28040 62710 28052
rect 62630 28020 62710 28040
rect 62740 28042 62940 28048
rect 62740 28008 62752 28042
rect 62928 28040 62940 28042
rect 63238 28042 63438 28048
rect 63238 28040 63250 28042
rect 62928 28030 63250 28040
rect 62928 28010 63060 28030
rect 62928 28008 62940 28010
rect 62740 28002 62940 28008
rect 63050 27970 63060 28010
rect 63120 28010 63250 28030
rect 63120 27970 63130 28010
rect 63238 28008 63250 28010
rect 63426 28008 63438 28042
rect 63470 28040 63480 28100
rect 63540 28040 63550 28100
rect 63470 28020 63550 28040
rect 63238 28002 63438 28008
rect 63050 27960 63130 27970
rect 62520 27360 62590 27940
rect 63600 27940 63610 28180
rect 63650 27940 63670 28180
rect 63600 27530 63670 27940
rect 63660 27400 63670 27440
rect 63600 27360 63670 27390
rect 63700 27360 63730 29920
rect 64050 29590 64110 29600
rect 63850 29530 64050 29550
rect 67220 29590 67280 29600
rect 63850 29520 64110 29530
rect 64230 29530 64290 29540
rect 63760 29140 63820 29150
rect 63760 29070 63820 29080
rect 63790 27360 63820 29070
rect 63850 27360 63880 29520
rect 63970 29470 64230 29490
rect 63970 29460 64290 29470
rect 67040 29530 67100 29540
rect 67280 29530 67480 29550
rect 67220 29520 67480 29530
rect 67100 29470 67360 29490
rect 67040 29460 67360 29470
rect 63970 27360 64000 29460
rect 64090 27360 64120 29070
rect 64210 27360 64240 29070
rect 64330 27360 64360 29070
rect 64450 27360 64480 29070
rect 64570 27360 64600 29070
rect 66730 27360 66760 29070
rect 66850 27360 66880 29070
rect 66970 27360 67000 29070
rect 67090 27360 67120 29070
rect 67210 27360 67240 29070
rect 67330 27360 67360 29460
rect 67450 27360 67480 29520
rect 68580 29140 68660 29150
rect 67510 29080 67520 29140
rect 67580 29080 67590 29140
rect 67510 29070 67590 29080
rect 68580 29080 68590 29140
rect 68650 29080 68660 29140
rect 68580 29070 68660 29080
rect 67510 28960 67580 29070
rect 67510 28950 68660 28960
rect 67510 28890 67520 28950
rect 67580 28900 68660 28950
rect 67580 28890 67590 28900
rect 67510 28880 67590 28890
rect 67510 28500 67580 28880
rect 67510 28260 67530 28500
rect 67570 28260 67580 28500
rect 68590 28500 68660 28900
rect 68040 28480 68120 28490
rect 67730 28440 67930 28446
rect 68040 28440 68050 28480
rect 67620 28410 67700 28430
rect 67620 28350 67630 28410
rect 67690 28396 67700 28410
rect 67730 28406 67742 28440
rect 67918 28420 68050 28440
rect 68110 28440 68120 28480
rect 68228 28440 68428 28446
rect 68110 28420 68240 28440
rect 67918 28410 68240 28420
rect 67918 28406 67930 28410
rect 67730 28400 67930 28406
rect 68228 28406 68240 28410
rect 68416 28406 68428 28440
rect 68228 28400 68428 28406
rect 68460 28410 68540 28430
rect 67692 28362 67700 28396
rect 67690 28350 67700 28362
rect 67620 28330 67700 28350
rect 67730 28352 67930 28358
rect 67730 28318 67742 28352
rect 67918 28350 67930 28352
rect 68228 28352 68428 28358
rect 68228 28350 68240 28352
rect 67918 28320 68240 28350
rect 67918 28318 67930 28320
rect 67730 28312 67930 28318
rect 67510 28200 67580 28260
rect 67510 27940 67530 28200
rect 67570 27940 67580 28200
rect 68040 28310 68120 28320
rect 68228 28318 68240 28320
rect 68416 28318 68428 28352
rect 68460 28350 68470 28410
rect 68530 28350 68540 28410
rect 68460 28330 68540 28350
rect 68228 28312 68428 28318
rect 68040 28250 68050 28310
rect 68110 28250 68120 28310
rect 68040 28200 68120 28250
rect 68040 28140 68050 28200
rect 68110 28140 68120 28200
rect 67730 28130 67930 28136
rect 68040 28130 68120 28140
rect 68590 28260 68600 28500
rect 68640 28260 68660 28500
rect 68590 28180 68660 28260
rect 68228 28130 68428 28136
rect 67620 28100 67700 28120
rect 67620 28040 67630 28100
rect 67690 28086 67700 28100
rect 67730 28096 67742 28130
rect 67918 28100 68240 28130
rect 67918 28096 67930 28100
rect 67730 28090 67930 28096
rect 68228 28096 68240 28100
rect 68416 28096 68428 28130
rect 68228 28090 68428 28096
rect 68460 28100 68540 28120
rect 67692 28052 67700 28086
rect 67690 28040 67700 28052
rect 67620 28020 67700 28040
rect 67730 28042 67930 28048
rect 67730 28008 67742 28042
rect 67918 28040 67930 28042
rect 68228 28042 68428 28048
rect 68228 28040 68240 28042
rect 67918 28030 68240 28040
rect 67918 28010 68050 28030
rect 67918 28008 67930 28010
rect 67730 28002 67930 28008
rect 68040 27970 68050 28010
rect 68110 28010 68240 28030
rect 68110 27970 68120 28010
rect 68228 28008 68240 28010
rect 68416 28008 68428 28042
rect 68460 28040 68470 28100
rect 68530 28040 68540 28100
rect 68460 28020 68540 28040
rect 68228 28002 68428 28008
rect 68040 27960 68120 27970
rect 67510 27360 67580 27940
rect 68590 27940 68600 28180
rect 68640 27940 68660 28180
rect 68590 27530 68660 27940
rect 68650 27400 68660 27440
rect 68590 27360 68660 27390
rect 68690 27360 68720 29920
rect 69040 29590 69100 29600
rect 68840 29530 69040 29550
rect 72210 29590 72270 29600
rect 68840 29520 69100 29530
rect 69220 29530 69280 29540
rect 68750 29140 68810 29150
rect 68750 29070 68810 29080
rect 68780 27360 68810 29070
rect 68840 27360 68870 29520
rect 68960 29470 69220 29490
rect 72270 29530 72470 29550
rect 72210 29520 72470 29530
rect 68960 29460 69280 29470
rect 68960 27360 68990 29460
rect 69080 27360 69110 29070
rect 69200 27360 69230 29070
rect 69320 27360 69350 29070
rect 69440 27360 69470 29070
rect 69560 27360 69590 29070
rect 71720 27360 71750 29070
rect 71840 27360 71870 29070
rect 71960 27360 71990 29070
rect 72080 27360 72110 29070
rect 72200 27360 72230 29070
rect 72320 27360 72350 29070
rect 72440 27360 72470 29520
rect 73570 29140 73650 29150
rect 72500 29080 72510 29140
rect 72570 29080 72580 29140
rect 72500 29070 72580 29080
rect 73570 29080 73580 29140
rect 73640 29080 73650 29140
rect 73570 29070 73650 29080
rect 72500 28960 72570 29070
rect 72500 28950 73650 28960
rect 72500 28890 72510 28950
rect 72570 28900 73650 28950
rect 72570 28890 72580 28900
rect 72500 28880 72580 28890
rect 72500 28500 72570 28880
rect 72500 28260 72520 28500
rect 72560 28260 72570 28500
rect 73580 28500 73650 28900
rect 73030 28480 73110 28490
rect 72720 28440 72920 28446
rect 73030 28440 73040 28480
rect 72610 28410 72690 28430
rect 72610 28350 72620 28410
rect 72680 28396 72690 28410
rect 72720 28406 72732 28440
rect 72908 28420 73040 28440
rect 73100 28440 73110 28480
rect 73218 28440 73418 28446
rect 73100 28420 73230 28440
rect 72908 28410 73230 28420
rect 72908 28406 72920 28410
rect 72720 28400 72920 28406
rect 73218 28406 73230 28410
rect 73406 28406 73418 28440
rect 73218 28400 73418 28406
rect 73450 28410 73530 28430
rect 72682 28362 72690 28396
rect 72680 28350 72690 28362
rect 72610 28330 72690 28350
rect 72720 28352 72920 28358
rect 72720 28318 72732 28352
rect 72908 28350 72920 28352
rect 73218 28352 73418 28358
rect 73218 28350 73230 28352
rect 72908 28320 73230 28350
rect 72908 28318 72920 28320
rect 72720 28312 72920 28318
rect 72500 28200 72570 28260
rect 72500 27940 72520 28200
rect 72560 27940 72570 28200
rect 73030 28310 73110 28320
rect 73218 28318 73230 28320
rect 73406 28318 73418 28352
rect 73450 28350 73460 28410
rect 73520 28350 73530 28410
rect 73450 28330 73530 28350
rect 73218 28312 73418 28318
rect 73030 28250 73040 28310
rect 73100 28250 73110 28310
rect 73030 28200 73110 28250
rect 73030 28140 73040 28200
rect 73100 28140 73110 28200
rect 72720 28130 72920 28136
rect 73030 28130 73110 28140
rect 73580 28260 73590 28500
rect 73630 28260 73650 28500
rect 73580 28180 73650 28260
rect 73218 28130 73418 28136
rect 72610 28100 72690 28120
rect 72610 28040 72620 28100
rect 72680 28086 72690 28100
rect 72720 28096 72732 28130
rect 72908 28100 73230 28130
rect 72908 28096 72920 28100
rect 72720 28090 72920 28096
rect 73218 28096 73230 28100
rect 73406 28096 73418 28130
rect 73218 28090 73418 28096
rect 73450 28100 73530 28120
rect 72682 28052 72690 28086
rect 72680 28040 72690 28052
rect 72610 28020 72690 28040
rect 72720 28042 72920 28048
rect 72720 28008 72732 28042
rect 72908 28040 72920 28042
rect 73218 28042 73418 28048
rect 73218 28040 73230 28042
rect 72908 28030 73230 28040
rect 72908 28010 73040 28030
rect 72908 28008 72920 28010
rect 72720 28002 72920 28008
rect 73030 27970 73040 28010
rect 73100 28010 73230 28030
rect 73100 27970 73110 28010
rect 73218 28008 73230 28010
rect 73406 28008 73418 28042
rect 73450 28040 73460 28100
rect 73520 28040 73530 28100
rect 73450 28020 73530 28040
rect 73218 28002 73418 28008
rect 73030 27960 73110 27970
rect 72500 27360 72570 27940
rect 73580 27940 73590 28180
rect 73630 27940 73650 28180
rect 73580 27530 73650 27940
rect 73640 27400 73650 27440
rect 73580 27360 73650 27390
rect 73680 27360 73710 29920
rect 74030 29590 74090 29600
rect 73830 29530 74030 29550
rect 73830 29520 74090 29530
rect 77200 29590 77260 29600
rect 77260 29530 77460 29550
rect 77200 29520 77460 29530
rect 73740 29140 73800 29150
rect 73740 29070 73800 29080
rect 73770 27360 73800 29070
rect 73830 27360 73860 29520
rect 73950 27360 73980 29070
rect 74070 27360 74100 29070
rect 74190 27360 74220 29070
rect 74310 27360 74340 29070
rect 74430 27360 74460 29070
rect 74550 27360 74580 29070
rect 76710 27360 76740 29070
rect 76830 27360 76860 29070
rect 76950 27360 76980 29070
rect 77070 27360 77100 29070
rect 77190 27360 77220 29070
rect 77310 27360 77340 29070
rect 77430 27360 77460 29520
rect 78560 29140 78640 29150
rect 77490 29080 77500 29140
rect 77560 29080 77570 29140
rect 77490 29070 77570 29080
rect 78560 29080 78570 29140
rect 78630 29080 78640 29140
rect 78560 29070 78640 29080
rect 77490 28960 77560 29070
rect 77490 28950 78640 28960
rect 77490 28890 77500 28950
rect 77560 28900 78640 28950
rect 77560 28890 77570 28900
rect 77490 28880 77570 28890
rect 77490 28500 77560 28880
rect 77490 28260 77510 28500
rect 77550 28260 77560 28500
rect 78570 28500 78640 28900
rect 78020 28480 78100 28490
rect 77710 28440 77910 28446
rect 78020 28440 78030 28480
rect 77600 28410 77680 28430
rect 77600 28350 77610 28410
rect 77670 28396 77680 28410
rect 77710 28406 77722 28440
rect 77898 28420 78030 28440
rect 78090 28440 78100 28480
rect 78208 28440 78408 28446
rect 78090 28420 78220 28440
rect 77898 28410 78220 28420
rect 77898 28406 77910 28410
rect 77710 28400 77910 28406
rect 78208 28406 78220 28410
rect 78396 28406 78408 28440
rect 78208 28400 78408 28406
rect 78440 28410 78520 28430
rect 77672 28362 77680 28396
rect 77670 28350 77680 28362
rect 77600 28330 77680 28350
rect 77710 28352 77910 28358
rect 77710 28318 77722 28352
rect 77898 28350 77910 28352
rect 78208 28352 78408 28358
rect 78208 28350 78220 28352
rect 77898 28320 78220 28350
rect 77898 28318 77910 28320
rect 77710 28312 77910 28318
rect 77490 28200 77560 28260
rect 77490 27940 77510 28200
rect 77550 27940 77560 28200
rect 78020 28310 78100 28320
rect 78208 28318 78220 28320
rect 78396 28318 78408 28352
rect 78440 28350 78450 28410
rect 78510 28350 78520 28410
rect 78440 28330 78520 28350
rect 78208 28312 78408 28318
rect 78020 28250 78030 28310
rect 78090 28250 78100 28310
rect 78020 28200 78100 28250
rect 78020 28140 78030 28200
rect 78090 28140 78100 28200
rect 77710 28130 77910 28136
rect 78020 28130 78100 28140
rect 78570 28260 78580 28500
rect 78620 28260 78640 28500
rect 78570 28180 78640 28260
rect 78208 28130 78408 28136
rect 77600 28100 77680 28120
rect 77600 28040 77610 28100
rect 77670 28086 77680 28100
rect 77710 28096 77722 28130
rect 77898 28100 78220 28130
rect 77898 28096 77910 28100
rect 77710 28090 77910 28096
rect 78208 28096 78220 28100
rect 78396 28096 78408 28130
rect 78208 28090 78408 28096
rect 78440 28100 78520 28120
rect 77672 28052 77680 28086
rect 77670 28040 77680 28052
rect 77600 28020 77680 28040
rect 77710 28042 77910 28048
rect 77710 28008 77722 28042
rect 77898 28040 77910 28042
rect 78208 28042 78408 28048
rect 78208 28040 78220 28042
rect 77898 28030 78220 28040
rect 77898 28010 78030 28030
rect 77898 28008 77910 28010
rect 77710 28002 77910 28008
rect 78020 27970 78030 28010
rect 78090 28010 78220 28030
rect 78090 27970 78100 28010
rect 78208 28008 78220 28010
rect 78396 28008 78408 28042
rect 78440 28040 78450 28100
rect 78510 28040 78520 28100
rect 78440 28020 78520 28040
rect 78208 28002 78408 28008
rect 78020 27960 78100 27970
rect 77490 27360 77560 27940
rect 78570 27940 78580 28180
rect 78620 27940 78640 28180
rect 78570 27530 78640 27940
rect 78630 27400 78640 27440
rect 78570 27360 78640 27390
rect 78670 27360 78700 29920
rect 79020 29590 79080 29600
rect 78820 29530 79020 29550
rect 78820 29520 79080 29530
rect 78730 29140 78790 29150
rect 78730 29070 78790 29080
rect 78760 27360 78790 29070
rect 78820 27360 78850 29520
rect 82210 29080 82220 29140
rect 82280 29080 82290 29140
rect 82210 29070 82290 29080
rect 78940 27360 78970 29070
rect 79060 27360 79090 29070
rect 79180 27360 79210 29070
rect 79300 27360 79330 29070
rect 79420 27360 79450 29070
rect 79540 27360 79570 29070
rect -940 25690 -930 25710
rect -2860 -1710 -2830 23940
rect -2740 -1710 -2710 23940
rect -2620 -1710 -2590 23940
rect -2500 -1710 -2470 23940
rect -2380 -1710 -2350 23940
rect -2260 -1710 -2230 23940
rect -2140 -1710 -2110 23940
rect -2080 23830 -2010 23940
rect -1010 23930 -930 23940
rect -1010 23870 -1000 23930
rect -940 23870 -930 23930
rect -1010 23860 -930 23870
rect -2080 23820 -930 23830
rect -2080 23760 -2070 23820
rect -2010 23770 -930 23820
rect -2010 23760 -2000 23770
rect -2080 23750 -2000 23760
rect -2080 23370 -2010 23750
rect -2080 23130 -2060 23370
rect -2020 23130 -2010 23370
rect -1000 23370 -930 23770
rect -1550 23350 -1470 23360
rect -1860 23310 -1660 23316
rect -1550 23310 -1540 23350
rect -1970 23280 -1890 23300
rect -1970 23220 -1960 23280
rect -1900 23266 -1890 23280
rect -1860 23276 -1848 23310
rect -1672 23290 -1540 23310
rect -1480 23310 -1470 23350
rect -1362 23310 -1162 23316
rect -1480 23290 -1350 23310
rect -1672 23280 -1350 23290
rect -1672 23276 -1660 23280
rect -1860 23270 -1660 23276
rect -1362 23276 -1350 23280
rect -1174 23276 -1162 23310
rect -1362 23270 -1162 23276
rect -1130 23280 -1050 23300
rect -1898 23232 -1890 23266
rect -1900 23220 -1890 23232
rect -1970 23200 -1890 23220
rect -1860 23222 -1660 23228
rect -1860 23188 -1848 23222
rect -1672 23220 -1660 23222
rect -1362 23222 -1162 23228
rect -1362 23220 -1350 23222
rect -1672 23190 -1350 23220
rect -1672 23188 -1660 23190
rect -1860 23182 -1660 23188
rect -2080 23070 -2010 23130
rect -2080 22810 -2060 23070
rect -2020 22810 -2010 23070
rect -1550 23180 -1470 23190
rect -1362 23188 -1350 23190
rect -1174 23188 -1162 23222
rect -1130 23220 -1120 23280
rect -1060 23220 -1050 23280
rect -1130 23200 -1050 23220
rect -1362 23182 -1162 23188
rect -1550 23120 -1540 23180
rect -1480 23120 -1470 23180
rect -1550 23070 -1470 23120
rect -1550 23010 -1540 23070
rect -1480 23010 -1470 23070
rect -1860 23000 -1660 23006
rect -1550 23000 -1470 23010
rect -1000 23130 -990 23370
rect -950 23130 -930 23370
rect -1000 23050 -930 23130
rect -1362 23000 -1162 23006
rect -1970 22970 -1890 22990
rect -1970 22910 -1960 22970
rect -1900 22956 -1890 22970
rect -1860 22966 -1848 23000
rect -1672 22970 -1350 23000
rect -1672 22966 -1660 22970
rect -1860 22960 -1660 22966
rect -1362 22966 -1350 22970
rect -1174 22966 -1162 23000
rect -1362 22960 -1162 22966
rect -1130 22970 -1050 22990
rect -1898 22922 -1890 22956
rect -1900 22910 -1890 22922
rect -1970 22890 -1890 22910
rect -1860 22912 -1660 22918
rect -1860 22878 -1848 22912
rect -1672 22910 -1660 22912
rect -1362 22912 -1162 22918
rect -1362 22910 -1350 22912
rect -1672 22900 -1350 22910
rect -1672 22880 -1540 22900
rect -1672 22878 -1660 22880
rect -1860 22872 -1660 22878
rect -1550 22840 -1540 22880
rect -1480 22880 -1350 22900
rect -1480 22840 -1470 22880
rect -1362 22878 -1350 22880
rect -1174 22878 -1162 22912
rect -1130 22910 -1120 22970
rect -1060 22910 -1050 22970
rect -1130 22890 -1050 22910
rect -1362 22872 -1162 22878
rect -1550 22830 -1470 22840
rect -2080 22120 -2010 22810
rect -1000 22810 -990 23050
rect -950 22810 -930 23050
rect -1000 22400 -930 22810
rect -1020 22360 -930 22370
rect -1020 22300 -1010 22360
rect -940 22300 -930 22360
rect -1020 22290 -930 22300
rect -1000 22230 -930 22290
rect -1010 22220 -930 22230
rect -1010 22160 -1000 22220
rect -940 22160 -930 22220
rect -1010 22150 -930 22160
rect -2080 22110 -930 22120
rect -2080 22050 -2070 22110
rect -2010 22060 -930 22110
rect -2010 22050 -2000 22060
rect -2080 22040 -2000 22050
rect -2080 21660 -2010 22040
rect -2080 21420 -2060 21660
rect -2020 21420 -2010 21660
rect -1000 21660 -930 22060
rect -1550 21640 -1470 21650
rect -1860 21600 -1660 21606
rect -1550 21600 -1540 21640
rect -1970 21570 -1890 21590
rect -1970 21510 -1960 21570
rect -1900 21556 -1890 21570
rect -1860 21566 -1848 21600
rect -1672 21580 -1540 21600
rect -1480 21600 -1470 21640
rect -1362 21600 -1162 21606
rect -1480 21580 -1350 21600
rect -1672 21570 -1350 21580
rect -1672 21566 -1660 21570
rect -1860 21560 -1660 21566
rect -1362 21566 -1350 21570
rect -1174 21566 -1162 21600
rect -1362 21560 -1162 21566
rect -1130 21570 -1050 21590
rect -1898 21522 -1890 21556
rect -1900 21510 -1890 21522
rect -1970 21490 -1890 21510
rect -1860 21512 -1660 21518
rect -1860 21478 -1848 21512
rect -1672 21510 -1660 21512
rect -1362 21512 -1162 21518
rect -1362 21510 -1350 21512
rect -1672 21480 -1350 21510
rect -1672 21478 -1660 21480
rect -1860 21472 -1660 21478
rect -2080 21360 -2010 21420
rect -2080 21100 -2060 21360
rect -2020 21100 -2010 21360
rect -1550 21470 -1470 21480
rect -1362 21478 -1350 21480
rect -1174 21478 -1162 21512
rect -1130 21510 -1120 21570
rect -1060 21510 -1050 21570
rect -1130 21490 -1050 21510
rect -1362 21472 -1162 21478
rect -1550 21410 -1540 21470
rect -1480 21410 -1470 21470
rect -1550 21360 -1470 21410
rect -1550 21300 -1540 21360
rect -1480 21300 -1470 21360
rect -1860 21290 -1660 21296
rect -1550 21290 -1470 21300
rect -1000 21420 -990 21660
rect -950 21420 -930 21660
rect -1000 21340 -930 21420
rect -1362 21290 -1162 21296
rect -1970 21260 -1890 21280
rect -1970 21200 -1960 21260
rect -1900 21246 -1890 21260
rect -1860 21256 -1848 21290
rect -1672 21260 -1350 21290
rect -1672 21256 -1660 21260
rect -1860 21250 -1660 21256
rect -1362 21256 -1350 21260
rect -1174 21256 -1162 21290
rect -1362 21250 -1162 21256
rect -1130 21260 -1050 21280
rect -1898 21212 -1890 21246
rect -1900 21200 -1890 21212
rect -1970 21180 -1890 21200
rect -1860 21202 -1660 21208
rect -1860 21168 -1848 21202
rect -1672 21200 -1660 21202
rect -1362 21202 -1162 21208
rect -1362 21200 -1350 21202
rect -1672 21190 -1350 21200
rect -1672 21170 -1540 21190
rect -1672 21168 -1660 21170
rect -1860 21162 -1660 21168
rect -1550 21130 -1540 21170
rect -1480 21170 -1350 21190
rect -1480 21130 -1470 21170
rect -1362 21168 -1350 21170
rect -1174 21168 -1162 21202
rect -1130 21200 -1120 21260
rect -1060 21200 -1050 21260
rect -1130 21180 -1050 21200
rect -1362 21162 -1162 21168
rect -1550 21120 -1470 21130
rect -2080 20410 -2010 21100
rect -1000 21100 -990 21340
rect -950 21100 -930 21340
rect -1000 20690 -930 21100
rect -1020 20650 -930 20660
rect -1020 20590 -1010 20650
rect -940 20590 -930 20650
rect -1020 20580 -930 20590
rect -1000 20520 -930 20580
rect -1010 20510 -930 20520
rect -1010 20450 -1000 20510
rect -940 20450 -930 20510
rect -1010 20440 -930 20450
rect -2080 20400 -930 20410
rect -2080 20340 -2070 20400
rect -2010 20350 -930 20400
rect -2010 20340 -2000 20350
rect -2080 20330 -2000 20340
rect -2080 19950 -2010 20330
rect -2080 19710 -2060 19950
rect -2020 19710 -2010 19950
rect -1000 19950 -930 20350
rect -1550 19930 -1470 19940
rect -1860 19890 -1660 19896
rect -1550 19890 -1540 19930
rect -1970 19860 -1890 19880
rect -1970 19800 -1960 19860
rect -1900 19846 -1890 19860
rect -1860 19856 -1848 19890
rect -1672 19870 -1540 19890
rect -1480 19890 -1470 19930
rect -1362 19890 -1162 19896
rect -1480 19870 -1350 19890
rect -1672 19860 -1350 19870
rect -1672 19856 -1660 19860
rect -1860 19850 -1660 19856
rect -1362 19856 -1350 19860
rect -1174 19856 -1162 19890
rect -1362 19850 -1162 19856
rect -1130 19860 -1050 19880
rect -1898 19812 -1890 19846
rect -1900 19800 -1890 19812
rect -1970 19780 -1890 19800
rect -1860 19802 -1660 19808
rect -1860 19768 -1848 19802
rect -1672 19800 -1660 19802
rect -1362 19802 -1162 19808
rect -1362 19800 -1350 19802
rect -1672 19770 -1350 19800
rect -1672 19768 -1660 19770
rect -1860 19762 -1660 19768
rect -2080 19650 -2010 19710
rect -2080 19390 -2060 19650
rect -2020 19390 -2010 19650
rect -1550 19760 -1470 19770
rect -1362 19768 -1350 19770
rect -1174 19768 -1162 19802
rect -1130 19800 -1120 19860
rect -1060 19800 -1050 19860
rect -1130 19780 -1050 19800
rect -1362 19762 -1162 19768
rect -1550 19700 -1540 19760
rect -1480 19700 -1470 19760
rect -1550 19650 -1470 19700
rect -1550 19590 -1540 19650
rect -1480 19590 -1470 19650
rect -1860 19580 -1660 19586
rect -1550 19580 -1470 19590
rect -1000 19710 -990 19950
rect -950 19710 -930 19950
rect -1000 19630 -930 19710
rect -1362 19580 -1162 19586
rect -1970 19550 -1890 19570
rect -1970 19490 -1960 19550
rect -1900 19536 -1890 19550
rect -1860 19546 -1848 19580
rect -1672 19550 -1350 19580
rect -1672 19546 -1660 19550
rect -1860 19540 -1660 19546
rect -1362 19546 -1350 19550
rect -1174 19546 -1162 19580
rect -1362 19540 -1162 19546
rect -1130 19550 -1050 19570
rect -1898 19502 -1890 19536
rect -1900 19490 -1890 19502
rect -1970 19470 -1890 19490
rect -1860 19492 -1660 19498
rect -1860 19458 -1848 19492
rect -1672 19490 -1660 19492
rect -1362 19492 -1162 19498
rect -1362 19490 -1350 19492
rect -1672 19480 -1350 19490
rect -1672 19460 -1540 19480
rect -1672 19458 -1660 19460
rect -1860 19452 -1660 19458
rect -1550 19420 -1540 19460
rect -1480 19460 -1350 19480
rect -1480 19420 -1470 19460
rect -1362 19458 -1350 19460
rect -1174 19458 -1162 19492
rect -1130 19490 -1120 19550
rect -1060 19490 -1050 19550
rect -1130 19470 -1050 19490
rect -1362 19452 -1162 19458
rect -1550 19410 -1470 19420
rect -2080 18700 -2010 19390
rect -1000 19390 -990 19630
rect -950 19390 -930 19630
rect -1000 18980 -930 19390
rect -1020 18940 -930 18950
rect -1020 18880 -1010 18940
rect -940 18880 -930 18940
rect -1020 18870 -930 18880
rect -1000 18810 -930 18870
rect -1010 18800 -930 18810
rect -1010 18740 -1000 18800
rect -940 18740 -930 18800
rect -1010 18730 -930 18740
rect -2080 18690 -930 18700
rect -2080 18630 -2070 18690
rect -2010 18640 -930 18690
rect -2010 18630 -2000 18640
rect -2080 18620 -2000 18630
rect -2080 18240 -2010 18620
rect -2080 18000 -2060 18240
rect -2020 18000 -2010 18240
rect -1000 18240 -930 18640
rect -1550 18220 -1470 18230
rect -1860 18180 -1660 18186
rect -1550 18180 -1540 18220
rect -1970 18150 -1890 18170
rect -1970 18090 -1960 18150
rect -1900 18136 -1890 18150
rect -1860 18146 -1848 18180
rect -1672 18160 -1540 18180
rect -1480 18180 -1470 18220
rect -1362 18180 -1162 18186
rect -1480 18160 -1350 18180
rect -1672 18150 -1350 18160
rect -1672 18146 -1660 18150
rect -1860 18140 -1660 18146
rect -1362 18146 -1350 18150
rect -1174 18146 -1162 18180
rect -1362 18140 -1162 18146
rect -1130 18150 -1050 18170
rect -1898 18102 -1890 18136
rect -1900 18090 -1890 18102
rect -1970 18070 -1890 18090
rect -1860 18092 -1660 18098
rect -1860 18058 -1848 18092
rect -1672 18090 -1660 18092
rect -1362 18092 -1162 18098
rect -1362 18090 -1350 18092
rect -1672 18060 -1350 18090
rect -1672 18058 -1660 18060
rect -1860 18052 -1660 18058
rect -2080 17940 -2010 18000
rect -2080 17680 -2060 17940
rect -2020 17680 -2010 17940
rect -1550 18050 -1470 18060
rect -1362 18058 -1350 18060
rect -1174 18058 -1162 18092
rect -1130 18090 -1120 18150
rect -1060 18090 -1050 18150
rect -1130 18070 -1050 18090
rect -1362 18052 -1162 18058
rect -1550 17990 -1540 18050
rect -1480 17990 -1470 18050
rect -1550 17940 -1470 17990
rect -1550 17880 -1540 17940
rect -1480 17880 -1470 17940
rect -1860 17870 -1660 17876
rect -1550 17870 -1470 17880
rect -1000 18000 -990 18240
rect -950 18000 -930 18240
rect -1000 17920 -930 18000
rect -1362 17870 -1162 17876
rect -1970 17840 -1890 17860
rect -1970 17780 -1960 17840
rect -1900 17826 -1890 17840
rect -1860 17836 -1848 17870
rect -1672 17840 -1350 17870
rect -1672 17836 -1660 17840
rect -1860 17830 -1660 17836
rect -1362 17836 -1350 17840
rect -1174 17836 -1162 17870
rect -1362 17830 -1162 17836
rect -1130 17840 -1050 17860
rect -1898 17792 -1890 17826
rect -1900 17780 -1890 17792
rect -1970 17760 -1890 17780
rect -1860 17782 -1660 17788
rect -1860 17748 -1848 17782
rect -1672 17780 -1660 17782
rect -1362 17782 -1162 17788
rect -1362 17780 -1350 17782
rect -1672 17770 -1350 17780
rect -1672 17750 -1540 17770
rect -1672 17748 -1660 17750
rect -1860 17742 -1660 17748
rect -1550 17710 -1540 17750
rect -1480 17750 -1350 17770
rect -1480 17710 -1470 17750
rect -1362 17748 -1350 17750
rect -1174 17748 -1162 17782
rect -1130 17780 -1120 17840
rect -1060 17780 -1050 17840
rect -1130 17760 -1050 17780
rect -1362 17742 -1162 17748
rect -1550 17700 -1470 17710
rect -2080 16990 -2010 17680
rect -1000 17680 -990 17920
rect -950 17680 -930 17920
rect -1000 17270 -930 17680
rect -1020 17230 -930 17240
rect -1020 17170 -1010 17230
rect -940 17170 -930 17230
rect -1020 17160 -930 17170
rect -1000 17100 -930 17160
rect -1010 17090 -930 17100
rect -1010 17030 -1000 17090
rect -940 17030 -930 17090
rect -1010 17020 -930 17030
rect -2080 16980 -930 16990
rect -2080 16920 -2070 16980
rect -2010 16930 -930 16980
rect -2010 16920 -2000 16930
rect -2080 16910 -2000 16920
rect -2080 16530 -2010 16910
rect -2080 16290 -2060 16530
rect -2020 16290 -2010 16530
rect -1000 16530 -930 16930
rect -1550 16510 -1470 16520
rect -1860 16470 -1660 16476
rect -1550 16470 -1540 16510
rect -1970 16440 -1890 16460
rect -1970 16380 -1960 16440
rect -1900 16426 -1890 16440
rect -1860 16436 -1848 16470
rect -1672 16450 -1540 16470
rect -1480 16470 -1470 16510
rect -1362 16470 -1162 16476
rect -1480 16450 -1350 16470
rect -1672 16440 -1350 16450
rect -1672 16436 -1660 16440
rect -1860 16430 -1660 16436
rect -1362 16436 -1350 16440
rect -1174 16436 -1162 16470
rect -1362 16430 -1162 16436
rect -1130 16440 -1050 16460
rect -1898 16392 -1890 16426
rect -1900 16380 -1890 16392
rect -1970 16360 -1890 16380
rect -1860 16382 -1660 16388
rect -1860 16348 -1848 16382
rect -1672 16380 -1660 16382
rect -1362 16382 -1162 16388
rect -1362 16380 -1350 16382
rect -1672 16350 -1350 16380
rect -1672 16348 -1660 16350
rect -1860 16342 -1660 16348
rect -2080 16230 -2010 16290
rect -2080 15970 -2060 16230
rect -2020 15970 -2010 16230
rect -1550 16340 -1470 16350
rect -1362 16348 -1350 16350
rect -1174 16348 -1162 16382
rect -1130 16380 -1120 16440
rect -1060 16380 -1050 16440
rect -1130 16360 -1050 16380
rect -1362 16342 -1162 16348
rect -1550 16280 -1540 16340
rect -1480 16280 -1470 16340
rect -1550 16230 -1470 16280
rect -1550 16170 -1540 16230
rect -1480 16170 -1470 16230
rect -1860 16160 -1660 16166
rect -1550 16160 -1470 16170
rect -1000 16290 -990 16530
rect -950 16290 -930 16530
rect -1000 16210 -930 16290
rect -1362 16160 -1162 16166
rect -1970 16130 -1890 16150
rect -1970 16070 -1960 16130
rect -1900 16116 -1890 16130
rect -1860 16126 -1848 16160
rect -1672 16130 -1350 16160
rect -1672 16126 -1660 16130
rect -1860 16120 -1660 16126
rect -1362 16126 -1350 16130
rect -1174 16126 -1162 16160
rect -1362 16120 -1162 16126
rect -1130 16130 -1050 16150
rect -1898 16082 -1890 16116
rect -1900 16070 -1890 16082
rect -1970 16050 -1890 16070
rect -1860 16072 -1660 16078
rect -1860 16038 -1848 16072
rect -1672 16070 -1660 16072
rect -1362 16072 -1162 16078
rect -1362 16070 -1350 16072
rect -1672 16060 -1350 16070
rect -1672 16040 -1540 16060
rect -1672 16038 -1660 16040
rect -1860 16032 -1660 16038
rect -1550 16000 -1540 16040
rect -1480 16040 -1350 16060
rect -1480 16000 -1470 16040
rect -1362 16038 -1350 16040
rect -1174 16038 -1162 16072
rect -1130 16070 -1120 16130
rect -1060 16070 -1050 16130
rect -1130 16050 -1050 16070
rect -1362 16032 -1162 16038
rect -1550 15990 -1470 16000
rect -2080 15280 -2010 15970
rect -1000 15970 -990 16210
rect -950 15970 -930 16210
rect -1000 15560 -930 15970
rect -1020 15520 -930 15530
rect -1020 15460 -1010 15520
rect -940 15460 -930 15520
rect -1020 15450 -930 15460
rect -1000 15390 -930 15450
rect -1010 15380 -930 15390
rect -1010 15320 -1000 15380
rect -940 15320 -930 15380
rect -1010 15310 -930 15320
rect -2080 15270 -930 15280
rect -2080 15210 -2070 15270
rect -2010 15220 -930 15270
rect -2010 15210 -2000 15220
rect -2080 15200 -2000 15210
rect -2080 14820 -2010 15200
rect -2080 14580 -2060 14820
rect -2020 14580 -2010 14820
rect -1000 14820 -930 15220
rect -1550 14800 -1470 14810
rect -1860 14760 -1660 14766
rect -1550 14760 -1540 14800
rect -1970 14730 -1890 14750
rect -1970 14670 -1960 14730
rect -1900 14716 -1890 14730
rect -1860 14726 -1848 14760
rect -1672 14740 -1540 14760
rect -1480 14760 -1470 14800
rect -1362 14760 -1162 14766
rect -1480 14740 -1350 14760
rect -1672 14730 -1350 14740
rect -1672 14726 -1660 14730
rect -1860 14720 -1660 14726
rect -1362 14726 -1350 14730
rect -1174 14726 -1162 14760
rect -1362 14720 -1162 14726
rect -1130 14730 -1050 14750
rect -1898 14682 -1890 14716
rect -1900 14670 -1890 14682
rect -1970 14650 -1890 14670
rect -1860 14672 -1660 14678
rect -1860 14638 -1848 14672
rect -1672 14670 -1660 14672
rect -1362 14672 -1162 14678
rect -1362 14670 -1350 14672
rect -1672 14640 -1350 14670
rect -1672 14638 -1660 14640
rect -1860 14632 -1660 14638
rect -2080 14520 -2010 14580
rect -2080 14260 -2060 14520
rect -2020 14260 -2010 14520
rect -1550 14630 -1470 14640
rect -1362 14638 -1350 14640
rect -1174 14638 -1162 14672
rect -1130 14670 -1120 14730
rect -1060 14670 -1050 14730
rect -1130 14650 -1050 14670
rect -1362 14632 -1162 14638
rect -1550 14570 -1540 14630
rect -1480 14570 -1470 14630
rect -1550 14520 -1470 14570
rect -1550 14460 -1540 14520
rect -1480 14460 -1470 14520
rect -1860 14450 -1660 14456
rect -1550 14450 -1470 14460
rect -1000 14580 -990 14820
rect -950 14580 -930 14820
rect -1000 14500 -930 14580
rect -1362 14450 -1162 14456
rect -1970 14420 -1890 14440
rect -1970 14360 -1960 14420
rect -1900 14406 -1890 14420
rect -1860 14416 -1848 14450
rect -1672 14420 -1350 14450
rect -1672 14416 -1660 14420
rect -1860 14410 -1660 14416
rect -1362 14416 -1350 14420
rect -1174 14416 -1162 14450
rect -1362 14410 -1162 14416
rect -1130 14420 -1050 14440
rect -1898 14372 -1890 14406
rect -1900 14360 -1890 14372
rect -1970 14340 -1890 14360
rect -1860 14362 -1660 14368
rect -1860 14328 -1848 14362
rect -1672 14360 -1660 14362
rect -1362 14362 -1162 14368
rect -1362 14360 -1350 14362
rect -1672 14350 -1350 14360
rect -1672 14330 -1540 14350
rect -1672 14328 -1660 14330
rect -1860 14322 -1660 14328
rect -1550 14290 -1540 14330
rect -1480 14330 -1350 14350
rect -1480 14290 -1470 14330
rect -1362 14328 -1350 14330
rect -1174 14328 -1162 14362
rect -1130 14360 -1120 14420
rect -1060 14360 -1050 14420
rect -1130 14340 -1050 14360
rect -1362 14322 -1162 14328
rect -1550 14280 -1470 14290
rect -2080 13570 -2010 14260
rect -1000 14260 -990 14500
rect -950 14260 -930 14500
rect -1000 13850 -930 14260
rect -1020 13810 -930 13820
rect -1020 13750 -1010 13810
rect -940 13750 -930 13810
rect -1020 13740 -930 13750
rect -1000 13680 -930 13740
rect -1010 13670 -930 13680
rect -1010 13610 -1000 13670
rect -940 13610 -930 13670
rect -1010 13600 -930 13610
rect -2080 13560 -930 13570
rect -2080 13500 -2070 13560
rect -2010 13510 -930 13560
rect -2010 13500 -2000 13510
rect -2080 13490 -2000 13500
rect -2080 13110 -2010 13490
rect -2080 12870 -2060 13110
rect -2020 12870 -2010 13110
rect -1000 13110 -930 13510
rect -1550 13090 -1470 13100
rect -1860 13050 -1660 13056
rect -1550 13050 -1540 13090
rect -1970 13020 -1890 13040
rect -1970 12960 -1960 13020
rect -1900 13006 -1890 13020
rect -1860 13016 -1848 13050
rect -1672 13030 -1540 13050
rect -1480 13050 -1470 13090
rect -1362 13050 -1162 13056
rect -1480 13030 -1350 13050
rect -1672 13020 -1350 13030
rect -1672 13016 -1660 13020
rect -1860 13010 -1660 13016
rect -1362 13016 -1350 13020
rect -1174 13016 -1162 13050
rect -1362 13010 -1162 13016
rect -1130 13020 -1050 13040
rect -1898 12972 -1890 13006
rect -1900 12960 -1890 12972
rect -1970 12940 -1890 12960
rect -1860 12962 -1660 12968
rect -1860 12928 -1848 12962
rect -1672 12960 -1660 12962
rect -1362 12962 -1162 12968
rect -1362 12960 -1350 12962
rect -1672 12930 -1350 12960
rect -1672 12928 -1660 12930
rect -1860 12922 -1660 12928
rect -2080 12810 -2010 12870
rect -2080 12550 -2060 12810
rect -2020 12550 -2010 12810
rect -1550 12920 -1470 12930
rect -1362 12928 -1350 12930
rect -1174 12928 -1162 12962
rect -1130 12960 -1120 13020
rect -1060 12960 -1050 13020
rect -1130 12940 -1050 12960
rect -1362 12922 -1162 12928
rect -1550 12860 -1540 12920
rect -1480 12860 -1470 12920
rect -1550 12810 -1470 12860
rect -1550 12750 -1540 12810
rect -1480 12750 -1470 12810
rect -1860 12740 -1660 12746
rect -1550 12740 -1470 12750
rect -1000 12870 -990 13110
rect -950 12870 -930 13110
rect -1000 12790 -930 12870
rect -1362 12740 -1162 12746
rect -1970 12710 -1890 12730
rect -1970 12650 -1960 12710
rect -1900 12696 -1890 12710
rect -1860 12706 -1848 12740
rect -1672 12710 -1350 12740
rect -1672 12706 -1660 12710
rect -1860 12700 -1660 12706
rect -1362 12706 -1350 12710
rect -1174 12706 -1162 12740
rect -1362 12700 -1162 12706
rect -1130 12710 -1050 12730
rect -1898 12662 -1890 12696
rect -1900 12650 -1890 12662
rect -1970 12630 -1890 12650
rect -1860 12652 -1660 12658
rect -1860 12618 -1848 12652
rect -1672 12650 -1660 12652
rect -1362 12652 -1162 12658
rect -1362 12650 -1350 12652
rect -1672 12640 -1350 12650
rect -1672 12620 -1540 12640
rect -1672 12618 -1660 12620
rect -1860 12612 -1660 12618
rect -1550 12580 -1540 12620
rect -1480 12620 -1350 12640
rect -1480 12580 -1470 12620
rect -1362 12618 -1350 12620
rect -1174 12618 -1162 12652
rect -1130 12650 -1120 12710
rect -1060 12650 -1050 12710
rect -1130 12630 -1050 12650
rect -1362 12612 -1162 12618
rect -1550 12570 -1470 12580
rect -2080 11860 -2010 12550
rect -1000 12550 -990 12790
rect -950 12550 -930 12790
rect -1000 12140 -930 12550
rect -1020 12100 -930 12110
rect -1020 12040 -1010 12100
rect -940 12040 -930 12100
rect -1020 12030 -930 12040
rect -1000 11970 -930 12030
rect -1010 11960 -930 11970
rect -1010 11900 -1000 11960
rect -940 11900 -930 11960
rect -1010 11890 -930 11900
rect -2080 11850 -930 11860
rect -2080 11790 -2070 11850
rect -2010 11800 -930 11850
rect -2010 11790 -2000 11800
rect -2080 11780 -2000 11790
rect -2080 11400 -2010 11780
rect -2080 11160 -2060 11400
rect -2020 11160 -2010 11400
rect -1000 11400 -930 11800
rect -1550 11380 -1470 11390
rect -1860 11340 -1660 11346
rect -1550 11340 -1540 11380
rect -1970 11310 -1890 11330
rect -1970 11250 -1960 11310
rect -1900 11296 -1890 11310
rect -1860 11306 -1848 11340
rect -1672 11320 -1540 11340
rect -1480 11340 -1470 11380
rect -1362 11340 -1162 11346
rect -1480 11320 -1350 11340
rect -1672 11310 -1350 11320
rect -1672 11306 -1660 11310
rect -1860 11300 -1660 11306
rect -1362 11306 -1350 11310
rect -1174 11306 -1162 11340
rect -1362 11300 -1162 11306
rect -1130 11310 -1050 11330
rect -1898 11262 -1890 11296
rect -1900 11250 -1890 11262
rect -1970 11230 -1890 11250
rect -1860 11252 -1660 11258
rect -1860 11218 -1848 11252
rect -1672 11250 -1660 11252
rect -1362 11252 -1162 11258
rect -1362 11250 -1350 11252
rect -1672 11220 -1350 11250
rect -1672 11218 -1660 11220
rect -1860 11212 -1660 11218
rect -2080 11100 -2010 11160
rect -2080 10840 -2060 11100
rect -2020 10840 -2010 11100
rect -1550 11210 -1470 11220
rect -1362 11218 -1350 11220
rect -1174 11218 -1162 11252
rect -1130 11250 -1120 11310
rect -1060 11250 -1050 11310
rect -1130 11230 -1050 11250
rect -1362 11212 -1162 11218
rect -1550 11150 -1540 11210
rect -1480 11150 -1470 11210
rect -1550 11100 -1470 11150
rect -1550 11040 -1540 11100
rect -1480 11040 -1470 11100
rect -1860 11030 -1660 11036
rect -1550 11030 -1470 11040
rect -1000 11160 -990 11400
rect -950 11160 -930 11400
rect -1000 11080 -930 11160
rect -1362 11030 -1162 11036
rect -1970 11000 -1890 11020
rect -1970 10940 -1960 11000
rect -1900 10986 -1890 11000
rect -1860 10996 -1848 11030
rect -1672 11000 -1350 11030
rect -1672 10996 -1660 11000
rect -1860 10990 -1660 10996
rect -1362 10996 -1350 11000
rect -1174 10996 -1162 11030
rect -1362 10990 -1162 10996
rect -1130 11000 -1050 11020
rect -1898 10952 -1890 10986
rect -1900 10940 -1890 10952
rect -1970 10920 -1890 10940
rect -1860 10942 -1660 10948
rect -1860 10908 -1848 10942
rect -1672 10940 -1660 10942
rect -1362 10942 -1162 10948
rect -1362 10940 -1350 10942
rect -1672 10930 -1350 10940
rect -1672 10910 -1540 10930
rect -1672 10908 -1660 10910
rect -1860 10902 -1660 10908
rect -1550 10870 -1540 10910
rect -1480 10910 -1350 10930
rect -1480 10870 -1470 10910
rect -1362 10908 -1350 10910
rect -1174 10908 -1162 10942
rect -1130 10940 -1120 11000
rect -1060 10940 -1050 11000
rect -1130 10920 -1050 10940
rect -1362 10902 -1162 10908
rect -1550 10860 -1470 10870
rect -2080 10150 -2010 10840
rect -1000 10840 -990 11080
rect -950 10840 -930 11080
rect -1000 10430 -930 10840
rect -1020 10390 -930 10400
rect -1020 10330 -1010 10390
rect -940 10330 -930 10390
rect -1020 10320 -930 10330
rect -1000 10260 -930 10320
rect -1010 10250 -930 10260
rect -1010 10190 -1000 10250
rect -940 10190 -930 10250
rect -1010 10180 -930 10190
rect -2080 10140 -930 10150
rect -2080 10080 -2070 10140
rect -2010 10090 -930 10140
rect -2010 10080 -2000 10090
rect -2080 10070 -2000 10080
rect -2080 9690 -2010 10070
rect -2080 9450 -2060 9690
rect -2020 9450 -2010 9690
rect -1000 9690 -930 10090
rect -1550 9670 -1470 9680
rect -1860 9630 -1660 9636
rect -1550 9630 -1540 9670
rect -1970 9600 -1890 9620
rect -1970 9540 -1960 9600
rect -1900 9586 -1890 9600
rect -1860 9596 -1848 9630
rect -1672 9610 -1540 9630
rect -1480 9630 -1470 9670
rect -1362 9630 -1162 9636
rect -1480 9610 -1350 9630
rect -1672 9600 -1350 9610
rect -1672 9596 -1660 9600
rect -1860 9590 -1660 9596
rect -1362 9596 -1350 9600
rect -1174 9596 -1162 9630
rect -1362 9590 -1162 9596
rect -1130 9600 -1050 9620
rect -1898 9552 -1890 9586
rect -1900 9540 -1890 9552
rect -1970 9520 -1890 9540
rect -1860 9542 -1660 9548
rect -1860 9508 -1848 9542
rect -1672 9540 -1660 9542
rect -1362 9542 -1162 9548
rect -1362 9540 -1350 9542
rect -1672 9510 -1350 9540
rect -1672 9508 -1660 9510
rect -1860 9502 -1660 9508
rect -2080 9390 -2010 9450
rect -2080 9130 -2060 9390
rect -2020 9130 -2010 9390
rect -1550 9500 -1470 9510
rect -1362 9508 -1350 9510
rect -1174 9508 -1162 9542
rect -1130 9540 -1120 9600
rect -1060 9540 -1050 9600
rect -1130 9520 -1050 9540
rect -1362 9502 -1162 9508
rect -1550 9440 -1540 9500
rect -1480 9440 -1470 9500
rect -1550 9390 -1470 9440
rect -1550 9330 -1540 9390
rect -1480 9330 -1470 9390
rect -1860 9320 -1660 9326
rect -1550 9320 -1470 9330
rect -1000 9450 -990 9690
rect -950 9450 -930 9690
rect -1000 9370 -930 9450
rect -1362 9320 -1162 9326
rect -1970 9290 -1890 9310
rect -1970 9230 -1960 9290
rect -1900 9276 -1890 9290
rect -1860 9286 -1848 9320
rect -1672 9290 -1350 9320
rect -1672 9286 -1660 9290
rect -1860 9280 -1660 9286
rect -1362 9286 -1350 9290
rect -1174 9286 -1162 9320
rect -1362 9280 -1162 9286
rect -1130 9290 -1050 9310
rect -1898 9242 -1890 9276
rect -1900 9230 -1890 9242
rect -1970 9210 -1890 9230
rect -1860 9232 -1660 9238
rect -1860 9198 -1848 9232
rect -1672 9230 -1660 9232
rect -1362 9232 -1162 9238
rect -1362 9230 -1350 9232
rect -1672 9220 -1350 9230
rect -1672 9200 -1540 9220
rect -1672 9198 -1660 9200
rect -1860 9192 -1660 9198
rect -1550 9160 -1540 9200
rect -1480 9200 -1350 9220
rect -1480 9160 -1470 9200
rect -1362 9198 -1350 9200
rect -1174 9198 -1162 9232
rect -1130 9230 -1120 9290
rect -1060 9230 -1050 9290
rect -1130 9210 -1050 9230
rect -1362 9192 -1162 9198
rect -1550 9150 -1470 9160
rect -2080 8440 -2010 9130
rect -1000 9130 -990 9370
rect -950 9130 -930 9370
rect -1000 8720 -930 9130
rect -1020 8680 -930 8690
rect -1020 8620 -1010 8680
rect -940 8620 -930 8680
rect -1020 8610 -930 8620
rect -1000 8550 -930 8610
rect -1010 8540 -930 8550
rect -1010 8480 -1000 8540
rect -940 8480 -930 8540
rect -1010 8470 -930 8480
rect -2080 8430 -930 8440
rect -2080 8370 -2070 8430
rect -2010 8380 -930 8430
rect -2010 8370 -2000 8380
rect -2080 8360 -2000 8370
rect -2080 7980 -2010 8360
rect -2080 7740 -2060 7980
rect -2020 7740 -2010 7980
rect -1000 7980 -930 8380
rect -1550 7960 -1470 7970
rect -1860 7920 -1660 7926
rect -1550 7920 -1540 7960
rect -1970 7890 -1890 7910
rect -1970 7830 -1960 7890
rect -1900 7876 -1890 7890
rect -1860 7886 -1848 7920
rect -1672 7900 -1540 7920
rect -1480 7920 -1470 7960
rect -1362 7920 -1162 7926
rect -1480 7900 -1350 7920
rect -1672 7890 -1350 7900
rect -1672 7886 -1660 7890
rect -1860 7880 -1660 7886
rect -1362 7886 -1350 7890
rect -1174 7886 -1162 7920
rect -1362 7880 -1162 7886
rect -1130 7890 -1050 7910
rect -1898 7842 -1890 7876
rect -1900 7830 -1890 7842
rect -1970 7810 -1890 7830
rect -1860 7832 -1660 7838
rect -1860 7798 -1848 7832
rect -1672 7830 -1660 7832
rect -1362 7832 -1162 7838
rect -1362 7830 -1350 7832
rect -1672 7800 -1350 7830
rect -1672 7798 -1660 7800
rect -1860 7792 -1660 7798
rect -2080 7680 -2010 7740
rect -2080 7420 -2060 7680
rect -2020 7420 -2010 7680
rect -1550 7790 -1470 7800
rect -1362 7798 -1350 7800
rect -1174 7798 -1162 7832
rect -1130 7830 -1120 7890
rect -1060 7830 -1050 7890
rect -1130 7810 -1050 7830
rect -1362 7792 -1162 7798
rect -1550 7730 -1540 7790
rect -1480 7730 -1470 7790
rect -1550 7680 -1470 7730
rect -1550 7620 -1540 7680
rect -1480 7620 -1470 7680
rect -1860 7610 -1660 7616
rect -1550 7610 -1470 7620
rect -1000 7740 -990 7980
rect -950 7740 -930 7980
rect -1000 7660 -930 7740
rect -1362 7610 -1162 7616
rect -1970 7580 -1890 7600
rect -1970 7520 -1960 7580
rect -1900 7566 -1890 7580
rect -1860 7576 -1848 7610
rect -1672 7580 -1350 7610
rect -1672 7576 -1660 7580
rect -1860 7570 -1660 7576
rect -1362 7576 -1350 7580
rect -1174 7576 -1162 7610
rect -1362 7570 -1162 7576
rect -1130 7580 -1050 7600
rect -1898 7532 -1890 7566
rect -1900 7520 -1890 7532
rect -1970 7500 -1890 7520
rect -1860 7522 -1660 7528
rect -1860 7488 -1848 7522
rect -1672 7520 -1660 7522
rect -1362 7522 -1162 7528
rect -1362 7520 -1350 7522
rect -1672 7510 -1350 7520
rect -1672 7490 -1540 7510
rect -1672 7488 -1660 7490
rect -1860 7482 -1660 7488
rect -1550 7450 -1540 7490
rect -1480 7490 -1350 7510
rect -1480 7450 -1470 7490
rect -1362 7488 -1350 7490
rect -1174 7488 -1162 7522
rect -1130 7520 -1120 7580
rect -1060 7520 -1050 7580
rect -1130 7500 -1050 7520
rect -1362 7482 -1162 7488
rect -1550 7440 -1470 7450
rect -2080 6730 -2010 7420
rect -1000 7420 -990 7660
rect -950 7420 -930 7660
rect -1000 7010 -930 7420
rect -1020 6970 -930 6980
rect -1020 6910 -1010 6970
rect -940 6910 -930 6970
rect -1020 6900 -930 6910
rect -1000 6840 -930 6900
rect -1010 6830 -930 6840
rect -1010 6770 -1000 6830
rect -940 6770 -930 6830
rect -1010 6760 -930 6770
rect -2080 6720 -930 6730
rect -2080 6660 -2070 6720
rect -2010 6670 -930 6720
rect -2010 6660 -2000 6670
rect -2080 6650 -2000 6660
rect -2080 6270 -2010 6650
rect -2080 6030 -2060 6270
rect -2020 6030 -2010 6270
rect -1000 6270 -930 6670
rect -1550 6250 -1470 6260
rect -1860 6210 -1660 6216
rect -1550 6210 -1540 6250
rect -1970 6180 -1890 6200
rect -1970 6120 -1960 6180
rect -1900 6166 -1890 6180
rect -1860 6176 -1848 6210
rect -1672 6190 -1540 6210
rect -1480 6210 -1470 6250
rect -1362 6210 -1162 6216
rect -1480 6190 -1350 6210
rect -1672 6180 -1350 6190
rect -1672 6176 -1660 6180
rect -1860 6170 -1660 6176
rect -1362 6176 -1350 6180
rect -1174 6176 -1162 6210
rect -1362 6170 -1162 6176
rect -1130 6180 -1050 6200
rect -1898 6132 -1890 6166
rect -1900 6120 -1890 6132
rect -1970 6100 -1890 6120
rect -1860 6122 -1660 6128
rect -1860 6088 -1848 6122
rect -1672 6120 -1660 6122
rect -1362 6122 -1162 6128
rect -1362 6120 -1350 6122
rect -1672 6090 -1350 6120
rect -1672 6088 -1660 6090
rect -1860 6082 -1660 6088
rect -2080 5970 -2010 6030
rect -2080 5710 -2060 5970
rect -2020 5710 -2010 5970
rect -1550 6080 -1470 6090
rect -1362 6088 -1350 6090
rect -1174 6088 -1162 6122
rect -1130 6120 -1120 6180
rect -1060 6120 -1050 6180
rect -1130 6100 -1050 6120
rect -1362 6082 -1162 6088
rect -1550 6020 -1540 6080
rect -1480 6020 -1470 6080
rect -1550 5970 -1470 6020
rect -1550 5910 -1540 5970
rect -1480 5910 -1470 5970
rect -1860 5900 -1660 5906
rect -1550 5900 -1470 5910
rect -1000 6030 -990 6270
rect -950 6030 -930 6270
rect -1000 5950 -930 6030
rect -1362 5900 -1162 5906
rect -1970 5870 -1890 5890
rect -1970 5810 -1960 5870
rect -1900 5856 -1890 5870
rect -1860 5866 -1848 5900
rect -1672 5870 -1350 5900
rect -1672 5866 -1660 5870
rect -1860 5860 -1660 5866
rect -1362 5866 -1350 5870
rect -1174 5866 -1162 5900
rect -1362 5860 -1162 5866
rect -1130 5870 -1050 5890
rect -1898 5822 -1890 5856
rect -1900 5810 -1890 5822
rect -1970 5790 -1890 5810
rect -1860 5812 -1660 5818
rect -1860 5778 -1848 5812
rect -1672 5810 -1660 5812
rect -1362 5812 -1162 5818
rect -1362 5810 -1350 5812
rect -1672 5800 -1350 5810
rect -1672 5780 -1540 5800
rect -1672 5778 -1660 5780
rect -1860 5772 -1660 5778
rect -1550 5740 -1540 5780
rect -1480 5780 -1350 5800
rect -1480 5740 -1470 5780
rect -1362 5778 -1350 5780
rect -1174 5778 -1162 5812
rect -1130 5810 -1120 5870
rect -1060 5810 -1050 5870
rect -1130 5790 -1050 5810
rect -1362 5772 -1162 5778
rect -1550 5730 -1470 5740
rect -2080 5020 -2010 5710
rect -1000 5710 -990 5950
rect -950 5710 -930 5950
rect -1000 5300 -930 5710
rect -1020 5260 -930 5270
rect -1020 5200 -1010 5260
rect -940 5200 -930 5260
rect -1020 5190 -930 5200
rect -1000 5130 -930 5190
rect -1010 5120 -930 5130
rect -1010 5060 -1000 5120
rect -940 5060 -930 5120
rect -1010 5050 -930 5060
rect -2080 5010 -930 5020
rect -2080 4950 -2070 5010
rect -2010 4960 -930 5010
rect -2010 4950 -2000 4960
rect -2080 4940 -2000 4950
rect -2080 4560 -2010 4940
rect -2080 4320 -2060 4560
rect -2020 4320 -2010 4560
rect -1000 4560 -930 4960
rect -1550 4540 -1470 4550
rect -1860 4500 -1660 4506
rect -1550 4500 -1540 4540
rect -1970 4470 -1890 4490
rect -1970 4410 -1960 4470
rect -1900 4456 -1890 4470
rect -1860 4466 -1848 4500
rect -1672 4480 -1540 4500
rect -1480 4500 -1470 4540
rect -1362 4500 -1162 4506
rect -1480 4480 -1350 4500
rect -1672 4470 -1350 4480
rect -1672 4466 -1660 4470
rect -1860 4460 -1660 4466
rect -1362 4466 -1350 4470
rect -1174 4466 -1162 4500
rect -1362 4460 -1162 4466
rect -1130 4470 -1050 4490
rect -1898 4422 -1890 4456
rect -1900 4410 -1890 4422
rect -1970 4390 -1890 4410
rect -1860 4412 -1660 4418
rect -1860 4378 -1848 4412
rect -1672 4410 -1660 4412
rect -1362 4412 -1162 4418
rect -1362 4410 -1350 4412
rect -1672 4380 -1350 4410
rect -1672 4378 -1660 4380
rect -1860 4372 -1660 4378
rect -2080 4260 -2010 4320
rect -2080 4000 -2060 4260
rect -2020 4000 -2010 4260
rect -1550 4370 -1470 4380
rect -1362 4378 -1350 4380
rect -1174 4378 -1162 4412
rect -1130 4410 -1120 4470
rect -1060 4410 -1050 4470
rect -1130 4390 -1050 4410
rect -1362 4372 -1162 4378
rect -1550 4310 -1540 4370
rect -1480 4310 -1470 4370
rect -1550 4260 -1470 4310
rect -1550 4200 -1540 4260
rect -1480 4200 -1470 4260
rect -1860 4190 -1660 4196
rect -1550 4190 -1470 4200
rect -1000 4320 -990 4560
rect -950 4320 -930 4560
rect -1000 4240 -930 4320
rect -1362 4190 -1162 4196
rect -1970 4160 -1890 4180
rect -1970 4100 -1960 4160
rect -1900 4146 -1890 4160
rect -1860 4156 -1848 4190
rect -1672 4160 -1350 4190
rect -1672 4156 -1660 4160
rect -1860 4150 -1660 4156
rect -1362 4156 -1350 4160
rect -1174 4156 -1162 4190
rect -1362 4150 -1162 4156
rect -1130 4160 -1050 4180
rect -1898 4112 -1890 4146
rect -1900 4100 -1890 4112
rect -1970 4080 -1890 4100
rect -1860 4102 -1660 4108
rect -1860 4068 -1848 4102
rect -1672 4100 -1660 4102
rect -1362 4102 -1162 4108
rect -1362 4100 -1350 4102
rect -1672 4090 -1350 4100
rect -1672 4070 -1540 4090
rect -1672 4068 -1660 4070
rect -1860 4062 -1660 4068
rect -1550 4030 -1540 4070
rect -1480 4070 -1350 4090
rect -1480 4030 -1470 4070
rect -1362 4068 -1350 4070
rect -1174 4068 -1162 4102
rect -1130 4100 -1120 4160
rect -1060 4100 -1050 4160
rect -1130 4080 -1050 4100
rect -1362 4062 -1162 4068
rect -1550 4020 -1470 4030
rect -2080 3310 -2010 4000
rect -1000 4000 -990 4240
rect -950 4000 -930 4240
rect -1000 3590 -930 4000
rect -1020 3550 -930 3560
rect -1020 3490 -1010 3550
rect -940 3490 -930 3550
rect -1020 3480 -930 3490
rect -1000 3420 -930 3480
rect -1010 3410 -930 3420
rect -1010 3350 -1000 3410
rect -940 3350 -930 3410
rect -1010 3340 -930 3350
rect -2080 3300 -930 3310
rect -2080 3240 -2070 3300
rect -2010 3250 -930 3300
rect -2010 3240 -2000 3250
rect -2080 3230 -2000 3240
rect -2080 2850 -2010 3230
rect -2080 2610 -2060 2850
rect -2020 2610 -2010 2850
rect -1000 2850 -930 3250
rect -1550 2830 -1470 2840
rect -1860 2790 -1660 2796
rect -1550 2790 -1540 2830
rect -1970 2760 -1890 2780
rect -1970 2700 -1960 2760
rect -1900 2746 -1890 2760
rect -1860 2756 -1848 2790
rect -1672 2770 -1540 2790
rect -1480 2790 -1470 2830
rect -1362 2790 -1162 2796
rect -1480 2770 -1350 2790
rect -1672 2760 -1350 2770
rect -1672 2756 -1660 2760
rect -1860 2750 -1660 2756
rect -1362 2756 -1350 2760
rect -1174 2756 -1162 2790
rect -1362 2750 -1162 2756
rect -1130 2760 -1050 2780
rect -1898 2712 -1890 2746
rect -1900 2700 -1890 2712
rect -1970 2680 -1890 2700
rect -1860 2702 -1660 2708
rect -1860 2668 -1848 2702
rect -1672 2700 -1660 2702
rect -1362 2702 -1162 2708
rect -1362 2700 -1350 2702
rect -1672 2670 -1350 2700
rect -1672 2668 -1660 2670
rect -1860 2662 -1660 2668
rect -2080 2550 -2010 2610
rect -2080 2290 -2060 2550
rect -2020 2290 -2010 2550
rect -1550 2660 -1470 2670
rect -1362 2668 -1350 2670
rect -1174 2668 -1162 2702
rect -1130 2700 -1120 2760
rect -1060 2700 -1050 2760
rect -1130 2680 -1050 2700
rect -1362 2662 -1162 2668
rect -1550 2600 -1540 2660
rect -1480 2600 -1470 2660
rect -1550 2550 -1470 2600
rect -1550 2490 -1540 2550
rect -1480 2490 -1470 2550
rect -1860 2480 -1660 2486
rect -1550 2480 -1470 2490
rect -1000 2610 -990 2850
rect -950 2610 -930 2850
rect -1000 2530 -930 2610
rect -1362 2480 -1162 2486
rect -1970 2450 -1890 2470
rect -1970 2390 -1960 2450
rect -1900 2436 -1890 2450
rect -1860 2446 -1848 2480
rect -1672 2450 -1350 2480
rect -1672 2446 -1660 2450
rect -1860 2440 -1660 2446
rect -1362 2446 -1350 2450
rect -1174 2446 -1162 2480
rect -1362 2440 -1162 2446
rect -1130 2450 -1050 2470
rect -1898 2402 -1890 2436
rect -1900 2390 -1890 2402
rect -1970 2370 -1890 2390
rect -1860 2392 -1660 2398
rect -1860 2358 -1848 2392
rect -1672 2390 -1660 2392
rect -1362 2392 -1162 2398
rect -1362 2390 -1350 2392
rect -1672 2380 -1350 2390
rect -1672 2360 -1540 2380
rect -1672 2358 -1660 2360
rect -1860 2352 -1660 2358
rect -1550 2320 -1540 2360
rect -1480 2360 -1350 2380
rect -1480 2320 -1470 2360
rect -1362 2358 -1350 2360
rect -1174 2358 -1162 2392
rect -1130 2390 -1120 2450
rect -1060 2390 -1050 2450
rect -1130 2370 -1050 2390
rect -1362 2352 -1162 2358
rect -1550 2310 -1470 2320
rect -2080 1600 -2010 2290
rect -1000 2290 -990 2530
rect -950 2290 -930 2530
rect -1000 1880 -930 2290
rect -1020 1840 -930 1850
rect -1020 1780 -1010 1840
rect -940 1780 -930 1840
rect -1020 1770 -930 1780
rect -1000 1710 -930 1770
rect -1010 1700 -930 1710
rect -1010 1640 -1000 1700
rect -940 1640 -930 1700
rect -1010 1630 -930 1640
rect -2080 1590 -930 1600
rect -2080 1530 -2070 1590
rect -2010 1540 -930 1590
rect -2010 1530 -2000 1540
rect -2080 1520 -2000 1530
rect -2080 1140 -2010 1520
rect -2080 900 -2060 1140
rect -2020 900 -2010 1140
rect -1000 1140 -930 1540
rect -1550 1120 -1470 1130
rect -1860 1080 -1660 1086
rect -1550 1080 -1540 1120
rect -1970 1050 -1890 1070
rect -1970 990 -1960 1050
rect -1900 1036 -1890 1050
rect -1860 1046 -1848 1080
rect -1672 1060 -1540 1080
rect -1480 1080 -1470 1120
rect -1362 1080 -1162 1086
rect -1480 1060 -1350 1080
rect -1672 1050 -1350 1060
rect -1672 1046 -1660 1050
rect -1860 1040 -1660 1046
rect -1362 1046 -1350 1050
rect -1174 1046 -1162 1080
rect -1362 1040 -1162 1046
rect -1130 1050 -1050 1070
rect -1898 1002 -1890 1036
rect -1900 990 -1890 1002
rect -1970 970 -1890 990
rect -1860 992 -1660 998
rect -1860 958 -1848 992
rect -1672 990 -1660 992
rect -1362 992 -1162 998
rect -1362 990 -1350 992
rect -1672 960 -1350 990
rect -1672 958 -1660 960
rect -1860 952 -1660 958
rect -2080 840 -2010 900
rect -2080 580 -2060 840
rect -2020 580 -2010 840
rect -1550 950 -1470 960
rect -1362 958 -1350 960
rect -1174 958 -1162 992
rect -1130 990 -1120 1050
rect -1060 990 -1050 1050
rect -1130 970 -1050 990
rect -1362 952 -1162 958
rect -1550 890 -1540 950
rect -1480 890 -1470 950
rect -1550 840 -1470 890
rect -1550 780 -1540 840
rect -1480 780 -1470 840
rect -1860 770 -1660 776
rect -1550 770 -1470 780
rect -1000 900 -990 1140
rect -950 900 -930 1140
rect -1000 820 -930 900
rect -1362 770 -1162 776
rect -1970 740 -1890 760
rect -1970 680 -1960 740
rect -1900 726 -1890 740
rect -1860 736 -1848 770
rect -1672 740 -1350 770
rect -1672 736 -1660 740
rect -1860 730 -1660 736
rect -1362 736 -1350 740
rect -1174 736 -1162 770
rect -1362 730 -1162 736
rect -1130 740 -1050 760
rect -1898 692 -1890 726
rect -1900 680 -1890 692
rect -1970 660 -1890 680
rect -1860 682 -1660 688
rect -1860 648 -1848 682
rect -1672 680 -1660 682
rect -1362 682 -1162 688
rect -1362 680 -1350 682
rect -1672 670 -1350 680
rect -1672 650 -1540 670
rect -1672 648 -1660 650
rect -1860 642 -1660 648
rect -1550 610 -1540 650
rect -1480 650 -1350 670
rect -1480 610 -1470 650
rect -1362 648 -1350 650
rect -1174 648 -1162 682
rect -1130 680 -1120 740
rect -1060 680 -1050 740
rect -1130 660 -1050 680
rect -1362 642 -1162 648
rect -1550 600 -1470 610
rect -2080 150 -2010 580
rect -1000 580 -990 820
rect -950 580 -930 820
rect -1000 170 -930 580
rect -2080 140 -2000 150
rect -900 140 -870 23940
rect -810 140 -780 23940
rect -750 140 -720 23940
rect -630 140 -600 23940
rect -510 140 -480 23940
rect -390 140 -360 23940
rect -270 140 -240 23940
rect -150 140 -120 23940
rect -30 140 0 23940
rect -2080 80 -2070 140
rect -2010 80 -2000 140
rect -2080 70 -2000 80
rect -1020 130 -930 140
rect -1020 70 -1010 130
rect -940 70 -930 130
rect -2080 -110 -2010 70
rect -1020 60 -930 70
rect -1000 0 -930 60
rect -1010 -10 -930 0
rect -1010 -70 -1000 -10
rect -940 -70 -930 -10
rect -1010 -80 -930 -70
rect -2080 -120 -930 -110
rect -2080 -180 -2070 -120
rect -2010 -170 -930 -120
rect -2010 -180 -2000 -170
rect -2080 -190 -2000 -180
rect -2080 -570 -2010 -190
rect -2080 -810 -2060 -570
rect -2020 -810 -2010 -570
rect -1000 -570 -930 -170
rect -1550 -590 -1470 -580
rect -1860 -630 -1660 -624
rect -1550 -630 -1540 -590
rect -1970 -660 -1890 -640
rect -1970 -720 -1960 -660
rect -1900 -674 -1890 -660
rect -1860 -664 -1848 -630
rect -1672 -650 -1540 -630
rect -1480 -630 -1470 -590
rect -1362 -630 -1162 -624
rect -1480 -650 -1350 -630
rect -1672 -660 -1350 -650
rect -1672 -664 -1660 -660
rect -1860 -670 -1660 -664
rect -1362 -664 -1350 -660
rect -1174 -664 -1162 -630
rect -1362 -670 -1162 -664
rect -1130 -660 -1050 -640
rect -1898 -708 -1890 -674
rect -1900 -720 -1890 -708
rect -1970 -740 -1890 -720
rect -1860 -718 -1660 -712
rect -1860 -752 -1848 -718
rect -1672 -720 -1660 -718
rect -1362 -718 -1162 -712
rect -1362 -720 -1350 -718
rect -1672 -750 -1350 -720
rect -1672 -752 -1660 -750
rect -1860 -758 -1660 -752
rect -2080 -870 -2010 -810
rect -2080 -1130 -2060 -870
rect -2020 -1130 -2010 -870
rect -1550 -760 -1470 -750
rect -1362 -752 -1350 -750
rect -1174 -752 -1162 -718
rect -1130 -720 -1120 -660
rect -1060 -720 -1050 -660
rect -1130 -740 -1050 -720
rect -1362 -758 -1162 -752
rect -1550 -820 -1540 -760
rect -1480 -820 -1470 -760
rect -1550 -870 -1470 -820
rect -1550 -930 -1540 -870
rect -1480 -930 -1470 -870
rect -1860 -940 -1660 -934
rect -1550 -940 -1470 -930
rect -1000 -810 -990 -570
rect -950 -810 -930 -570
rect -1000 -890 -930 -810
rect -1362 -940 -1162 -934
rect -1970 -970 -1890 -950
rect -1970 -1030 -1960 -970
rect -1900 -984 -1890 -970
rect -1860 -974 -1848 -940
rect -1672 -970 -1350 -940
rect -1672 -974 -1660 -970
rect -1860 -980 -1660 -974
rect -1362 -974 -1350 -970
rect -1174 -974 -1162 -940
rect -1362 -980 -1162 -974
rect -1130 -970 -1050 -950
rect -1898 -1018 -1890 -984
rect -1900 -1030 -1890 -1018
rect -1970 -1050 -1890 -1030
rect -1860 -1028 -1660 -1022
rect -1860 -1062 -1848 -1028
rect -1672 -1030 -1660 -1028
rect -1362 -1028 -1162 -1022
rect -1362 -1030 -1350 -1028
rect -1672 -1040 -1350 -1030
rect -1672 -1060 -1540 -1040
rect -1672 -1062 -1660 -1060
rect -1860 -1068 -1660 -1062
rect -1550 -1100 -1540 -1060
rect -1480 -1060 -1350 -1040
rect -1480 -1100 -1470 -1060
rect -1362 -1062 -1350 -1060
rect -1174 -1062 -1162 -1028
rect -1130 -1030 -1120 -970
rect -1060 -1030 -1050 -970
rect -1130 -1050 -1050 -1030
rect -1362 -1068 -1162 -1062
rect -1550 -1110 -1470 -1100
rect -2080 -1710 -2010 -1130
rect -1000 -1130 -990 -890
rect -950 -1130 -930 -890
rect -1000 -1540 -930 -1130
rect -1020 -1580 -930 -1570
rect -1020 -1640 -1010 -1580
rect -940 -1640 -930 -1580
rect -1020 -1650 -930 -1640
rect -1000 -1710 -930 -1650
rect -900 -1710 -870 -110
rect -810 -1710 -780 -110
rect -750 -1710 -720 -110
rect -630 -1710 -600 -110
rect -510 -1710 -480 -110
rect -390 -1710 -360 -110
rect -270 -1710 -240 -110
rect -150 -1710 -120 -110
rect -30 -1710 0 -110
rect 1860 -1710 1890 150
rect 1980 -1710 2010 150
rect 2100 -1710 2130 150
rect 2220 -1710 2250 150
rect 2340 -1710 2370 150
rect 2460 -1710 2490 150
rect 2580 -1710 2610 150
rect 2640 140 2720 150
rect 2640 80 2650 140
rect 2710 80 2720 140
rect 2640 70 2720 80
rect 2640 -110 2710 70
rect 2640 -120 3790 -110
rect 2640 -180 2650 -120
rect 2710 -170 3790 -120
rect 2710 -180 2720 -170
rect 2640 -190 2720 -180
rect 2640 -570 2710 -190
rect 2640 -810 2660 -570
rect 2700 -810 2710 -570
rect 3720 -570 3790 -170
rect 3170 -590 3250 -580
rect 2860 -630 3060 -624
rect 3170 -630 3180 -590
rect 2750 -660 2830 -640
rect 2750 -720 2760 -660
rect 2820 -674 2830 -660
rect 2860 -664 2872 -630
rect 3048 -650 3180 -630
rect 3240 -630 3250 -590
rect 3358 -630 3558 -624
rect 3240 -650 3370 -630
rect 3048 -660 3370 -650
rect 3048 -664 3060 -660
rect 2860 -670 3060 -664
rect 3358 -664 3370 -660
rect 3546 -664 3558 -630
rect 3358 -670 3558 -664
rect 3590 -660 3670 -640
rect 2822 -708 2830 -674
rect 2820 -720 2830 -708
rect 2750 -740 2830 -720
rect 2860 -718 3060 -712
rect 2860 -752 2872 -718
rect 3048 -720 3060 -718
rect 3358 -718 3558 -712
rect 3358 -720 3370 -718
rect 3048 -750 3370 -720
rect 3048 -752 3060 -750
rect 2860 -758 3060 -752
rect 2640 -870 2710 -810
rect 2640 -1130 2660 -870
rect 2700 -1130 2710 -870
rect 3170 -760 3250 -750
rect 3358 -752 3370 -750
rect 3546 -752 3558 -718
rect 3590 -720 3600 -660
rect 3660 -720 3670 -660
rect 3590 -740 3670 -720
rect 3358 -758 3558 -752
rect 3170 -820 3180 -760
rect 3240 -820 3250 -760
rect 3170 -870 3250 -820
rect 3170 -930 3180 -870
rect 3240 -930 3250 -870
rect 2860 -940 3060 -934
rect 3170 -940 3250 -930
rect 3720 -810 3730 -570
rect 3770 -810 3790 -570
rect 3720 -890 3790 -810
rect 3358 -940 3558 -934
rect 2750 -970 2830 -950
rect 2750 -1030 2760 -970
rect 2820 -984 2830 -970
rect 2860 -974 2872 -940
rect 3048 -970 3370 -940
rect 3048 -974 3060 -970
rect 2860 -980 3060 -974
rect 3358 -974 3370 -970
rect 3546 -974 3558 -940
rect 3358 -980 3558 -974
rect 3590 -970 3670 -950
rect 2822 -1018 2830 -984
rect 2820 -1030 2830 -1018
rect 2750 -1050 2830 -1030
rect 2860 -1028 3060 -1022
rect 2860 -1062 2872 -1028
rect 3048 -1030 3060 -1028
rect 3358 -1028 3558 -1022
rect 3358 -1030 3370 -1028
rect 3048 -1040 3370 -1030
rect 3048 -1060 3180 -1040
rect 3048 -1062 3060 -1060
rect 2860 -1068 3060 -1062
rect 3170 -1100 3180 -1060
rect 3240 -1060 3370 -1040
rect 3240 -1100 3250 -1060
rect 3358 -1062 3370 -1060
rect 3546 -1062 3558 -1028
rect 3590 -1030 3600 -970
rect 3660 -1030 3670 -970
rect 3590 -1050 3670 -1030
rect 3358 -1068 3558 -1062
rect 3170 -1110 3250 -1100
rect 2640 -1710 2710 -1130
rect 3720 -1130 3730 -890
rect 3770 -1130 3790 -890
rect 3720 -1600 3790 -1130
rect 3710 -1640 3790 -1630
rect 3710 -1700 3720 -1640
rect 3780 -1700 3790 -1640
rect 3710 -1710 3790 -1700
rect 3820 -1710 3850 0
rect 3910 -1710 3940 0
rect 3970 -1710 4000 0
rect 4090 -1710 4120 0
rect 4210 -1710 4240 0
rect 4330 -1710 4360 0
rect 4450 -1710 4480 0
rect 4570 -1710 4600 0
rect 4690 -1710 4720 0
rect 6850 -1710 6880 150
rect 6970 -1710 7000 150
rect 7090 -1710 7120 150
rect 7210 -1710 7240 150
rect 7330 -1710 7360 150
rect 7450 -1710 7480 150
rect 7570 -1710 7600 150
rect 7630 140 7710 150
rect 7630 80 7640 140
rect 7700 80 7710 140
rect 7630 70 7710 80
rect 7630 -110 7700 70
rect 8710 0 8780 130
rect 7630 -120 8780 -110
rect 7630 -180 7640 -120
rect 7700 -170 8780 -120
rect 7700 -180 7710 -170
rect 7630 -190 7710 -180
rect 7630 -570 7700 -190
rect 7630 -810 7650 -570
rect 7690 -810 7700 -570
rect 8710 -570 8780 -170
rect 8160 -590 8240 -580
rect 7850 -630 8050 -624
rect 8160 -630 8170 -590
rect 7740 -660 7820 -640
rect 7740 -720 7750 -660
rect 7810 -674 7820 -660
rect 7850 -664 7862 -630
rect 8038 -650 8170 -630
rect 8230 -630 8240 -590
rect 8348 -630 8548 -624
rect 8230 -650 8360 -630
rect 8038 -660 8360 -650
rect 8038 -664 8050 -660
rect 7850 -670 8050 -664
rect 8348 -664 8360 -660
rect 8536 -664 8548 -630
rect 8348 -670 8548 -664
rect 8580 -660 8660 -640
rect 7812 -708 7820 -674
rect 7810 -720 7820 -708
rect 7740 -740 7820 -720
rect 7850 -718 8050 -712
rect 7850 -752 7862 -718
rect 8038 -720 8050 -718
rect 8348 -718 8548 -712
rect 8348 -720 8360 -718
rect 8038 -750 8360 -720
rect 8038 -752 8050 -750
rect 7850 -758 8050 -752
rect 7630 -870 7700 -810
rect 7630 -1130 7650 -870
rect 7690 -1130 7700 -870
rect 8160 -760 8240 -750
rect 8348 -752 8360 -750
rect 8536 -752 8548 -718
rect 8580 -720 8590 -660
rect 8650 -720 8660 -660
rect 8580 -740 8660 -720
rect 8348 -758 8548 -752
rect 8160 -820 8170 -760
rect 8230 -820 8240 -760
rect 8160 -870 8240 -820
rect 8160 -930 8170 -870
rect 8230 -930 8240 -870
rect 7850 -940 8050 -934
rect 8160 -940 8240 -930
rect 8710 -810 8720 -570
rect 8760 -810 8780 -570
rect 8710 -890 8780 -810
rect 8348 -940 8548 -934
rect 7740 -970 7820 -950
rect 7740 -1030 7750 -970
rect 7810 -984 7820 -970
rect 7850 -974 7862 -940
rect 8038 -970 8360 -940
rect 8038 -974 8050 -970
rect 7850 -980 8050 -974
rect 8348 -974 8360 -970
rect 8536 -974 8548 -940
rect 8348 -980 8548 -974
rect 8580 -970 8660 -950
rect 7812 -1018 7820 -984
rect 7810 -1030 7820 -1018
rect 7740 -1050 7820 -1030
rect 7850 -1028 8050 -1022
rect 7850 -1062 7862 -1028
rect 8038 -1030 8050 -1028
rect 8348 -1028 8548 -1022
rect 8348 -1030 8360 -1028
rect 8038 -1040 8360 -1030
rect 8038 -1060 8170 -1040
rect 8038 -1062 8050 -1060
rect 7850 -1068 8050 -1062
rect 8160 -1100 8170 -1060
rect 8230 -1060 8360 -1040
rect 8230 -1100 8240 -1060
rect 8348 -1062 8360 -1060
rect 8536 -1062 8548 -1028
rect 8580 -1030 8590 -970
rect 8650 -1030 8660 -970
rect 8580 -1050 8660 -1030
rect 8348 -1068 8548 -1062
rect 8160 -1110 8240 -1100
rect 7630 -1710 7700 -1130
rect 8710 -1130 8720 -890
rect 8760 -1130 8780 -890
rect 8710 -1600 8780 -1130
rect 8700 -1640 8780 -1630
rect 8700 -1700 8710 -1640
rect 8770 -1700 8780 -1640
rect 8700 -1710 8780 -1700
rect 8810 -1710 8840 130
rect 8900 -1710 8930 130
rect 8960 -1710 8990 130
rect 9080 -1710 9110 130
rect 9200 -1710 9230 130
rect 9320 -1710 9350 130
rect 9440 -1710 9470 130
rect 9560 -1710 9590 130
rect 9680 -1710 9710 130
rect 11840 -1710 11870 150
rect 11960 -1710 11990 150
rect 12080 -1710 12110 150
rect 12200 -1710 12230 150
rect 12320 -1710 12350 150
rect 12440 -1710 12470 150
rect 12560 -1710 12590 150
rect 12620 140 12700 150
rect 12620 80 12630 140
rect 12690 80 12700 140
rect 12620 70 12700 80
rect 12620 -110 12690 70
rect 13700 0 13770 130
rect 12620 -120 13770 -110
rect 12620 -180 12630 -120
rect 12690 -170 13770 -120
rect 12690 -180 12700 -170
rect 12620 -190 12700 -180
rect 12620 -570 12690 -190
rect 12620 -810 12640 -570
rect 12680 -810 12690 -570
rect 13700 -570 13770 -170
rect 13150 -590 13230 -580
rect 12840 -630 13040 -624
rect 13150 -630 13160 -590
rect 12730 -660 12810 -640
rect 12730 -720 12740 -660
rect 12800 -674 12810 -660
rect 12840 -664 12852 -630
rect 13028 -650 13160 -630
rect 13220 -630 13230 -590
rect 13338 -630 13538 -624
rect 13220 -650 13350 -630
rect 13028 -660 13350 -650
rect 13028 -664 13040 -660
rect 12840 -670 13040 -664
rect 13338 -664 13350 -660
rect 13526 -664 13538 -630
rect 13338 -670 13538 -664
rect 13570 -660 13650 -640
rect 12802 -708 12810 -674
rect 12800 -720 12810 -708
rect 12730 -740 12810 -720
rect 12840 -718 13040 -712
rect 12840 -752 12852 -718
rect 13028 -720 13040 -718
rect 13338 -718 13538 -712
rect 13338 -720 13350 -718
rect 13028 -750 13350 -720
rect 13028 -752 13040 -750
rect 12840 -758 13040 -752
rect 12620 -870 12690 -810
rect 12620 -1130 12640 -870
rect 12680 -1130 12690 -870
rect 13150 -760 13230 -750
rect 13338 -752 13350 -750
rect 13526 -752 13538 -718
rect 13570 -720 13580 -660
rect 13640 -720 13650 -660
rect 13570 -740 13650 -720
rect 13338 -758 13538 -752
rect 13150 -820 13160 -760
rect 13220 -820 13230 -760
rect 13150 -870 13230 -820
rect 13150 -930 13160 -870
rect 13220 -930 13230 -870
rect 12840 -940 13040 -934
rect 13150 -940 13230 -930
rect 13700 -810 13710 -570
rect 13750 -810 13770 -570
rect 13700 -890 13770 -810
rect 13338 -940 13538 -934
rect 12730 -970 12810 -950
rect 12730 -1030 12740 -970
rect 12800 -984 12810 -970
rect 12840 -974 12852 -940
rect 13028 -970 13350 -940
rect 13028 -974 13040 -970
rect 12840 -980 13040 -974
rect 13338 -974 13350 -970
rect 13526 -974 13538 -940
rect 13338 -980 13538 -974
rect 13570 -970 13650 -950
rect 12802 -1018 12810 -984
rect 12800 -1030 12810 -1018
rect 12730 -1050 12810 -1030
rect 12840 -1028 13040 -1022
rect 12840 -1062 12852 -1028
rect 13028 -1030 13040 -1028
rect 13338 -1028 13538 -1022
rect 13338 -1030 13350 -1028
rect 13028 -1040 13350 -1030
rect 13028 -1060 13160 -1040
rect 13028 -1062 13040 -1060
rect 12840 -1068 13040 -1062
rect 13150 -1100 13160 -1060
rect 13220 -1060 13350 -1040
rect 13220 -1100 13230 -1060
rect 13338 -1062 13350 -1060
rect 13526 -1062 13538 -1028
rect 13570 -1030 13580 -970
rect 13640 -1030 13650 -970
rect 13570 -1050 13650 -1030
rect 13338 -1068 13538 -1062
rect 13150 -1110 13230 -1100
rect 12620 -1710 12690 -1130
rect 13700 -1130 13710 -890
rect 13750 -1130 13770 -890
rect 13700 -1600 13770 -1130
rect 13690 -1640 13770 -1630
rect 13690 -1700 13700 -1640
rect 13760 -1700 13770 -1640
rect 13690 -1710 13770 -1700
rect 13800 -1710 13830 130
rect 13890 -1710 13920 130
rect 13950 -1710 13980 130
rect 14070 -1710 14100 130
rect 14190 -1710 14220 130
rect 14310 -1710 14340 130
rect 14430 -1710 14460 130
rect 14550 -1710 14580 130
rect 14670 -1710 14700 130
rect 16830 -1710 16860 150
rect 16950 -1710 16980 150
rect 17070 -1710 17100 150
rect 17190 -1710 17220 150
rect 17310 -1710 17340 150
rect 17430 -1710 17460 150
rect 17550 -1710 17580 150
rect 17610 140 17690 150
rect 17610 80 17620 140
rect 17680 80 17690 140
rect 17610 70 17690 80
rect 17610 -110 17680 70
rect 18690 0 18760 130
rect 17610 -120 18760 -110
rect 17610 -180 17620 -120
rect 17680 -170 18760 -120
rect 17680 -180 17690 -170
rect 17610 -190 17690 -180
rect 17610 -570 17680 -190
rect 17610 -810 17630 -570
rect 17670 -810 17680 -570
rect 18690 -570 18760 -170
rect 18140 -590 18220 -580
rect 17830 -630 18030 -624
rect 18140 -630 18150 -590
rect 17720 -660 17800 -640
rect 17720 -720 17730 -660
rect 17790 -674 17800 -660
rect 17830 -664 17842 -630
rect 18018 -650 18150 -630
rect 18210 -630 18220 -590
rect 18328 -630 18528 -624
rect 18210 -650 18340 -630
rect 18018 -660 18340 -650
rect 18018 -664 18030 -660
rect 17830 -670 18030 -664
rect 18328 -664 18340 -660
rect 18516 -664 18528 -630
rect 18328 -670 18528 -664
rect 18560 -660 18640 -640
rect 17792 -708 17800 -674
rect 17790 -720 17800 -708
rect 17720 -740 17800 -720
rect 17830 -718 18030 -712
rect 17830 -752 17842 -718
rect 18018 -720 18030 -718
rect 18328 -718 18528 -712
rect 18328 -720 18340 -718
rect 18018 -750 18340 -720
rect 18018 -752 18030 -750
rect 17830 -758 18030 -752
rect 17610 -870 17680 -810
rect 17610 -1130 17630 -870
rect 17670 -1130 17680 -870
rect 18140 -760 18220 -750
rect 18328 -752 18340 -750
rect 18516 -752 18528 -718
rect 18560 -720 18570 -660
rect 18630 -720 18640 -660
rect 18560 -740 18640 -720
rect 18328 -758 18528 -752
rect 18140 -820 18150 -760
rect 18210 -820 18220 -760
rect 18140 -870 18220 -820
rect 18140 -930 18150 -870
rect 18210 -930 18220 -870
rect 17830 -940 18030 -934
rect 18140 -940 18220 -930
rect 18690 -810 18700 -570
rect 18740 -810 18760 -570
rect 18690 -890 18760 -810
rect 18328 -940 18528 -934
rect 17720 -970 17800 -950
rect 17720 -1030 17730 -970
rect 17790 -984 17800 -970
rect 17830 -974 17842 -940
rect 18018 -970 18340 -940
rect 18018 -974 18030 -970
rect 17830 -980 18030 -974
rect 18328 -974 18340 -970
rect 18516 -974 18528 -940
rect 18328 -980 18528 -974
rect 18560 -970 18640 -950
rect 17792 -1018 17800 -984
rect 17790 -1030 17800 -1018
rect 17720 -1050 17800 -1030
rect 17830 -1028 18030 -1022
rect 17830 -1062 17842 -1028
rect 18018 -1030 18030 -1028
rect 18328 -1028 18528 -1022
rect 18328 -1030 18340 -1028
rect 18018 -1040 18340 -1030
rect 18018 -1060 18150 -1040
rect 18018 -1062 18030 -1060
rect 17830 -1068 18030 -1062
rect 18140 -1100 18150 -1060
rect 18210 -1060 18340 -1040
rect 18210 -1100 18220 -1060
rect 18328 -1062 18340 -1060
rect 18516 -1062 18528 -1028
rect 18560 -1030 18570 -970
rect 18630 -1030 18640 -970
rect 18560 -1050 18640 -1030
rect 18328 -1068 18528 -1062
rect 18140 -1110 18220 -1100
rect 17610 -1710 17680 -1130
rect 18690 -1130 18700 -890
rect 18740 -1130 18760 -890
rect 18690 -1600 18760 -1130
rect 18680 -1640 18760 -1630
rect 18680 -1700 18690 -1640
rect 18750 -1700 18760 -1640
rect 18680 -1710 18760 -1700
rect 18790 -1710 18820 130
rect 18880 -1710 18910 130
rect 18940 -1710 18970 130
rect 19060 -1710 19090 130
rect 19180 -1710 19210 130
rect 19300 -1710 19330 130
rect 19420 -1710 19450 130
rect 19540 -1710 19570 130
rect 19660 -1710 19690 130
rect 21820 -1710 21850 150
rect 21940 -1710 21970 150
rect 22060 -1710 22090 150
rect 22180 -1710 22210 150
rect 22300 -1710 22330 150
rect 22420 -1710 22450 150
rect 22540 -1710 22570 150
rect 22600 140 22680 150
rect 22600 80 22610 140
rect 22670 80 22680 140
rect 22600 70 22680 80
rect 22600 -110 22670 70
rect 23680 0 23750 130
rect 22600 -120 23750 -110
rect 22600 -180 22610 -120
rect 22670 -170 23750 -120
rect 22670 -180 22680 -170
rect 22600 -190 22680 -180
rect 22600 -570 22670 -190
rect 22600 -810 22620 -570
rect 22660 -810 22670 -570
rect 23680 -570 23750 -170
rect 23130 -590 23210 -580
rect 22820 -630 23020 -624
rect 23130 -630 23140 -590
rect 22710 -660 22790 -640
rect 22710 -720 22720 -660
rect 22780 -674 22790 -660
rect 22820 -664 22832 -630
rect 23008 -650 23140 -630
rect 23200 -630 23210 -590
rect 23318 -630 23518 -624
rect 23200 -650 23330 -630
rect 23008 -660 23330 -650
rect 23008 -664 23020 -660
rect 22820 -670 23020 -664
rect 23318 -664 23330 -660
rect 23506 -664 23518 -630
rect 23318 -670 23518 -664
rect 23550 -660 23630 -640
rect 22782 -708 22790 -674
rect 22780 -720 22790 -708
rect 22710 -740 22790 -720
rect 22820 -718 23020 -712
rect 22820 -752 22832 -718
rect 23008 -720 23020 -718
rect 23318 -718 23518 -712
rect 23318 -720 23330 -718
rect 23008 -750 23330 -720
rect 23008 -752 23020 -750
rect 22820 -758 23020 -752
rect 22600 -870 22670 -810
rect 22600 -1130 22620 -870
rect 22660 -1130 22670 -870
rect 23130 -760 23210 -750
rect 23318 -752 23330 -750
rect 23506 -752 23518 -718
rect 23550 -720 23560 -660
rect 23620 -720 23630 -660
rect 23550 -740 23630 -720
rect 23318 -758 23518 -752
rect 23130 -820 23140 -760
rect 23200 -820 23210 -760
rect 23130 -870 23210 -820
rect 23130 -930 23140 -870
rect 23200 -930 23210 -870
rect 22820 -940 23020 -934
rect 23130 -940 23210 -930
rect 23680 -810 23690 -570
rect 23730 -810 23750 -570
rect 23680 -890 23750 -810
rect 23318 -940 23518 -934
rect 22710 -970 22790 -950
rect 22710 -1030 22720 -970
rect 22780 -984 22790 -970
rect 22820 -974 22832 -940
rect 23008 -970 23330 -940
rect 23008 -974 23020 -970
rect 22820 -980 23020 -974
rect 23318 -974 23330 -970
rect 23506 -974 23518 -940
rect 23318 -980 23518 -974
rect 23550 -970 23630 -950
rect 22782 -1018 22790 -984
rect 22780 -1030 22790 -1018
rect 22710 -1050 22790 -1030
rect 22820 -1028 23020 -1022
rect 22820 -1062 22832 -1028
rect 23008 -1030 23020 -1028
rect 23318 -1028 23518 -1022
rect 23318 -1030 23330 -1028
rect 23008 -1040 23330 -1030
rect 23008 -1060 23140 -1040
rect 23008 -1062 23020 -1060
rect 22820 -1068 23020 -1062
rect 23130 -1100 23140 -1060
rect 23200 -1060 23330 -1040
rect 23200 -1100 23210 -1060
rect 23318 -1062 23330 -1060
rect 23506 -1062 23518 -1028
rect 23550 -1030 23560 -970
rect 23620 -1030 23630 -970
rect 23550 -1050 23630 -1030
rect 23318 -1068 23518 -1062
rect 23130 -1110 23210 -1100
rect 22600 -1710 22670 -1130
rect 23680 -1130 23690 -890
rect 23730 -1130 23750 -890
rect 23680 -1600 23750 -1130
rect 23670 -1640 23750 -1630
rect 23670 -1700 23680 -1640
rect 23740 -1700 23750 -1640
rect 23670 -1710 23750 -1700
rect 23780 -1710 23810 130
rect 23870 -1710 23900 130
rect 23930 -1710 23960 130
rect 24050 -1710 24080 130
rect 24170 -1710 24200 130
rect 24290 -1710 24320 130
rect 24410 -1710 24440 130
rect 24530 -1710 24560 130
rect 24650 -1710 24680 130
rect 26810 -1710 26840 150
rect 26930 -1710 26960 150
rect 27050 -1710 27080 150
rect 27170 -1710 27200 150
rect 27290 -1710 27320 150
rect 27410 -1710 27440 150
rect 27530 -1710 27560 150
rect 27590 140 27670 150
rect 27590 80 27600 140
rect 27660 80 27670 140
rect 27590 70 27670 80
rect 27590 -110 27660 70
rect 28670 0 28740 130
rect 27590 -120 28740 -110
rect 27590 -180 27600 -120
rect 27660 -170 28740 -120
rect 27660 -180 27670 -170
rect 27590 -190 27670 -180
rect 27590 -570 27660 -190
rect 27590 -810 27610 -570
rect 27650 -810 27660 -570
rect 28670 -570 28740 -170
rect 28120 -590 28200 -580
rect 27810 -630 28010 -624
rect 28120 -630 28130 -590
rect 27700 -660 27780 -640
rect 27700 -720 27710 -660
rect 27770 -674 27780 -660
rect 27810 -664 27822 -630
rect 27998 -650 28130 -630
rect 28190 -630 28200 -590
rect 28308 -630 28508 -624
rect 28190 -650 28320 -630
rect 27998 -660 28320 -650
rect 27998 -664 28010 -660
rect 27810 -670 28010 -664
rect 28308 -664 28320 -660
rect 28496 -664 28508 -630
rect 28308 -670 28508 -664
rect 28540 -660 28620 -640
rect 27772 -708 27780 -674
rect 27770 -720 27780 -708
rect 27700 -740 27780 -720
rect 27810 -718 28010 -712
rect 27810 -752 27822 -718
rect 27998 -720 28010 -718
rect 28308 -718 28508 -712
rect 28308 -720 28320 -718
rect 27998 -750 28320 -720
rect 27998 -752 28010 -750
rect 27810 -758 28010 -752
rect 27590 -870 27660 -810
rect 27590 -1130 27610 -870
rect 27650 -1130 27660 -870
rect 28120 -760 28200 -750
rect 28308 -752 28320 -750
rect 28496 -752 28508 -718
rect 28540 -720 28550 -660
rect 28610 -720 28620 -660
rect 28540 -740 28620 -720
rect 28308 -758 28508 -752
rect 28120 -820 28130 -760
rect 28190 -820 28200 -760
rect 28120 -870 28200 -820
rect 28120 -930 28130 -870
rect 28190 -930 28200 -870
rect 27810 -940 28010 -934
rect 28120 -940 28200 -930
rect 28670 -810 28680 -570
rect 28720 -810 28740 -570
rect 28670 -890 28740 -810
rect 28308 -940 28508 -934
rect 27700 -970 27780 -950
rect 27700 -1030 27710 -970
rect 27770 -984 27780 -970
rect 27810 -974 27822 -940
rect 27998 -970 28320 -940
rect 27998 -974 28010 -970
rect 27810 -980 28010 -974
rect 28308 -974 28320 -970
rect 28496 -974 28508 -940
rect 28308 -980 28508 -974
rect 28540 -970 28620 -950
rect 27772 -1018 27780 -984
rect 27770 -1030 27780 -1018
rect 27700 -1050 27780 -1030
rect 27810 -1028 28010 -1022
rect 27810 -1062 27822 -1028
rect 27998 -1030 28010 -1028
rect 28308 -1028 28508 -1022
rect 28308 -1030 28320 -1028
rect 27998 -1040 28320 -1030
rect 27998 -1060 28130 -1040
rect 27998 -1062 28010 -1060
rect 27810 -1068 28010 -1062
rect 28120 -1100 28130 -1060
rect 28190 -1060 28320 -1040
rect 28190 -1100 28200 -1060
rect 28308 -1062 28320 -1060
rect 28496 -1062 28508 -1028
rect 28540 -1030 28550 -970
rect 28610 -1030 28620 -970
rect 28540 -1050 28620 -1030
rect 28308 -1068 28508 -1062
rect 28120 -1110 28200 -1100
rect 27590 -1710 27660 -1130
rect 28670 -1130 28680 -890
rect 28720 -1130 28740 -890
rect 28670 -1600 28740 -1130
rect 28660 -1640 28740 -1630
rect 28660 -1700 28670 -1640
rect 28730 -1700 28740 -1640
rect 28660 -1710 28740 -1700
rect 28770 -1710 28800 130
rect 28860 -1710 28890 130
rect 28920 -1710 28950 130
rect 29040 -1710 29070 130
rect 29160 -1710 29190 130
rect 29280 -1710 29310 130
rect 29400 -1710 29430 130
rect 29520 -1710 29550 130
rect 29640 -1710 29670 130
rect 31800 -1710 31830 150
rect 31920 -1710 31950 150
rect 32040 -1710 32070 150
rect 32160 -1710 32190 150
rect 32280 -1710 32310 150
rect 32400 -1710 32430 150
rect 32520 -1710 32550 150
rect 32580 140 32660 150
rect 32580 80 32590 140
rect 32650 80 32660 140
rect 32580 70 32660 80
rect 32580 -110 32650 70
rect 33660 0 33730 130
rect 32580 -120 33730 -110
rect 32580 -180 32590 -120
rect 32650 -170 33730 -120
rect 32650 -180 32660 -170
rect 32580 -190 32660 -180
rect 32580 -570 32650 -190
rect 32580 -810 32600 -570
rect 32640 -810 32650 -570
rect 33660 -570 33730 -170
rect 33110 -590 33190 -580
rect 32800 -630 33000 -624
rect 33110 -630 33120 -590
rect 32690 -660 32770 -640
rect 32690 -720 32700 -660
rect 32760 -674 32770 -660
rect 32800 -664 32812 -630
rect 32988 -650 33120 -630
rect 33180 -630 33190 -590
rect 33298 -630 33498 -624
rect 33180 -650 33310 -630
rect 32988 -660 33310 -650
rect 32988 -664 33000 -660
rect 32800 -670 33000 -664
rect 33298 -664 33310 -660
rect 33486 -664 33498 -630
rect 33298 -670 33498 -664
rect 33530 -660 33610 -640
rect 32762 -708 32770 -674
rect 32760 -720 32770 -708
rect 32690 -740 32770 -720
rect 32800 -718 33000 -712
rect 32800 -752 32812 -718
rect 32988 -720 33000 -718
rect 33298 -718 33498 -712
rect 33298 -720 33310 -718
rect 32988 -750 33310 -720
rect 32988 -752 33000 -750
rect 32800 -758 33000 -752
rect 32580 -870 32650 -810
rect 32580 -1130 32600 -870
rect 32640 -1130 32650 -870
rect 33110 -760 33190 -750
rect 33298 -752 33310 -750
rect 33486 -752 33498 -718
rect 33530 -720 33540 -660
rect 33600 -720 33610 -660
rect 33530 -740 33610 -720
rect 33298 -758 33498 -752
rect 33110 -820 33120 -760
rect 33180 -820 33190 -760
rect 33110 -870 33190 -820
rect 33110 -930 33120 -870
rect 33180 -930 33190 -870
rect 32800 -940 33000 -934
rect 33110 -940 33190 -930
rect 33660 -810 33670 -570
rect 33710 -810 33730 -570
rect 33660 -890 33730 -810
rect 33298 -940 33498 -934
rect 32690 -970 32770 -950
rect 32690 -1030 32700 -970
rect 32760 -984 32770 -970
rect 32800 -974 32812 -940
rect 32988 -970 33310 -940
rect 32988 -974 33000 -970
rect 32800 -980 33000 -974
rect 33298 -974 33310 -970
rect 33486 -974 33498 -940
rect 33298 -980 33498 -974
rect 33530 -970 33610 -950
rect 32762 -1018 32770 -984
rect 32760 -1030 32770 -1018
rect 32690 -1050 32770 -1030
rect 32800 -1028 33000 -1022
rect 32800 -1062 32812 -1028
rect 32988 -1030 33000 -1028
rect 33298 -1028 33498 -1022
rect 33298 -1030 33310 -1028
rect 32988 -1040 33310 -1030
rect 32988 -1060 33120 -1040
rect 32988 -1062 33000 -1060
rect 32800 -1068 33000 -1062
rect 33110 -1100 33120 -1060
rect 33180 -1060 33310 -1040
rect 33180 -1100 33190 -1060
rect 33298 -1062 33310 -1060
rect 33486 -1062 33498 -1028
rect 33530 -1030 33540 -970
rect 33600 -1030 33610 -970
rect 33530 -1050 33610 -1030
rect 33298 -1068 33498 -1062
rect 33110 -1110 33190 -1100
rect 32580 -1710 32650 -1130
rect 33660 -1130 33670 -890
rect 33710 -1130 33730 -890
rect 33660 -1600 33730 -1130
rect 33650 -1640 33730 -1630
rect 33650 -1700 33660 -1640
rect 33720 -1700 33730 -1640
rect 33650 -1710 33730 -1700
rect 33760 -1710 33790 130
rect 33850 -1710 33880 130
rect 33910 -1710 33940 130
rect 34030 -1710 34060 130
rect 34150 -1710 34180 130
rect 34270 -1710 34300 130
rect 34390 -1710 34420 130
rect 34510 -1710 34540 130
rect 34630 -1710 34660 130
rect 36790 -1710 36820 150
rect 36910 -1710 36940 150
rect 37030 -1710 37060 150
rect 37150 -1710 37180 150
rect 37270 -1710 37300 150
rect 37390 -1710 37420 150
rect 37510 -1710 37540 150
rect 37570 140 37650 150
rect 37570 80 37580 140
rect 37640 80 37650 140
rect 37570 70 37650 80
rect 37570 -110 37640 70
rect 38650 0 38720 130
rect 37570 -120 38720 -110
rect 37570 -180 37580 -120
rect 37640 -170 38720 -120
rect 37640 -180 37650 -170
rect 37570 -190 37650 -180
rect 37570 -570 37640 -190
rect 37570 -810 37590 -570
rect 37630 -810 37640 -570
rect 38650 -570 38720 -170
rect 38100 -590 38180 -580
rect 37790 -630 37990 -624
rect 38100 -630 38110 -590
rect 37680 -660 37760 -640
rect 37680 -720 37690 -660
rect 37750 -674 37760 -660
rect 37790 -664 37802 -630
rect 37978 -650 38110 -630
rect 38170 -630 38180 -590
rect 38288 -630 38488 -624
rect 38170 -650 38300 -630
rect 37978 -660 38300 -650
rect 37978 -664 37990 -660
rect 37790 -670 37990 -664
rect 38288 -664 38300 -660
rect 38476 -664 38488 -630
rect 38288 -670 38488 -664
rect 38520 -660 38600 -640
rect 37752 -708 37760 -674
rect 37750 -720 37760 -708
rect 37680 -740 37760 -720
rect 37790 -718 37990 -712
rect 37790 -752 37802 -718
rect 37978 -720 37990 -718
rect 38288 -718 38488 -712
rect 38288 -720 38300 -718
rect 37978 -750 38300 -720
rect 37978 -752 37990 -750
rect 37790 -758 37990 -752
rect 37570 -870 37640 -810
rect 37570 -1130 37590 -870
rect 37630 -1130 37640 -870
rect 38100 -760 38180 -750
rect 38288 -752 38300 -750
rect 38476 -752 38488 -718
rect 38520 -720 38530 -660
rect 38590 -720 38600 -660
rect 38520 -740 38600 -720
rect 38288 -758 38488 -752
rect 38100 -820 38110 -760
rect 38170 -820 38180 -760
rect 38100 -870 38180 -820
rect 38100 -930 38110 -870
rect 38170 -930 38180 -870
rect 37790 -940 37990 -934
rect 38100 -940 38180 -930
rect 38650 -810 38660 -570
rect 38700 -810 38720 -570
rect 38650 -890 38720 -810
rect 38288 -940 38488 -934
rect 37680 -970 37760 -950
rect 37680 -1030 37690 -970
rect 37750 -984 37760 -970
rect 37790 -974 37802 -940
rect 37978 -970 38300 -940
rect 37978 -974 37990 -970
rect 37790 -980 37990 -974
rect 38288 -974 38300 -970
rect 38476 -974 38488 -940
rect 38288 -980 38488 -974
rect 38520 -970 38600 -950
rect 37752 -1018 37760 -984
rect 37750 -1030 37760 -1018
rect 37680 -1050 37760 -1030
rect 37790 -1028 37990 -1022
rect 37790 -1062 37802 -1028
rect 37978 -1030 37990 -1028
rect 38288 -1028 38488 -1022
rect 38288 -1030 38300 -1028
rect 37978 -1040 38300 -1030
rect 37978 -1060 38110 -1040
rect 37978 -1062 37990 -1060
rect 37790 -1068 37990 -1062
rect 38100 -1100 38110 -1060
rect 38170 -1060 38300 -1040
rect 38170 -1100 38180 -1060
rect 38288 -1062 38300 -1060
rect 38476 -1062 38488 -1028
rect 38520 -1030 38530 -970
rect 38590 -1030 38600 -970
rect 38520 -1050 38600 -1030
rect 38288 -1068 38488 -1062
rect 38100 -1110 38180 -1100
rect 37570 -1710 37640 -1130
rect 38650 -1130 38660 -890
rect 38700 -1130 38720 -890
rect 38650 -1600 38720 -1130
rect 38640 -1640 38720 -1630
rect 38640 -1700 38650 -1640
rect 38710 -1700 38720 -1640
rect 38640 -1710 38720 -1700
rect 38750 -1710 38780 130
rect 38840 -1710 38870 130
rect 38900 -1710 38930 130
rect 39020 -1710 39050 130
rect 39140 -1710 39170 130
rect 39260 -1710 39290 130
rect 39380 -1710 39410 130
rect 39500 -1710 39530 130
rect 39620 -1710 39650 130
rect 41780 -1710 41810 150
rect 41900 -1710 41930 150
rect 42020 -1710 42050 150
rect 42140 -1710 42170 150
rect 42260 -1710 42290 150
rect 42380 -1710 42410 150
rect 42500 -1710 42530 150
rect 42560 140 42640 150
rect 42560 80 42570 140
rect 42630 80 42640 140
rect 42560 70 42640 80
rect 42560 -110 42630 70
rect 43640 0 43710 130
rect 42560 -120 43710 -110
rect 42560 -180 42570 -120
rect 42630 -170 43710 -120
rect 42630 -180 42640 -170
rect 42560 -190 42640 -180
rect 42560 -570 42630 -190
rect 42560 -810 42580 -570
rect 42620 -810 42630 -570
rect 43640 -570 43710 -170
rect 43090 -590 43170 -580
rect 42780 -630 42980 -624
rect 43090 -630 43100 -590
rect 42670 -660 42750 -640
rect 42670 -720 42680 -660
rect 42740 -674 42750 -660
rect 42780 -664 42792 -630
rect 42968 -650 43100 -630
rect 43160 -630 43170 -590
rect 43278 -630 43478 -624
rect 43160 -650 43290 -630
rect 42968 -660 43290 -650
rect 42968 -664 42980 -660
rect 42780 -670 42980 -664
rect 43278 -664 43290 -660
rect 43466 -664 43478 -630
rect 43278 -670 43478 -664
rect 43510 -660 43590 -640
rect 42742 -708 42750 -674
rect 42740 -720 42750 -708
rect 42670 -740 42750 -720
rect 42780 -718 42980 -712
rect 42780 -752 42792 -718
rect 42968 -720 42980 -718
rect 43278 -718 43478 -712
rect 43278 -720 43290 -718
rect 42968 -750 43290 -720
rect 42968 -752 42980 -750
rect 42780 -758 42980 -752
rect 42560 -870 42630 -810
rect 42560 -1130 42580 -870
rect 42620 -1130 42630 -870
rect 43090 -760 43170 -750
rect 43278 -752 43290 -750
rect 43466 -752 43478 -718
rect 43510 -720 43520 -660
rect 43580 -720 43590 -660
rect 43510 -740 43590 -720
rect 43278 -758 43478 -752
rect 43090 -820 43100 -760
rect 43160 -820 43170 -760
rect 43090 -870 43170 -820
rect 43090 -930 43100 -870
rect 43160 -930 43170 -870
rect 42780 -940 42980 -934
rect 43090 -940 43170 -930
rect 43640 -810 43650 -570
rect 43690 -810 43710 -570
rect 43640 -890 43710 -810
rect 43278 -940 43478 -934
rect 42670 -970 42750 -950
rect 42670 -1030 42680 -970
rect 42740 -984 42750 -970
rect 42780 -974 42792 -940
rect 42968 -970 43290 -940
rect 42968 -974 42980 -970
rect 42780 -980 42980 -974
rect 43278 -974 43290 -970
rect 43466 -974 43478 -940
rect 43278 -980 43478 -974
rect 43510 -970 43590 -950
rect 42742 -1018 42750 -984
rect 42740 -1030 42750 -1018
rect 42670 -1050 42750 -1030
rect 42780 -1028 42980 -1022
rect 42780 -1062 42792 -1028
rect 42968 -1030 42980 -1028
rect 43278 -1028 43478 -1022
rect 43278 -1030 43290 -1028
rect 42968 -1040 43290 -1030
rect 42968 -1060 43100 -1040
rect 42968 -1062 42980 -1060
rect 42780 -1068 42980 -1062
rect 43090 -1100 43100 -1060
rect 43160 -1060 43290 -1040
rect 43160 -1100 43170 -1060
rect 43278 -1062 43290 -1060
rect 43466 -1062 43478 -1028
rect 43510 -1030 43520 -970
rect 43580 -1030 43590 -970
rect 43510 -1050 43590 -1030
rect 43278 -1068 43478 -1062
rect 43090 -1110 43170 -1100
rect 42560 -1710 42630 -1130
rect 43640 -1130 43650 -890
rect 43690 -1130 43710 -890
rect 43640 -1600 43710 -1130
rect 43630 -1640 43710 -1630
rect 43630 -1700 43640 -1640
rect 43700 -1700 43710 -1640
rect 43630 -1710 43710 -1700
rect 43740 -1710 43770 130
rect 43830 -1710 43860 130
rect 43890 -1710 43920 130
rect 44010 -1710 44040 130
rect 44130 -1710 44160 130
rect 44250 -1710 44280 130
rect 44370 -1710 44400 130
rect 44490 -1710 44520 130
rect 44610 -1710 44640 130
rect 46770 -1710 46800 150
rect 46890 -1710 46920 150
rect 47010 -1710 47040 150
rect 47130 -1710 47160 150
rect 47250 -1710 47280 150
rect 47370 -1710 47400 150
rect 47490 -1710 47520 150
rect 47550 140 47630 150
rect 47550 80 47560 140
rect 47620 80 47630 140
rect 47550 70 47630 80
rect 47550 -110 47620 70
rect 48630 0 48700 130
rect 47550 -120 48700 -110
rect 47550 -180 47560 -120
rect 47620 -170 48700 -120
rect 47620 -180 47630 -170
rect 47550 -190 47630 -180
rect 47550 -570 47620 -190
rect 47550 -810 47570 -570
rect 47610 -810 47620 -570
rect 48630 -570 48700 -170
rect 48080 -590 48160 -580
rect 47770 -630 47970 -624
rect 48080 -630 48090 -590
rect 47660 -660 47740 -640
rect 47660 -720 47670 -660
rect 47730 -674 47740 -660
rect 47770 -664 47782 -630
rect 47958 -650 48090 -630
rect 48150 -630 48160 -590
rect 48268 -630 48468 -624
rect 48150 -650 48280 -630
rect 47958 -660 48280 -650
rect 47958 -664 47970 -660
rect 47770 -670 47970 -664
rect 48268 -664 48280 -660
rect 48456 -664 48468 -630
rect 48268 -670 48468 -664
rect 48500 -660 48580 -640
rect 47732 -708 47740 -674
rect 47730 -720 47740 -708
rect 47660 -740 47740 -720
rect 47770 -718 47970 -712
rect 47770 -752 47782 -718
rect 47958 -720 47970 -718
rect 48268 -718 48468 -712
rect 48268 -720 48280 -718
rect 47958 -750 48280 -720
rect 47958 -752 47970 -750
rect 47770 -758 47970 -752
rect 47550 -870 47620 -810
rect 47550 -1130 47570 -870
rect 47610 -1130 47620 -870
rect 48080 -760 48160 -750
rect 48268 -752 48280 -750
rect 48456 -752 48468 -718
rect 48500 -720 48510 -660
rect 48570 -720 48580 -660
rect 48500 -740 48580 -720
rect 48268 -758 48468 -752
rect 48080 -820 48090 -760
rect 48150 -820 48160 -760
rect 48080 -870 48160 -820
rect 48080 -930 48090 -870
rect 48150 -930 48160 -870
rect 47770 -940 47970 -934
rect 48080 -940 48160 -930
rect 48630 -810 48640 -570
rect 48680 -810 48700 -570
rect 48630 -890 48700 -810
rect 48268 -940 48468 -934
rect 47660 -970 47740 -950
rect 47660 -1030 47670 -970
rect 47730 -984 47740 -970
rect 47770 -974 47782 -940
rect 47958 -970 48280 -940
rect 47958 -974 47970 -970
rect 47770 -980 47970 -974
rect 48268 -974 48280 -970
rect 48456 -974 48468 -940
rect 48268 -980 48468 -974
rect 48500 -970 48580 -950
rect 47732 -1018 47740 -984
rect 47730 -1030 47740 -1018
rect 47660 -1050 47740 -1030
rect 47770 -1028 47970 -1022
rect 47770 -1062 47782 -1028
rect 47958 -1030 47970 -1028
rect 48268 -1028 48468 -1022
rect 48268 -1030 48280 -1028
rect 47958 -1040 48280 -1030
rect 47958 -1060 48090 -1040
rect 47958 -1062 47970 -1060
rect 47770 -1068 47970 -1062
rect 48080 -1100 48090 -1060
rect 48150 -1060 48280 -1040
rect 48150 -1100 48160 -1060
rect 48268 -1062 48280 -1060
rect 48456 -1062 48468 -1028
rect 48500 -1030 48510 -970
rect 48570 -1030 48580 -970
rect 48500 -1050 48580 -1030
rect 48268 -1068 48468 -1062
rect 48080 -1110 48160 -1100
rect 47550 -1710 47620 -1130
rect 48630 -1130 48640 -890
rect 48680 -1130 48700 -890
rect 48630 -1600 48700 -1130
rect 48620 -1640 48700 -1630
rect 48620 -1700 48630 -1640
rect 48690 -1700 48700 -1640
rect 48620 -1710 48700 -1700
rect 48730 -1710 48760 130
rect 48820 -1710 48850 130
rect 48880 -1710 48910 130
rect 49000 -1710 49030 130
rect 49120 -1710 49150 130
rect 49240 -1710 49270 130
rect 49360 -1710 49390 130
rect 49480 -1710 49510 130
rect 49600 -1710 49630 130
rect 51760 -1710 51790 150
rect 51880 -1710 51910 150
rect 52000 -1710 52030 150
rect 52120 -1710 52150 150
rect 52240 -1710 52270 150
rect 52360 -1710 52390 150
rect 52480 -1710 52510 150
rect 52540 140 52620 150
rect 52540 80 52550 140
rect 52610 80 52620 140
rect 52540 70 52620 80
rect 52540 -110 52610 70
rect 53620 0 53690 130
rect 52540 -120 53690 -110
rect 52540 -180 52550 -120
rect 52610 -170 53690 -120
rect 52610 -180 52620 -170
rect 52540 -190 52620 -180
rect 52540 -570 52610 -190
rect 52540 -810 52560 -570
rect 52600 -810 52610 -570
rect 53620 -570 53690 -170
rect 53070 -590 53150 -580
rect 52760 -630 52960 -624
rect 53070 -630 53080 -590
rect 52650 -660 52730 -640
rect 52650 -720 52660 -660
rect 52720 -674 52730 -660
rect 52760 -664 52772 -630
rect 52948 -650 53080 -630
rect 53140 -630 53150 -590
rect 53258 -630 53458 -624
rect 53140 -650 53270 -630
rect 52948 -660 53270 -650
rect 52948 -664 52960 -660
rect 52760 -670 52960 -664
rect 53258 -664 53270 -660
rect 53446 -664 53458 -630
rect 53258 -670 53458 -664
rect 53490 -660 53570 -640
rect 52722 -708 52730 -674
rect 52720 -720 52730 -708
rect 52650 -740 52730 -720
rect 52760 -718 52960 -712
rect 52760 -752 52772 -718
rect 52948 -720 52960 -718
rect 53258 -718 53458 -712
rect 53258 -720 53270 -718
rect 52948 -750 53270 -720
rect 52948 -752 52960 -750
rect 52760 -758 52960 -752
rect 52540 -870 52610 -810
rect 52540 -1130 52560 -870
rect 52600 -1130 52610 -870
rect 53070 -760 53150 -750
rect 53258 -752 53270 -750
rect 53446 -752 53458 -718
rect 53490 -720 53500 -660
rect 53560 -720 53570 -660
rect 53490 -740 53570 -720
rect 53258 -758 53458 -752
rect 53070 -820 53080 -760
rect 53140 -820 53150 -760
rect 53070 -870 53150 -820
rect 53070 -930 53080 -870
rect 53140 -930 53150 -870
rect 52760 -940 52960 -934
rect 53070 -940 53150 -930
rect 53620 -810 53630 -570
rect 53670 -810 53690 -570
rect 53620 -890 53690 -810
rect 53258 -940 53458 -934
rect 52650 -970 52730 -950
rect 52650 -1030 52660 -970
rect 52720 -984 52730 -970
rect 52760 -974 52772 -940
rect 52948 -970 53270 -940
rect 52948 -974 52960 -970
rect 52760 -980 52960 -974
rect 53258 -974 53270 -970
rect 53446 -974 53458 -940
rect 53258 -980 53458 -974
rect 53490 -970 53570 -950
rect 52722 -1018 52730 -984
rect 52720 -1030 52730 -1018
rect 52650 -1050 52730 -1030
rect 52760 -1028 52960 -1022
rect 52760 -1062 52772 -1028
rect 52948 -1030 52960 -1028
rect 53258 -1028 53458 -1022
rect 53258 -1030 53270 -1028
rect 52948 -1040 53270 -1030
rect 52948 -1060 53080 -1040
rect 52948 -1062 52960 -1060
rect 52760 -1068 52960 -1062
rect 53070 -1100 53080 -1060
rect 53140 -1060 53270 -1040
rect 53140 -1100 53150 -1060
rect 53258 -1062 53270 -1060
rect 53446 -1062 53458 -1028
rect 53490 -1030 53500 -970
rect 53560 -1030 53570 -970
rect 53490 -1050 53570 -1030
rect 53258 -1068 53458 -1062
rect 53070 -1110 53150 -1100
rect 52540 -1710 52610 -1130
rect 53620 -1130 53630 -890
rect 53670 -1130 53690 -890
rect 53620 -1600 53690 -1130
rect 53610 -1640 53690 -1630
rect 53610 -1700 53620 -1640
rect 53680 -1700 53690 -1640
rect 53610 -1710 53690 -1700
rect 53720 -1710 53750 130
rect 53810 -1710 53840 130
rect 53870 -1710 53900 130
rect 53990 -1710 54020 130
rect 54110 -1710 54140 130
rect 54230 -1710 54260 130
rect 54350 -1710 54380 130
rect 54470 -1710 54500 130
rect 54590 -1710 54620 130
rect 56750 -1710 56780 150
rect 56870 -1710 56900 150
rect 56990 -1710 57020 150
rect 57110 -1710 57140 150
rect 57230 -1710 57260 150
rect 57350 -1710 57380 150
rect 57470 -1710 57500 150
rect 57530 140 57610 150
rect 57530 80 57540 140
rect 57600 80 57610 140
rect 57530 70 57610 80
rect 57530 -110 57600 70
rect 58610 0 58680 130
rect 57530 -120 58680 -110
rect 57530 -180 57540 -120
rect 57600 -170 58680 -120
rect 57600 -180 57610 -170
rect 57530 -190 57610 -180
rect 57530 -570 57600 -190
rect 57530 -810 57550 -570
rect 57590 -810 57600 -570
rect 58610 -570 58680 -170
rect 58060 -590 58140 -580
rect 57750 -630 57950 -624
rect 58060 -630 58070 -590
rect 57640 -660 57720 -640
rect 57640 -720 57650 -660
rect 57710 -674 57720 -660
rect 57750 -664 57762 -630
rect 57938 -650 58070 -630
rect 58130 -630 58140 -590
rect 58248 -630 58448 -624
rect 58130 -650 58260 -630
rect 57938 -660 58260 -650
rect 57938 -664 57950 -660
rect 57750 -670 57950 -664
rect 58248 -664 58260 -660
rect 58436 -664 58448 -630
rect 58248 -670 58448 -664
rect 58480 -660 58560 -640
rect 57712 -708 57720 -674
rect 57710 -720 57720 -708
rect 57640 -740 57720 -720
rect 57750 -718 57950 -712
rect 57750 -752 57762 -718
rect 57938 -720 57950 -718
rect 58248 -718 58448 -712
rect 58248 -720 58260 -718
rect 57938 -750 58260 -720
rect 57938 -752 57950 -750
rect 57750 -758 57950 -752
rect 57530 -870 57600 -810
rect 57530 -1130 57550 -870
rect 57590 -1130 57600 -870
rect 58060 -760 58140 -750
rect 58248 -752 58260 -750
rect 58436 -752 58448 -718
rect 58480 -720 58490 -660
rect 58550 -720 58560 -660
rect 58480 -740 58560 -720
rect 58248 -758 58448 -752
rect 58060 -820 58070 -760
rect 58130 -820 58140 -760
rect 58060 -870 58140 -820
rect 58060 -930 58070 -870
rect 58130 -930 58140 -870
rect 57750 -940 57950 -934
rect 58060 -940 58140 -930
rect 58610 -810 58620 -570
rect 58660 -810 58680 -570
rect 58610 -890 58680 -810
rect 58248 -940 58448 -934
rect 57640 -970 57720 -950
rect 57640 -1030 57650 -970
rect 57710 -984 57720 -970
rect 57750 -974 57762 -940
rect 57938 -970 58260 -940
rect 57938 -974 57950 -970
rect 57750 -980 57950 -974
rect 58248 -974 58260 -970
rect 58436 -974 58448 -940
rect 58248 -980 58448 -974
rect 58480 -970 58560 -950
rect 57712 -1018 57720 -984
rect 57710 -1030 57720 -1018
rect 57640 -1050 57720 -1030
rect 57750 -1028 57950 -1022
rect 57750 -1062 57762 -1028
rect 57938 -1030 57950 -1028
rect 58248 -1028 58448 -1022
rect 58248 -1030 58260 -1028
rect 57938 -1040 58260 -1030
rect 57938 -1060 58070 -1040
rect 57938 -1062 57950 -1060
rect 57750 -1068 57950 -1062
rect 58060 -1100 58070 -1060
rect 58130 -1060 58260 -1040
rect 58130 -1100 58140 -1060
rect 58248 -1062 58260 -1060
rect 58436 -1062 58448 -1028
rect 58480 -1030 58490 -970
rect 58550 -1030 58560 -970
rect 58480 -1050 58560 -1030
rect 58248 -1068 58448 -1062
rect 58060 -1110 58140 -1100
rect 57530 -1710 57600 -1130
rect 58610 -1130 58620 -890
rect 58660 -1130 58680 -890
rect 58610 -1600 58680 -1130
rect 58600 -1640 58680 -1630
rect 58600 -1700 58610 -1640
rect 58670 -1700 58680 -1640
rect 58600 -1710 58680 -1700
rect 58710 -1710 58740 130
rect 58800 -1710 58830 130
rect 58860 -1710 58890 130
rect 58980 -1710 59010 130
rect 59100 -1710 59130 130
rect 59220 -1710 59250 130
rect 59340 -1710 59370 130
rect 59460 -1710 59490 130
rect 59580 -1710 59610 130
rect 61740 -1710 61770 150
rect 61860 -1710 61890 150
rect 61980 -1710 62010 150
rect 62100 -1710 62130 150
rect 62220 -1710 62250 150
rect 62340 -1710 62370 150
rect 62460 -1710 62490 150
rect 62520 140 62600 150
rect 62520 80 62530 140
rect 62590 80 62600 140
rect 62520 70 62600 80
rect 62520 -110 62590 70
rect 63600 0 63670 130
rect 62520 -120 63670 -110
rect 62520 -180 62530 -120
rect 62590 -170 63670 -120
rect 62590 -180 62600 -170
rect 62520 -190 62600 -180
rect 62520 -570 62590 -190
rect 62520 -810 62540 -570
rect 62580 -810 62590 -570
rect 63600 -570 63670 -170
rect 63050 -590 63130 -580
rect 62740 -630 62940 -624
rect 63050 -630 63060 -590
rect 62630 -660 62710 -640
rect 62630 -720 62640 -660
rect 62700 -674 62710 -660
rect 62740 -664 62752 -630
rect 62928 -650 63060 -630
rect 63120 -630 63130 -590
rect 63238 -630 63438 -624
rect 63120 -650 63250 -630
rect 62928 -660 63250 -650
rect 62928 -664 62940 -660
rect 62740 -670 62940 -664
rect 63238 -664 63250 -660
rect 63426 -664 63438 -630
rect 63238 -670 63438 -664
rect 63470 -660 63550 -640
rect 62702 -708 62710 -674
rect 62700 -720 62710 -708
rect 62630 -740 62710 -720
rect 62740 -718 62940 -712
rect 62740 -752 62752 -718
rect 62928 -720 62940 -718
rect 63238 -718 63438 -712
rect 63238 -720 63250 -718
rect 62928 -750 63250 -720
rect 62928 -752 62940 -750
rect 62740 -758 62940 -752
rect 62520 -870 62590 -810
rect 62520 -1130 62540 -870
rect 62580 -1130 62590 -870
rect 63050 -760 63130 -750
rect 63238 -752 63250 -750
rect 63426 -752 63438 -718
rect 63470 -720 63480 -660
rect 63540 -720 63550 -660
rect 63470 -740 63550 -720
rect 63238 -758 63438 -752
rect 63050 -820 63060 -760
rect 63120 -820 63130 -760
rect 63050 -870 63130 -820
rect 63050 -930 63060 -870
rect 63120 -930 63130 -870
rect 62740 -940 62940 -934
rect 63050 -940 63130 -930
rect 63600 -810 63610 -570
rect 63650 -810 63670 -570
rect 63600 -890 63670 -810
rect 63238 -940 63438 -934
rect 62630 -970 62710 -950
rect 62630 -1030 62640 -970
rect 62700 -984 62710 -970
rect 62740 -974 62752 -940
rect 62928 -970 63250 -940
rect 62928 -974 62940 -970
rect 62740 -980 62940 -974
rect 63238 -974 63250 -970
rect 63426 -974 63438 -940
rect 63238 -980 63438 -974
rect 63470 -970 63550 -950
rect 62702 -1018 62710 -984
rect 62700 -1030 62710 -1018
rect 62630 -1050 62710 -1030
rect 62740 -1028 62940 -1022
rect 62740 -1062 62752 -1028
rect 62928 -1030 62940 -1028
rect 63238 -1028 63438 -1022
rect 63238 -1030 63250 -1028
rect 62928 -1040 63250 -1030
rect 62928 -1060 63060 -1040
rect 62928 -1062 62940 -1060
rect 62740 -1068 62940 -1062
rect 63050 -1100 63060 -1060
rect 63120 -1060 63250 -1040
rect 63120 -1100 63130 -1060
rect 63238 -1062 63250 -1060
rect 63426 -1062 63438 -1028
rect 63470 -1030 63480 -970
rect 63540 -1030 63550 -970
rect 63470 -1050 63550 -1030
rect 63238 -1068 63438 -1062
rect 63050 -1110 63130 -1100
rect 62520 -1710 62590 -1130
rect 63600 -1130 63610 -890
rect 63650 -1130 63670 -890
rect 63600 -1600 63670 -1130
rect 63590 -1640 63670 -1630
rect 63590 -1700 63600 -1640
rect 63660 -1700 63670 -1640
rect 63590 -1710 63670 -1700
rect 63700 -1710 63730 130
rect 63790 -1710 63820 130
rect 63850 -1710 63880 130
rect 63970 -1710 64000 130
rect 64090 -1710 64120 130
rect 64210 -1710 64240 130
rect 64330 -1710 64360 130
rect 64450 -1710 64480 130
rect 64570 -1710 64600 130
rect 66730 -1710 66760 150
rect 66850 -1710 66880 150
rect 66970 -1710 67000 150
rect 67090 -1710 67120 150
rect 67210 -1710 67240 150
rect 67330 -1710 67360 150
rect 67450 -1710 67480 150
rect 67510 140 67590 150
rect 67510 80 67520 140
rect 67580 80 67590 140
rect 67510 70 67590 80
rect 67510 -110 67580 70
rect 68590 0 68660 130
rect 67510 -120 68660 -110
rect 67510 -180 67520 -120
rect 67580 -170 68660 -120
rect 67580 -180 67590 -170
rect 67510 -190 67590 -180
rect 67510 -570 67580 -190
rect 67510 -810 67530 -570
rect 67570 -810 67580 -570
rect 68590 -570 68660 -170
rect 68040 -590 68120 -580
rect 67730 -630 67930 -624
rect 68040 -630 68050 -590
rect 67620 -660 67700 -640
rect 67620 -720 67630 -660
rect 67690 -674 67700 -660
rect 67730 -664 67742 -630
rect 67918 -650 68050 -630
rect 68110 -630 68120 -590
rect 68228 -630 68428 -624
rect 68110 -650 68240 -630
rect 67918 -660 68240 -650
rect 67918 -664 67930 -660
rect 67730 -670 67930 -664
rect 68228 -664 68240 -660
rect 68416 -664 68428 -630
rect 68228 -670 68428 -664
rect 68460 -660 68540 -640
rect 67692 -708 67700 -674
rect 67690 -720 67700 -708
rect 67620 -740 67700 -720
rect 67730 -718 67930 -712
rect 67730 -752 67742 -718
rect 67918 -720 67930 -718
rect 68228 -718 68428 -712
rect 68228 -720 68240 -718
rect 67918 -750 68240 -720
rect 67918 -752 67930 -750
rect 67730 -758 67930 -752
rect 67510 -870 67580 -810
rect 67510 -1130 67530 -870
rect 67570 -1130 67580 -870
rect 68040 -760 68120 -750
rect 68228 -752 68240 -750
rect 68416 -752 68428 -718
rect 68460 -720 68470 -660
rect 68530 -720 68540 -660
rect 68460 -740 68540 -720
rect 68228 -758 68428 -752
rect 68040 -820 68050 -760
rect 68110 -820 68120 -760
rect 68040 -870 68120 -820
rect 68040 -930 68050 -870
rect 68110 -930 68120 -870
rect 67730 -940 67930 -934
rect 68040 -940 68120 -930
rect 68590 -810 68600 -570
rect 68640 -810 68660 -570
rect 68590 -890 68660 -810
rect 68228 -940 68428 -934
rect 67620 -970 67700 -950
rect 67620 -1030 67630 -970
rect 67690 -984 67700 -970
rect 67730 -974 67742 -940
rect 67918 -970 68240 -940
rect 67918 -974 67930 -970
rect 67730 -980 67930 -974
rect 68228 -974 68240 -970
rect 68416 -974 68428 -940
rect 68228 -980 68428 -974
rect 68460 -970 68540 -950
rect 67692 -1018 67700 -984
rect 67690 -1030 67700 -1018
rect 67620 -1050 67700 -1030
rect 67730 -1028 67930 -1022
rect 67730 -1062 67742 -1028
rect 67918 -1030 67930 -1028
rect 68228 -1028 68428 -1022
rect 68228 -1030 68240 -1028
rect 67918 -1040 68240 -1030
rect 67918 -1060 68050 -1040
rect 67918 -1062 67930 -1060
rect 67730 -1068 67930 -1062
rect 68040 -1100 68050 -1060
rect 68110 -1060 68240 -1040
rect 68110 -1100 68120 -1060
rect 68228 -1062 68240 -1060
rect 68416 -1062 68428 -1028
rect 68460 -1030 68470 -970
rect 68530 -1030 68540 -970
rect 68460 -1050 68540 -1030
rect 68228 -1068 68428 -1062
rect 68040 -1110 68120 -1100
rect 67510 -1710 67580 -1130
rect 68590 -1130 68600 -890
rect 68640 -1130 68660 -890
rect 68590 -1600 68660 -1130
rect 68580 -1640 68660 -1630
rect 68580 -1700 68590 -1640
rect 68650 -1700 68660 -1640
rect 68580 -1710 68660 -1700
rect 68690 -1710 68720 130
rect 68780 -1710 68810 130
rect 68840 -1710 68870 130
rect 68960 -1710 68990 130
rect 69080 -1710 69110 130
rect 69200 -1710 69230 130
rect 69320 -1710 69350 130
rect 69440 -1710 69470 130
rect 69560 -1710 69590 130
rect 71720 -1710 71750 150
rect 71840 -1710 71870 150
rect 71960 -1710 71990 150
rect 72080 -1710 72110 150
rect 72200 -1710 72230 150
rect 72320 -1710 72350 150
rect 72440 -1710 72470 150
rect 72500 140 72580 150
rect 72500 80 72510 140
rect 72570 80 72580 140
rect 72500 70 72580 80
rect 72500 -110 72570 70
rect 73580 0 73650 130
rect 72500 -120 73650 -110
rect 72500 -180 72510 -120
rect 72570 -170 73650 -120
rect 72570 -180 72580 -170
rect 72500 -190 72580 -180
rect 72500 -570 72570 -190
rect 72500 -810 72520 -570
rect 72560 -810 72570 -570
rect 73580 -570 73650 -170
rect 73030 -590 73110 -580
rect 72720 -630 72920 -624
rect 73030 -630 73040 -590
rect 72610 -660 72690 -640
rect 72610 -720 72620 -660
rect 72680 -674 72690 -660
rect 72720 -664 72732 -630
rect 72908 -650 73040 -630
rect 73100 -630 73110 -590
rect 73218 -630 73418 -624
rect 73100 -650 73230 -630
rect 72908 -660 73230 -650
rect 72908 -664 72920 -660
rect 72720 -670 72920 -664
rect 73218 -664 73230 -660
rect 73406 -664 73418 -630
rect 73218 -670 73418 -664
rect 73450 -660 73530 -640
rect 72682 -708 72690 -674
rect 72680 -720 72690 -708
rect 72610 -740 72690 -720
rect 72720 -718 72920 -712
rect 72720 -752 72732 -718
rect 72908 -720 72920 -718
rect 73218 -718 73418 -712
rect 73218 -720 73230 -718
rect 72908 -750 73230 -720
rect 72908 -752 72920 -750
rect 72720 -758 72920 -752
rect 72500 -870 72570 -810
rect 72500 -1130 72520 -870
rect 72560 -1130 72570 -870
rect 73030 -760 73110 -750
rect 73218 -752 73230 -750
rect 73406 -752 73418 -718
rect 73450 -720 73460 -660
rect 73520 -720 73530 -660
rect 73450 -740 73530 -720
rect 73218 -758 73418 -752
rect 73030 -820 73040 -760
rect 73100 -820 73110 -760
rect 73030 -870 73110 -820
rect 73030 -930 73040 -870
rect 73100 -930 73110 -870
rect 72720 -940 72920 -934
rect 73030 -940 73110 -930
rect 73580 -810 73590 -570
rect 73630 -810 73650 -570
rect 73580 -890 73650 -810
rect 73218 -940 73418 -934
rect 72610 -970 72690 -950
rect 72610 -1030 72620 -970
rect 72680 -984 72690 -970
rect 72720 -974 72732 -940
rect 72908 -970 73230 -940
rect 72908 -974 72920 -970
rect 72720 -980 72920 -974
rect 73218 -974 73230 -970
rect 73406 -974 73418 -940
rect 73218 -980 73418 -974
rect 73450 -970 73530 -950
rect 72682 -1018 72690 -984
rect 72680 -1030 72690 -1018
rect 72610 -1050 72690 -1030
rect 72720 -1028 72920 -1022
rect 72720 -1062 72732 -1028
rect 72908 -1030 72920 -1028
rect 73218 -1028 73418 -1022
rect 73218 -1030 73230 -1028
rect 72908 -1040 73230 -1030
rect 72908 -1060 73040 -1040
rect 72908 -1062 72920 -1060
rect 72720 -1068 72920 -1062
rect 73030 -1100 73040 -1060
rect 73100 -1060 73230 -1040
rect 73100 -1100 73110 -1060
rect 73218 -1062 73230 -1060
rect 73406 -1062 73418 -1028
rect 73450 -1030 73460 -970
rect 73520 -1030 73530 -970
rect 73450 -1050 73530 -1030
rect 73218 -1068 73418 -1062
rect 73030 -1110 73110 -1100
rect 72500 -1710 72570 -1130
rect 73580 -1130 73590 -890
rect 73630 -1130 73650 -890
rect 73580 -1600 73650 -1130
rect 73570 -1640 73650 -1630
rect 73570 -1700 73580 -1640
rect 73640 -1700 73650 -1640
rect 73570 -1710 73650 -1700
rect 73680 -1710 73710 130
rect 73770 -1710 73800 130
rect 73830 -1710 73860 130
rect 73950 -1710 73980 130
rect 74070 -1710 74100 130
rect 74190 -1710 74220 130
rect 74310 -1710 74340 130
rect 74430 -1710 74460 130
rect 74550 -1710 74580 130
rect 76710 -1710 76740 150
rect 76830 -1710 76860 150
rect 76950 -1710 76980 150
rect 77070 -1710 77100 150
rect 77190 -1710 77220 150
rect 77310 -1710 77340 150
rect 77430 -1710 77460 150
rect 77490 140 77570 150
rect 77490 80 77500 140
rect 77560 80 77570 140
rect 77490 70 77570 80
rect 77490 -110 77560 70
rect 77490 -120 78640 -110
rect 77490 -180 77500 -120
rect 77560 -170 78640 -120
rect 77560 -180 77570 -170
rect 77490 -190 77570 -180
rect 77490 -570 77560 -190
rect 77490 -810 77510 -570
rect 77550 -810 77560 -570
rect 78570 -570 78640 -170
rect 78020 -590 78100 -580
rect 77710 -630 77910 -624
rect 78020 -630 78030 -590
rect 77600 -660 77680 -640
rect 77600 -720 77610 -660
rect 77670 -674 77680 -660
rect 77710 -664 77722 -630
rect 77898 -650 78030 -630
rect 78090 -630 78100 -590
rect 78208 -630 78408 -624
rect 78090 -650 78220 -630
rect 77898 -660 78220 -650
rect 77898 -664 77910 -660
rect 77710 -670 77910 -664
rect 78208 -664 78220 -660
rect 78396 -664 78408 -630
rect 78208 -670 78408 -664
rect 78440 -660 78520 -640
rect 77672 -708 77680 -674
rect 77670 -720 77680 -708
rect 77600 -740 77680 -720
rect 77710 -718 77910 -712
rect 77710 -752 77722 -718
rect 77898 -720 77910 -718
rect 78208 -718 78408 -712
rect 78208 -720 78220 -718
rect 77898 -750 78220 -720
rect 77898 -752 77910 -750
rect 77710 -758 77910 -752
rect 77490 -870 77560 -810
rect 77490 -1130 77510 -870
rect 77550 -1130 77560 -870
rect 78020 -760 78100 -750
rect 78208 -752 78220 -750
rect 78396 -752 78408 -718
rect 78440 -720 78450 -660
rect 78510 -720 78520 -660
rect 78440 -740 78520 -720
rect 78208 -758 78408 -752
rect 78020 -820 78030 -760
rect 78090 -820 78100 -760
rect 78020 -870 78100 -820
rect 78020 -930 78030 -870
rect 78090 -930 78100 -870
rect 77710 -940 77910 -934
rect 78020 -940 78100 -930
rect 78570 -810 78580 -570
rect 78620 -810 78640 -570
rect 78570 -890 78640 -810
rect 78208 -940 78408 -934
rect 77600 -970 77680 -950
rect 77600 -1030 77610 -970
rect 77670 -984 77680 -970
rect 77710 -974 77722 -940
rect 77898 -970 78220 -940
rect 77898 -974 77910 -970
rect 77710 -980 77910 -974
rect 78208 -974 78220 -970
rect 78396 -974 78408 -940
rect 78208 -980 78408 -974
rect 78440 -970 78520 -950
rect 77672 -1018 77680 -984
rect 77670 -1030 77680 -1018
rect 77600 -1050 77680 -1030
rect 77710 -1028 77910 -1022
rect 77710 -1062 77722 -1028
rect 77898 -1030 77910 -1028
rect 78208 -1028 78408 -1022
rect 78208 -1030 78220 -1028
rect 77898 -1040 78220 -1030
rect 77898 -1060 78030 -1040
rect 77898 -1062 77910 -1060
rect 77710 -1068 77910 -1062
rect 78020 -1100 78030 -1060
rect 78090 -1060 78220 -1040
rect 78090 -1100 78100 -1060
rect 78208 -1062 78220 -1060
rect 78396 -1062 78408 -1028
rect 78440 -1030 78450 -970
rect 78510 -1030 78520 -970
rect 78440 -1050 78520 -1030
rect 78208 -1068 78408 -1062
rect 78020 -1110 78100 -1100
rect 77490 -1710 77560 -1130
rect 78570 -1130 78580 -890
rect 78620 -1130 78640 -890
rect 78570 -1600 78640 -1130
rect 78560 -1640 78640 -1630
rect 78560 -1700 78570 -1640
rect 78630 -1700 78640 -1640
rect 78560 -1710 78640 -1700
rect 78670 -1710 78700 -260
rect 78760 -1710 78790 -260
rect 78820 -1710 78850 -260
rect 78940 -1710 78970 -260
rect 79060 -1710 79090 -260
rect 79180 -1710 79210 -260
rect 79300 -1710 79330 -260
rect 79420 -1710 79450 -260
rect 79540 -1710 79570 -260
rect 81430 -1710 81460 29070
rect 81550 -1710 81580 29070
rect 81670 -1710 81700 29070
rect 81790 -1710 81820 29070
rect 81910 -1710 81940 29070
rect 82030 -1710 82060 29070
rect 82150 -1710 82180 29070
rect 82210 28960 82280 29070
rect 83280 29060 83360 29070
rect 83280 29000 83290 29060
rect 83350 29000 83360 29060
rect 83280 28990 83360 29000
rect 82210 28950 83360 28960
rect 82210 28890 82220 28950
rect 82280 28900 83360 28950
rect 82280 28890 82290 28900
rect 82210 28880 82290 28890
rect 82210 28500 82280 28880
rect 82210 28260 82230 28500
rect 82270 28260 82280 28500
rect 83290 28500 83360 28900
rect 82740 28480 82820 28490
rect 82430 28440 82630 28446
rect 82740 28440 82750 28480
rect 82320 28410 82400 28430
rect 82320 28350 82330 28410
rect 82390 28396 82400 28410
rect 82430 28406 82442 28440
rect 82618 28420 82750 28440
rect 82810 28440 82820 28480
rect 82928 28440 83128 28446
rect 82810 28420 82940 28440
rect 82618 28410 82940 28420
rect 82618 28406 82630 28410
rect 82430 28400 82630 28406
rect 82928 28406 82940 28410
rect 83116 28406 83128 28440
rect 82928 28400 83128 28406
rect 83160 28410 83240 28430
rect 82392 28362 82400 28396
rect 82390 28350 82400 28362
rect 82320 28330 82400 28350
rect 82430 28352 82630 28358
rect 82430 28318 82442 28352
rect 82618 28350 82630 28352
rect 82928 28352 83128 28358
rect 82928 28350 82940 28352
rect 82618 28320 82940 28350
rect 82618 28318 82630 28320
rect 82430 28312 82630 28318
rect 82210 28200 82280 28260
rect 82210 27940 82230 28200
rect 82270 27940 82280 28200
rect 82740 28310 82820 28320
rect 82928 28318 82940 28320
rect 83116 28318 83128 28352
rect 83160 28350 83170 28410
rect 83230 28350 83240 28410
rect 83160 28330 83240 28350
rect 82928 28312 83128 28318
rect 82740 28250 82750 28310
rect 82810 28250 82820 28310
rect 82740 28200 82820 28250
rect 82740 28140 82750 28200
rect 82810 28140 82820 28200
rect 82430 28130 82630 28136
rect 82740 28130 82820 28140
rect 83290 28260 83300 28500
rect 83340 28260 83360 28500
rect 83290 28180 83360 28260
rect 82928 28130 83128 28136
rect 82320 28100 82400 28120
rect 82320 28040 82330 28100
rect 82390 28086 82400 28100
rect 82430 28096 82442 28130
rect 82618 28100 82940 28130
rect 82618 28096 82630 28100
rect 82430 28090 82630 28096
rect 82928 28096 82940 28100
rect 83116 28096 83128 28130
rect 82928 28090 83128 28096
rect 83160 28100 83240 28120
rect 82392 28052 82400 28086
rect 82390 28040 82400 28052
rect 82320 28020 82400 28040
rect 82430 28042 82630 28048
rect 82430 28008 82442 28042
rect 82618 28040 82630 28042
rect 82928 28042 83128 28048
rect 82928 28040 82940 28042
rect 82618 28030 82940 28040
rect 82618 28010 82750 28030
rect 82618 28008 82630 28010
rect 82430 28002 82630 28008
rect 82740 27970 82750 28010
rect 82810 28010 82940 28030
rect 82810 27970 82820 28010
rect 82928 28008 82940 28010
rect 83116 28008 83128 28042
rect 83160 28040 83170 28100
rect 83230 28040 83240 28100
rect 83160 28020 83240 28040
rect 82928 28002 83128 28008
rect 82740 27960 82820 27970
rect 82210 27250 82280 27940
rect 83290 27940 83300 28180
rect 83340 27940 83360 28180
rect 83290 27530 83360 27940
rect 83270 27490 83360 27500
rect 83270 27430 83280 27490
rect 83350 27430 83360 27490
rect 83270 27420 83360 27430
rect 83290 27360 83360 27420
rect 83280 27350 83360 27360
rect 83280 27290 83290 27350
rect 83350 27290 83360 27350
rect 83280 27280 83360 27290
rect 82210 27240 83360 27250
rect 82210 27180 82220 27240
rect 82280 27190 83360 27240
rect 82280 27180 82290 27190
rect 82210 27170 82290 27180
rect 82210 26790 82280 27170
rect 82210 26550 82230 26790
rect 82270 26550 82280 26790
rect 83290 26790 83360 27190
rect 82740 26770 82820 26780
rect 82430 26730 82630 26736
rect 82740 26730 82750 26770
rect 82320 26700 82400 26720
rect 82320 26640 82330 26700
rect 82390 26686 82400 26700
rect 82430 26696 82442 26730
rect 82618 26710 82750 26730
rect 82810 26730 82820 26770
rect 82928 26730 83128 26736
rect 82810 26710 82940 26730
rect 82618 26700 82940 26710
rect 82618 26696 82630 26700
rect 82430 26690 82630 26696
rect 82928 26696 82940 26700
rect 83116 26696 83128 26730
rect 82928 26690 83128 26696
rect 83160 26700 83240 26720
rect 82392 26652 82400 26686
rect 82390 26640 82400 26652
rect 82320 26620 82400 26640
rect 82430 26642 82630 26648
rect 82430 26608 82442 26642
rect 82618 26640 82630 26642
rect 82928 26642 83128 26648
rect 82928 26640 82940 26642
rect 82618 26610 82940 26640
rect 82618 26608 82630 26610
rect 82430 26602 82630 26608
rect 82210 26490 82280 26550
rect 82210 26230 82230 26490
rect 82270 26230 82280 26490
rect 82740 26600 82820 26610
rect 82928 26608 82940 26610
rect 83116 26608 83128 26642
rect 83160 26640 83170 26700
rect 83230 26640 83240 26700
rect 83160 26620 83240 26640
rect 82928 26602 83128 26608
rect 82740 26540 82750 26600
rect 82810 26540 82820 26600
rect 82740 26490 82820 26540
rect 82740 26430 82750 26490
rect 82810 26430 82820 26490
rect 82430 26420 82630 26426
rect 82740 26420 82820 26430
rect 83290 26550 83300 26790
rect 83340 26550 83360 26790
rect 83290 26470 83360 26550
rect 82928 26420 83128 26426
rect 82320 26390 82400 26410
rect 82320 26330 82330 26390
rect 82390 26376 82400 26390
rect 82430 26386 82442 26420
rect 82618 26390 82940 26420
rect 82618 26386 82630 26390
rect 82430 26380 82630 26386
rect 82928 26386 82940 26390
rect 83116 26386 83128 26420
rect 82928 26380 83128 26386
rect 83160 26390 83240 26410
rect 82392 26342 82400 26376
rect 82390 26330 82400 26342
rect 82320 26310 82400 26330
rect 82430 26332 82630 26338
rect 82430 26298 82442 26332
rect 82618 26330 82630 26332
rect 82928 26332 83128 26338
rect 82928 26330 82940 26332
rect 82618 26320 82940 26330
rect 82618 26300 82750 26320
rect 82618 26298 82630 26300
rect 82430 26292 82630 26298
rect 82740 26260 82750 26300
rect 82810 26300 82940 26320
rect 82810 26260 82820 26300
rect 82928 26298 82940 26300
rect 83116 26298 83128 26332
rect 83160 26330 83170 26390
rect 83230 26330 83240 26390
rect 83160 26310 83240 26330
rect 82928 26292 83128 26298
rect 82740 26250 82820 26260
rect 82210 25540 82280 26230
rect 83290 26230 83300 26470
rect 83340 26230 83360 26470
rect 83290 25820 83360 26230
rect 83270 25780 83360 25790
rect 83270 25720 83280 25780
rect 83350 25720 83360 25780
rect 83270 25710 83360 25720
rect 83290 25650 83360 25710
rect 83280 25640 83360 25650
rect 83280 25580 83290 25640
rect 83350 25580 83360 25640
rect 83280 25570 83360 25580
rect 82210 25530 83360 25540
rect 82210 25470 82220 25530
rect 82280 25480 83360 25530
rect 82280 25470 82290 25480
rect 82210 25460 82290 25470
rect 82210 25080 82280 25460
rect 82210 24840 82230 25080
rect 82270 24840 82280 25080
rect 83290 25080 83360 25480
rect 82740 25060 82820 25070
rect 82430 25020 82630 25026
rect 82740 25020 82750 25060
rect 82320 24990 82400 25010
rect 82320 24930 82330 24990
rect 82390 24976 82400 24990
rect 82430 24986 82442 25020
rect 82618 25000 82750 25020
rect 82810 25020 82820 25060
rect 82928 25020 83128 25026
rect 82810 25000 82940 25020
rect 82618 24990 82940 25000
rect 82618 24986 82630 24990
rect 82430 24980 82630 24986
rect 82928 24986 82940 24990
rect 83116 24986 83128 25020
rect 82928 24980 83128 24986
rect 83160 24990 83240 25010
rect 82392 24942 82400 24976
rect 82390 24930 82400 24942
rect 82320 24910 82400 24930
rect 82430 24932 82630 24938
rect 82430 24898 82442 24932
rect 82618 24930 82630 24932
rect 82928 24932 83128 24938
rect 82928 24930 82940 24932
rect 82618 24900 82940 24930
rect 82618 24898 82630 24900
rect 82430 24892 82630 24898
rect 82210 24780 82280 24840
rect 82210 24520 82230 24780
rect 82270 24520 82280 24780
rect 82740 24890 82820 24900
rect 82928 24898 82940 24900
rect 83116 24898 83128 24932
rect 83160 24930 83170 24990
rect 83230 24930 83240 24990
rect 83160 24910 83240 24930
rect 82928 24892 83128 24898
rect 82740 24830 82750 24890
rect 82810 24830 82820 24890
rect 82740 24780 82820 24830
rect 82740 24720 82750 24780
rect 82810 24720 82820 24780
rect 82430 24710 82630 24716
rect 82740 24710 82820 24720
rect 83290 24840 83300 25080
rect 83340 24840 83360 25080
rect 83290 24760 83360 24840
rect 82928 24710 83128 24716
rect 82320 24680 82400 24700
rect 82320 24620 82330 24680
rect 82390 24666 82400 24680
rect 82430 24676 82442 24710
rect 82618 24680 82940 24710
rect 82618 24676 82630 24680
rect 82430 24670 82630 24676
rect 82928 24676 82940 24680
rect 83116 24676 83128 24710
rect 82928 24670 83128 24676
rect 83160 24680 83240 24700
rect 82392 24632 82400 24666
rect 82390 24620 82400 24632
rect 82320 24600 82400 24620
rect 82430 24622 82630 24628
rect 82430 24588 82442 24622
rect 82618 24620 82630 24622
rect 82928 24622 83128 24628
rect 82928 24620 82940 24622
rect 82618 24610 82940 24620
rect 82618 24590 82750 24610
rect 82618 24588 82630 24590
rect 82430 24582 82630 24588
rect 82740 24550 82750 24590
rect 82810 24590 82940 24610
rect 82810 24550 82820 24590
rect 82928 24588 82940 24590
rect 83116 24588 83128 24622
rect 83160 24620 83170 24680
rect 83230 24620 83240 24680
rect 83160 24600 83240 24620
rect 82928 24582 83128 24588
rect 82740 24540 82820 24550
rect 82210 23830 82280 24520
rect 83290 24520 83300 24760
rect 83340 24520 83360 24760
rect 83290 24110 83360 24520
rect 83270 24070 83360 24080
rect 83270 24010 83280 24070
rect 83350 24010 83360 24070
rect 83270 24000 83360 24010
rect 83290 23940 83360 24000
rect 83280 23930 83360 23940
rect 83280 23870 83290 23930
rect 83350 23870 83360 23930
rect 83280 23860 83360 23870
rect 82210 23820 83360 23830
rect 82210 23760 82220 23820
rect 82280 23770 83360 23820
rect 82280 23760 82290 23770
rect 82210 23750 82290 23760
rect 82210 23370 82280 23750
rect 82210 23130 82230 23370
rect 82270 23130 82280 23370
rect 83290 23370 83360 23770
rect 82740 23350 82820 23360
rect 82430 23310 82630 23316
rect 82740 23310 82750 23350
rect 82320 23280 82400 23300
rect 82320 23220 82330 23280
rect 82390 23266 82400 23280
rect 82430 23276 82442 23310
rect 82618 23290 82750 23310
rect 82810 23310 82820 23350
rect 82928 23310 83128 23316
rect 82810 23290 82940 23310
rect 82618 23280 82940 23290
rect 82618 23276 82630 23280
rect 82430 23270 82630 23276
rect 82928 23276 82940 23280
rect 83116 23276 83128 23310
rect 82928 23270 83128 23276
rect 83160 23280 83240 23300
rect 82392 23232 82400 23266
rect 82390 23220 82400 23232
rect 82320 23200 82400 23220
rect 82430 23222 82630 23228
rect 82430 23188 82442 23222
rect 82618 23220 82630 23222
rect 82928 23222 83128 23228
rect 82928 23220 82940 23222
rect 82618 23190 82940 23220
rect 82618 23188 82630 23190
rect 82430 23182 82630 23188
rect 82210 23070 82280 23130
rect 82210 22810 82230 23070
rect 82270 22810 82280 23070
rect 82740 23180 82820 23190
rect 82928 23188 82940 23190
rect 83116 23188 83128 23222
rect 83160 23220 83170 23280
rect 83230 23220 83240 23280
rect 83160 23200 83240 23220
rect 82928 23182 83128 23188
rect 82740 23120 82750 23180
rect 82810 23120 82820 23180
rect 82740 23070 82820 23120
rect 82740 23010 82750 23070
rect 82810 23010 82820 23070
rect 82430 23000 82630 23006
rect 82740 23000 82820 23010
rect 83290 23130 83300 23370
rect 83340 23130 83360 23370
rect 83290 23050 83360 23130
rect 82928 23000 83128 23006
rect 82320 22970 82400 22990
rect 82320 22910 82330 22970
rect 82390 22956 82400 22970
rect 82430 22966 82442 23000
rect 82618 22970 82940 23000
rect 82618 22966 82630 22970
rect 82430 22960 82630 22966
rect 82928 22966 82940 22970
rect 83116 22966 83128 23000
rect 82928 22960 83128 22966
rect 83160 22970 83240 22990
rect 82392 22922 82400 22956
rect 82390 22910 82400 22922
rect 82320 22890 82400 22910
rect 82430 22912 82630 22918
rect 82430 22878 82442 22912
rect 82618 22910 82630 22912
rect 82928 22912 83128 22918
rect 82928 22910 82940 22912
rect 82618 22900 82940 22910
rect 82618 22880 82750 22900
rect 82618 22878 82630 22880
rect 82430 22872 82630 22878
rect 82740 22840 82750 22880
rect 82810 22880 82940 22900
rect 82810 22840 82820 22880
rect 82928 22878 82940 22880
rect 83116 22878 83128 22912
rect 83160 22910 83170 22970
rect 83230 22910 83240 22970
rect 83160 22890 83240 22910
rect 82928 22872 83128 22878
rect 82740 22830 82820 22840
rect 82210 22120 82280 22810
rect 83290 22810 83300 23050
rect 83340 22810 83360 23050
rect 83290 22400 83360 22810
rect 83270 22360 83360 22370
rect 83270 22300 83280 22360
rect 83350 22300 83360 22360
rect 83270 22290 83360 22300
rect 83290 22230 83360 22290
rect 83280 22220 83360 22230
rect 83280 22160 83290 22220
rect 83350 22160 83360 22220
rect 83280 22150 83360 22160
rect 82210 22110 83360 22120
rect 82210 22050 82220 22110
rect 82280 22060 83360 22110
rect 82280 22050 82290 22060
rect 82210 22040 82290 22050
rect 82210 21660 82280 22040
rect 82210 21420 82230 21660
rect 82270 21420 82280 21660
rect 83290 21660 83360 22060
rect 82740 21640 82820 21650
rect 82430 21600 82630 21606
rect 82740 21600 82750 21640
rect 82320 21570 82400 21590
rect 82320 21510 82330 21570
rect 82390 21556 82400 21570
rect 82430 21566 82442 21600
rect 82618 21580 82750 21600
rect 82810 21600 82820 21640
rect 82928 21600 83128 21606
rect 82810 21580 82940 21600
rect 82618 21570 82940 21580
rect 82618 21566 82630 21570
rect 82430 21560 82630 21566
rect 82928 21566 82940 21570
rect 83116 21566 83128 21600
rect 82928 21560 83128 21566
rect 83160 21570 83240 21590
rect 82392 21522 82400 21556
rect 82390 21510 82400 21522
rect 82320 21490 82400 21510
rect 82430 21512 82630 21518
rect 82430 21478 82442 21512
rect 82618 21510 82630 21512
rect 82928 21512 83128 21518
rect 82928 21510 82940 21512
rect 82618 21480 82940 21510
rect 82618 21478 82630 21480
rect 82430 21472 82630 21478
rect 82210 21360 82280 21420
rect 82210 21100 82230 21360
rect 82270 21100 82280 21360
rect 82740 21470 82820 21480
rect 82928 21478 82940 21480
rect 83116 21478 83128 21512
rect 83160 21510 83170 21570
rect 83230 21510 83240 21570
rect 83160 21490 83240 21510
rect 82928 21472 83128 21478
rect 82740 21410 82750 21470
rect 82810 21410 82820 21470
rect 82740 21360 82820 21410
rect 82740 21300 82750 21360
rect 82810 21300 82820 21360
rect 82430 21290 82630 21296
rect 82740 21290 82820 21300
rect 83290 21420 83300 21660
rect 83340 21420 83360 21660
rect 83290 21340 83360 21420
rect 82928 21290 83128 21296
rect 82320 21260 82400 21280
rect 82320 21200 82330 21260
rect 82390 21246 82400 21260
rect 82430 21256 82442 21290
rect 82618 21260 82940 21290
rect 82618 21256 82630 21260
rect 82430 21250 82630 21256
rect 82928 21256 82940 21260
rect 83116 21256 83128 21290
rect 82928 21250 83128 21256
rect 83160 21260 83240 21280
rect 82392 21212 82400 21246
rect 82390 21200 82400 21212
rect 82320 21180 82400 21200
rect 82430 21202 82630 21208
rect 82430 21168 82442 21202
rect 82618 21200 82630 21202
rect 82928 21202 83128 21208
rect 82928 21200 82940 21202
rect 82618 21190 82940 21200
rect 82618 21170 82750 21190
rect 82618 21168 82630 21170
rect 82430 21162 82630 21168
rect 82740 21130 82750 21170
rect 82810 21170 82940 21190
rect 82810 21130 82820 21170
rect 82928 21168 82940 21170
rect 83116 21168 83128 21202
rect 83160 21200 83170 21260
rect 83230 21200 83240 21260
rect 83160 21180 83240 21200
rect 82928 21162 83128 21168
rect 82740 21120 82820 21130
rect 82210 20410 82280 21100
rect 83290 21100 83300 21340
rect 83340 21100 83360 21340
rect 83290 20690 83360 21100
rect 83270 20650 83360 20660
rect 83270 20590 83280 20650
rect 83350 20590 83360 20650
rect 83270 20580 83360 20590
rect 83290 20520 83360 20580
rect 83280 20510 83360 20520
rect 83280 20450 83290 20510
rect 83350 20450 83360 20510
rect 83280 20440 83360 20450
rect 82210 20400 83360 20410
rect 82210 20340 82220 20400
rect 82280 20350 83360 20400
rect 82280 20340 82290 20350
rect 82210 20330 82290 20340
rect 82210 19950 82280 20330
rect 82210 19710 82230 19950
rect 82270 19710 82280 19950
rect 83290 19950 83360 20350
rect 82740 19930 82820 19940
rect 82430 19890 82630 19896
rect 82740 19890 82750 19930
rect 82320 19860 82400 19880
rect 82320 19800 82330 19860
rect 82390 19846 82400 19860
rect 82430 19856 82442 19890
rect 82618 19870 82750 19890
rect 82810 19890 82820 19930
rect 82928 19890 83128 19896
rect 82810 19870 82940 19890
rect 82618 19860 82940 19870
rect 82618 19856 82630 19860
rect 82430 19850 82630 19856
rect 82928 19856 82940 19860
rect 83116 19856 83128 19890
rect 82928 19850 83128 19856
rect 83160 19860 83240 19880
rect 82392 19812 82400 19846
rect 82390 19800 82400 19812
rect 82320 19780 82400 19800
rect 82430 19802 82630 19808
rect 82430 19768 82442 19802
rect 82618 19800 82630 19802
rect 82928 19802 83128 19808
rect 82928 19800 82940 19802
rect 82618 19770 82940 19800
rect 82618 19768 82630 19770
rect 82430 19762 82630 19768
rect 82210 19650 82280 19710
rect 82210 19390 82230 19650
rect 82270 19390 82280 19650
rect 82740 19760 82820 19770
rect 82928 19768 82940 19770
rect 83116 19768 83128 19802
rect 83160 19800 83170 19860
rect 83230 19800 83240 19860
rect 83160 19780 83240 19800
rect 82928 19762 83128 19768
rect 82740 19700 82750 19760
rect 82810 19700 82820 19760
rect 82740 19650 82820 19700
rect 82740 19590 82750 19650
rect 82810 19590 82820 19650
rect 82430 19580 82630 19586
rect 82740 19580 82820 19590
rect 83290 19710 83300 19950
rect 83340 19710 83360 19950
rect 83290 19630 83360 19710
rect 82928 19580 83128 19586
rect 82320 19550 82400 19570
rect 82320 19490 82330 19550
rect 82390 19536 82400 19550
rect 82430 19546 82442 19580
rect 82618 19550 82940 19580
rect 82618 19546 82630 19550
rect 82430 19540 82630 19546
rect 82928 19546 82940 19550
rect 83116 19546 83128 19580
rect 82928 19540 83128 19546
rect 83160 19550 83240 19570
rect 82392 19502 82400 19536
rect 82390 19490 82400 19502
rect 82320 19470 82400 19490
rect 82430 19492 82630 19498
rect 82430 19458 82442 19492
rect 82618 19490 82630 19492
rect 82928 19492 83128 19498
rect 82928 19490 82940 19492
rect 82618 19480 82940 19490
rect 82618 19460 82750 19480
rect 82618 19458 82630 19460
rect 82430 19452 82630 19458
rect 82740 19420 82750 19460
rect 82810 19460 82940 19480
rect 82810 19420 82820 19460
rect 82928 19458 82940 19460
rect 83116 19458 83128 19492
rect 83160 19490 83170 19550
rect 83230 19490 83240 19550
rect 83160 19470 83240 19490
rect 82928 19452 83128 19458
rect 82740 19410 82820 19420
rect 82210 18700 82280 19390
rect 83290 19390 83300 19630
rect 83340 19390 83360 19630
rect 83290 18980 83360 19390
rect 83270 18940 83360 18950
rect 83270 18880 83280 18940
rect 83350 18880 83360 18940
rect 83270 18870 83360 18880
rect 83290 18810 83360 18870
rect 83280 18800 83360 18810
rect 83280 18740 83290 18800
rect 83350 18740 83360 18800
rect 83280 18730 83360 18740
rect 82210 18690 83360 18700
rect 82210 18630 82220 18690
rect 82280 18640 83360 18690
rect 82280 18630 82290 18640
rect 82210 18620 82290 18630
rect 82210 18240 82280 18620
rect 82210 18000 82230 18240
rect 82270 18000 82280 18240
rect 83290 18240 83360 18640
rect 82740 18220 82820 18230
rect 82430 18180 82630 18186
rect 82740 18180 82750 18220
rect 82320 18150 82400 18170
rect 82320 18090 82330 18150
rect 82390 18136 82400 18150
rect 82430 18146 82442 18180
rect 82618 18160 82750 18180
rect 82810 18180 82820 18220
rect 82928 18180 83128 18186
rect 82810 18160 82940 18180
rect 82618 18150 82940 18160
rect 82618 18146 82630 18150
rect 82430 18140 82630 18146
rect 82928 18146 82940 18150
rect 83116 18146 83128 18180
rect 82928 18140 83128 18146
rect 83160 18150 83240 18170
rect 82392 18102 82400 18136
rect 82390 18090 82400 18102
rect 82320 18070 82400 18090
rect 82430 18092 82630 18098
rect 82430 18058 82442 18092
rect 82618 18090 82630 18092
rect 82928 18092 83128 18098
rect 82928 18090 82940 18092
rect 82618 18060 82940 18090
rect 82618 18058 82630 18060
rect 82430 18052 82630 18058
rect 82210 17940 82280 18000
rect 82210 17680 82230 17940
rect 82270 17680 82280 17940
rect 82740 18050 82820 18060
rect 82928 18058 82940 18060
rect 83116 18058 83128 18092
rect 83160 18090 83170 18150
rect 83230 18090 83240 18150
rect 83160 18070 83240 18090
rect 82928 18052 83128 18058
rect 82740 17990 82750 18050
rect 82810 17990 82820 18050
rect 82740 17940 82820 17990
rect 82740 17880 82750 17940
rect 82810 17880 82820 17940
rect 82430 17870 82630 17876
rect 82740 17870 82820 17880
rect 83290 18000 83300 18240
rect 83340 18000 83360 18240
rect 83290 17920 83360 18000
rect 82928 17870 83128 17876
rect 82320 17840 82400 17860
rect 82320 17780 82330 17840
rect 82390 17826 82400 17840
rect 82430 17836 82442 17870
rect 82618 17840 82940 17870
rect 82618 17836 82630 17840
rect 82430 17830 82630 17836
rect 82928 17836 82940 17840
rect 83116 17836 83128 17870
rect 82928 17830 83128 17836
rect 83160 17840 83240 17860
rect 82392 17792 82400 17826
rect 82390 17780 82400 17792
rect 82320 17760 82400 17780
rect 82430 17782 82630 17788
rect 82430 17748 82442 17782
rect 82618 17780 82630 17782
rect 82928 17782 83128 17788
rect 82928 17780 82940 17782
rect 82618 17770 82940 17780
rect 82618 17750 82750 17770
rect 82618 17748 82630 17750
rect 82430 17742 82630 17748
rect 82740 17710 82750 17750
rect 82810 17750 82940 17770
rect 82810 17710 82820 17750
rect 82928 17748 82940 17750
rect 83116 17748 83128 17782
rect 83160 17780 83170 17840
rect 83230 17780 83240 17840
rect 83160 17760 83240 17780
rect 82928 17742 83128 17748
rect 82740 17700 82820 17710
rect 82210 16990 82280 17680
rect 83290 17680 83300 17920
rect 83340 17680 83360 17920
rect 83290 17270 83360 17680
rect 83270 17230 83360 17240
rect 83270 17170 83280 17230
rect 83350 17170 83360 17230
rect 83270 17160 83360 17170
rect 83290 17100 83360 17160
rect 83280 17090 83360 17100
rect 83280 17030 83290 17090
rect 83350 17030 83360 17090
rect 83280 17020 83360 17030
rect 82210 16980 83360 16990
rect 82210 16920 82220 16980
rect 82280 16930 83360 16980
rect 82280 16920 82290 16930
rect 82210 16910 82290 16920
rect 82210 16530 82280 16910
rect 82210 16290 82230 16530
rect 82270 16290 82280 16530
rect 83290 16530 83360 16930
rect 82740 16510 82820 16520
rect 82430 16470 82630 16476
rect 82740 16470 82750 16510
rect 82320 16440 82400 16460
rect 82320 16380 82330 16440
rect 82390 16426 82400 16440
rect 82430 16436 82442 16470
rect 82618 16450 82750 16470
rect 82810 16470 82820 16510
rect 82928 16470 83128 16476
rect 82810 16450 82940 16470
rect 82618 16440 82940 16450
rect 82618 16436 82630 16440
rect 82430 16430 82630 16436
rect 82928 16436 82940 16440
rect 83116 16436 83128 16470
rect 82928 16430 83128 16436
rect 83160 16440 83240 16460
rect 82392 16392 82400 16426
rect 82390 16380 82400 16392
rect 82320 16360 82400 16380
rect 82430 16382 82630 16388
rect 82430 16348 82442 16382
rect 82618 16380 82630 16382
rect 82928 16382 83128 16388
rect 82928 16380 82940 16382
rect 82618 16350 82940 16380
rect 82618 16348 82630 16350
rect 82430 16342 82630 16348
rect 82210 16230 82280 16290
rect 82210 15970 82230 16230
rect 82270 15970 82280 16230
rect 82740 16340 82820 16350
rect 82928 16348 82940 16350
rect 83116 16348 83128 16382
rect 83160 16380 83170 16440
rect 83230 16380 83240 16440
rect 83160 16360 83240 16380
rect 82928 16342 83128 16348
rect 82740 16280 82750 16340
rect 82810 16280 82820 16340
rect 82740 16230 82820 16280
rect 82740 16170 82750 16230
rect 82810 16170 82820 16230
rect 82430 16160 82630 16166
rect 82740 16160 82820 16170
rect 83290 16290 83300 16530
rect 83340 16290 83360 16530
rect 83290 16210 83360 16290
rect 82928 16160 83128 16166
rect 82320 16130 82400 16150
rect 82320 16070 82330 16130
rect 82390 16116 82400 16130
rect 82430 16126 82442 16160
rect 82618 16130 82940 16160
rect 82618 16126 82630 16130
rect 82430 16120 82630 16126
rect 82928 16126 82940 16130
rect 83116 16126 83128 16160
rect 82928 16120 83128 16126
rect 83160 16130 83240 16150
rect 82392 16082 82400 16116
rect 82390 16070 82400 16082
rect 82320 16050 82400 16070
rect 82430 16072 82630 16078
rect 82430 16038 82442 16072
rect 82618 16070 82630 16072
rect 82928 16072 83128 16078
rect 82928 16070 82940 16072
rect 82618 16060 82940 16070
rect 82618 16040 82750 16060
rect 82618 16038 82630 16040
rect 82430 16032 82630 16038
rect 82740 16000 82750 16040
rect 82810 16040 82940 16060
rect 82810 16000 82820 16040
rect 82928 16038 82940 16040
rect 83116 16038 83128 16072
rect 83160 16070 83170 16130
rect 83230 16070 83240 16130
rect 83160 16050 83240 16070
rect 82928 16032 83128 16038
rect 82740 15990 82820 16000
rect 82210 15280 82280 15970
rect 83290 15970 83300 16210
rect 83340 15970 83360 16210
rect 83290 15560 83360 15970
rect 83270 15520 83360 15530
rect 83270 15460 83280 15520
rect 83350 15460 83360 15520
rect 83270 15450 83360 15460
rect 83290 15390 83360 15450
rect 83280 15380 83360 15390
rect 83280 15320 83290 15380
rect 83350 15320 83360 15380
rect 83280 15310 83360 15320
rect 82210 15270 83360 15280
rect 82210 15210 82220 15270
rect 82280 15220 83360 15270
rect 82280 15210 82290 15220
rect 82210 15200 82290 15210
rect 82210 14820 82280 15200
rect 82210 14580 82230 14820
rect 82270 14580 82280 14820
rect 83290 14820 83360 15220
rect 82740 14800 82820 14810
rect 82430 14760 82630 14766
rect 82740 14760 82750 14800
rect 82320 14730 82400 14750
rect 82320 14670 82330 14730
rect 82390 14716 82400 14730
rect 82430 14726 82442 14760
rect 82618 14740 82750 14760
rect 82810 14760 82820 14800
rect 82928 14760 83128 14766
rect 82810 14740 82940 14760
rect 82618 14730 82940 14740
rect 82618 14726 82630 14730
rect 82430 14720 82630 14726
rect 82928 14726 82940 14730
rect 83116 14726 83128 14760
rect 82928 14720 83128 14726
rect 83160 14730 83240 14750
rect 82392 14682 82400 14716
rect 82390 14670 82400 14682
rect 82320 14650 82400 14670
rect 82430 14672 82630 14678
rect 82430 14638 82442 14672
rect 82618 14670 82630 14672
rect 82928 14672 83128 14678
rect 82928 14670 82940 14672
rect 82618 14640 82940 14670
rect 82618 14638 82630 14640
rect 82430 14632 82630 14638
rect 82210 14520 82280 14580
rect 82210 14260 82230 14520
rect 82270 14260 82280 14520
rect 82740 14630 82820 14640
rect 82928 14638 82940 14640
rect 83116 14638 83128 14672
rect 83160 14670 83170 14730
rect 83230 14670 83240 14730
rect 83160 14650 83240 14670
rect 82928 14632 83128 14638
rect 82740 14570 82750 14630
rect 82810 14570 82820 14630
rect 82740 14520 82820 14570
rect 82740 14460 82750 14520
rect 82810 14460 82820 14520
rect 82430 14450 82630 14456
rect 82740 14450 82820 14460
rect 83290 14580 83300 14820
rect 83340 14580 83360 14820
rect 83290 14500 83360 14580
rect 82928 14450 83128 14456
rect 82320 14420 82400 14440
rect 82320 14360 82330 14420
rect 82390 14406 82400 14420
rect 82430 14416 82442 14450
rect 82618 14420 82940 14450
rect 82618 14416 82630 14420
rect 82430 14410 82630 14416
rect 82928 14416 82940 14420
rect 83116 14416 83128 14450
rect 82928 14410 83128 14416
rect 83160 14420 83240 14440
rect 82392 14372 82400 14406
rect 82390 14360 82400 14372
rect 82320 14340 82400 14360
rect 82430 14362 82630 14368
rect 82430 14328 82442 14362
rect 82618 14360 82630 14362
rect 82928 14362 83128 14368
rect 82928 14360 82940 14362
rect 82618 14350 82940 14360
rect 82618 14330 82750 14350
rect 82618 14328 82630 14330
rect 82430 14322 82630 14328
rect 82740 14290 82750 14330
rect 82810 14330 82940 14350
rect 82810 14290 82820 14330
rect 82928 14328 82940 14330
rect 83116 14328 83128 14362
rect 83160 14360 83170 14420
rect 83230 14360 83240 14420
rect 83160 14340 83240 14360
rect 82928 14322 83128 14328
rect 82740 14280 82820 14290
rect 82210 13570 82280 14260
rect 83290 14260 83300 14500
rect 83340 14260 83360 14500
rect 83290 13850 83360 14260
rect 83270 13810 83360 13820
rect 83270 13750 83280 13810
rect 83350 13750 83360 13810
rect 83270 13740 83360 13750
rect 83290 13680 83360 13740
rect 83280 13670 83360 13680
rect 83280 13610 83290 13670
rect 83350 13610 83360 13670
rect 83280 13600 83360 13610
rect 82210 13560 83360 13570
rect 82210 13500 82220 13560
rect 82280 13510 83360 13560
rect 82280 13500 82290 13510
rect 82210 13490 82290 13500
rect 82210 13110 82280 13490
rect 82210 12870 82230 13110
rect 82270 12870 82280 13110
rect 83290 13110 83360 13510
rect 82740 13090 82820 13100
rect 82430 13050 82630 13056
rect 82740 13050 82750 13090
rect 82320 13020 82400 13040
rect 82320 12960 82330 13020
rect 82390 13006 82400 13020
rect 82430 13016 82442 13050
rect 82618 13030 82750 13050
rect 82810 13050 82820 13090
rect 82928 13050 83128 13056
rect 82810 13030 82940 13050
rect 82618 13020 82940 13030
rect 82618 13016 82630 13020
rect 82430 13010 82630 13016
rect 82928 13016 82940 13020
rect 83116 13016 83128 13050
rect 82928 13010 83128 13016
rect 83160 13020 83240 13040
rect 82392 12972 82400 13006
rect 82390 12960 82400 12972
rect 82320 12940 82400 12960
rect 82430 12962 82630 12968
rect 82430 12928 82442 12962
rect 82618 12960 82630 12962
rect 82928 12962 83128 12968
rect 82928 12960 82940 12962
rect 82618 12930 82940 12960
rect 82618 12928 82630 12930
rect 82430 12922 82630 12928
rect 82210 12810 82280 12870
rect 82210 12550 82230 12810
rect 82270 12550 82280 12810
rect 82740 12920 82820 12930
rect 82928 12928 82940 12930
rect 83116 12928 83128 12962
rect 83160 12960 83170 13020
rect 83230 12960 83240 13020
rect 83160 12940 83240 12960
rect 82928 12922 83128 12928
rect 82740 12860 82750 12920
rect 82810 12860 82820 12920
rect 82740 12810 82820 12860
rect 82740 12750 82750 12810
rect 82810 12750 82820 12810
rect 82430 12740 82630 12746
rect 82740 12740 82820 12750
rect 83290 12870 83300 13110
rect 83340 12870 83360 13110
rect 83290 12790 83360 12870
rect 82928 12740 83128 12746
rect 82320 12710 82400 12730
rect 82320 12650 82330 12710
rect 82390 12696 82400 12710
rect 82430 12706 82442 12740
rect 82618 12710 82940 12740
rect 82618 12706 82630 12710
rect 82430 12700 82630 12706
rect 82928 12706 82940 12710
rect 83116 12706 83128 12740
rect 82928 12700 83128 12706
rect 83160 12710 83240 12730
rect 82392 12662 82400 12696
rect 82390 12650 82400 12662
rect 82320 12630 82400 12650
rect 82430 12652 82630 12658
rect 82430 12618 82442 12652
rect 82618 12650 82630 12652
rect 82928 12652 83128 12658
rect 82928 12650 82940 12652
rect 82618 12640 82940 12650
rect 82618 12620 82750 12640
rect 82618 12618 82630 12620
rect 82430 12612 82630 12618
rect 82740 12580 82750 12620
rect 82810 12620 82940 12640
rect 82810 12580 82820 12620
rect 82928 12618 82940 12620
rect 83116 12618 83128 12652
rect 83160 12650 83170 12710
rect 83230 12650 83240 12710
rect 83160 12630 83240 12650
rect 82928 12612 83128 12618
rect 82740 12570 82820 12580
rect 82210 11860 82280 12550
rect 83290 12550 83300 12790
rect 83340 12550 83360 12790
rect 83290 12140 83360 12550
rect 83270 12100 83360 12110
rect 83270 12040 83280 12100
rect 83350 12040 83360 12100
rect 83270 12030 83360 12040
rect 83290 11970 83360 12030
rect 83280 11960 83360 11970
rect 83280 11900 83290 11960
rect 83350 11900 83360 11960
rect 83280 11890 83360 11900
rect 82210 11850 83360 11860
rect 82210 11790 82220 11850
rect 82280 11800 83360 11850
rect 82280 11790 82290 11800
rect 82210 11780 82290 11790
rect 82210 11400 82280 11780
rect 82210 11160 82230 11400
rect 82270 11160 82280 11400
rect 83290 11400 83360 11800
rect 82740 11380 82820 11390
rect 82430 11340 82630 11346
rect 82740 11340 82750 11380
rect 82320 11310 82400 11330
rect 82320 11250 82330 11310
rect 82390 11296 82400 11310
rect 82430 11306 82442 11340
rect 82618 11320 82750 11340
rect 82810 11340 82820 11380
rect 82928 11340 83128 11346
rect 82810 11320 82940 11340
rect 82618 11310 82940 11320
rect 82618 11306 82630 11310
rect 82430 11300 82630 11306
rect 82928 11306 82940 11310
rect 83116 11306 83128 11340
rect 82928 11300 83128 11306
rect 83160 11310 83240 11330
rect 82392 11262 82400 11296
rect 82390 11250 82400 11262
rect 82320 11230 82400 11250
rect 82430 11252 82630 11258
rect 82430 11218 82442 11252
rect 82618 11250 82630 11252
rect 82928 11252 83128 11258
rect 82928 11250 82940 11252
rect 82618 11220 82940 11250
rect 82618 11218 82630 11220
rect 82430 11212 82630 11218
rect 82210 11100 82280 11160
rect 82210 10840 82230 11100
rect 82270 10840 82280 11100
rect 82740 11210 82820 11220
rect 82928 11218 82940 11220
rect 83116 11218 83128 11252
rect 83160 11250 83170 11310
rect 83230 11250 83240 11310
rect 83160 11230 83240 11250
rect 82928 11212 83128 11218
rect 82740 11150 82750 11210
rect 82810 11150 82820 11210
rect 82740 11100 82820 11150
rect 82740 11040 82750 11100
rect 82810 11040 82820 11100
rect 82430 11030 82630 11036
rect 82740 11030 82820 11040
rect 83290 11160 83300 11400
rect 83340 11160 83360 11400
rect 83290 11080 83360 11160
rect 82928 11030 83128 11036
rect 82320 11000 82400 11020
rect 82320 10940 82330 11000
rect 82390 10986 82400 11000
rect 82430 10996 82442 11030
rect 82618 11000 82940 11030
rect 82618 10996 82630 11000
rect 82430 10990 82630 10996
rect 82928 10996 82940 11000
rect 83116 10996 83128 11030
rect 82928 10990 83128 10996
rect 83160 11000 83240 11020
rect 82392 10952 82400 10986
rect 82390 10940 82400 10952
rect 82320 10920 82400 10940
rect 82430 10942 82630 10948
rect 82430 10908 82442 10942
rect 82618 10940 82630 10942
rect 82928 10942 83128 10948
rect 82928 10940 82940 10942
rect 82618 10930 82940 10940
rect 82618 10910 82750 10930
rect 82618 10908 82630 10910
rect 82430 10902 82630 10908
rect 82740 10870 82750 10910
rect 82810 10910 82940 10930
rect 82810 10870 82820 10910
rect 82928 10908 82940 10910
rect 83116 10908 83128 10942
rect 83160 10940 83170 11000
rect 83230 10940 83240 11000
rect 83160 10920 83240 10940
rect 82928 10902 83128 10908
rect 82740 10860 82820 10870
rect 82210 10150 82280 10840
rect 83290 10840 83300 11080
rect 83340 10840 83360 11080
rect 83290 10430 83360 10840
rect 83270 10390 83360 10400
rect 83270 10330 83280 10390
rect 83350 10330 83360 10390
rect 83270 10320 83360 10330
rect 83290 10260 83360 10320
rect 83280 10250 83360 10260
rect 83280 10190 83290 10250
rect 83350 10190 83360 10250
rect 83280 10180 83360 10190
rect 82210 10140 83360 10150
rect 82210 10080 82220 10140
rect 82280 10090 83360 10140
rect 82280 10080 82290 10090
rect 82210 10070 82290 10080
rect 82210 9690 82280 10070
rect 82210 9450 82230 9690
rect 82270 9450 82280 9690
rect 83290 9690 83360 10090
rect 82740 9670 82820 9680
rect 82430 9630 82630 9636
rect 82740 9630 82750 9670
rect 82320 9600 82400 9620
rect 82320 9540 82330 9600
rect 82390 9586 82400 9600
rect 82430 9596 82442 9630
rect 82618 9610 82750 9630
rect 82810 9630 82820 9670
rect 82928 9630 83128 9636
rect 82810 9610 82940 9630
rect 82618 9600 82940 9610
rect 82618 9596 82630 9600
rect 82430 9590 82630 9596
rect 82928 9596 82940 9600
rect 83116 9596 83128 9630
rect 82928 9590 83128 9596
rect 83160 9600 83240 9620
rect 82392 9552 82400 9586
rect 82390 9540 82400 9552
rect 82320 9520 82400 9540
rect 82430 9542 82630 9548
rect 82430 9508 82442 9542
rect 82618 9540 82630 9542
rect 82928 9542 83128 9548
rect 82928 9540 82940 9542
rect 82618 9510 82940 9540
rect 82618 9508 82630 9510
rect 82430 9502 82630 9508
rect 82210 9390 82280 9450
rect 82210 9130 82230 9390
rect 82270 9130 82280 9390
rect 82740 9500 82820 9510
rect 82928 9508 82940 9510
rect 83116 9508 83128 9542
rect 83160 9540 83170 9600
rect 83230 9540 83240 9600
rect 83160 9520 83240 9540
rect 82928 9502 83128 9508
rect 82740 9440 82750 9500
rect 82810 9440 82820 9500
rect 82740 9390 82820 9440
rect 82740 9330 82750 9390
rect 82810 9330 82820 9390
rect 82430 9320 82630 9326
rect 82740 9320 82820 9330
rect 83290 9450 83300 9690
rect 83340 9450 83360 9690
rect 83290 9370 83360 9450
rect 82928 9320 83128 9326
rect 82320 9290 82400 9310
rect 82320 9230 82330 9290
rect 82390 9276 82400 9290
rect 82430 9286 82442 9320
rect 82618 9290 82940 9320
rect 82618 9286 82630 9290
rect 82430 9280 82630 9286
rect 82928 9286 82940 9290
rect 83116 9286 83128 9320
rect 82928 9280 83128 9286
rect 83160 9290 83240 9310
rect 82392 9242 82400 9276
rect 82390 9230 82400 9242
rect 82320 9210 82400 9230
rect 82430 9232 82630 9238
rect 82430 9198 82442 9232
rect 82618 9230 82630 9232
rect 82928 9232 83128 9238
rect 82928 9230 82940 9232
rect 82618 9220 82940 9230
rect 82618 9200 82750 9220
rect 82618 9198 82630 9200
rect 82430 9192 82630 9198
rect 82740 9160 82750 9200
rect 82810 9200 82940 9220
rect 82810 9160 82820 9200
rect 82928 9198 82940 9200
rect 83116 9198 83128 9232
rect 83160 9230 83170 9290
rect 83230 9230 83240 9290
rect 83160 9210 83240 9230
rect 82928 9192 83128 9198
rect 82740 9150 82820 9160
rect 82210 8440 82280 9130
rect 83290 9130 83300 9370
rect 83340 9130 83360 9370
rect 83290 8720 83360 9130
rect 83270 8680 83360 8690
rect 83270 8620 83280 8680
rect 83350 8620 83360 8680
rect 83270 8610 83360 8620
rect 83290 8550 83360 8610
rect 83280 8540 83360 8550
rect 83280 8480 83290 8540
rect 83350 8480 83360 8540
rect 83280 8470 83360 8480
rect 82210 8430 83360 8440
rect 82210 8370 82220 8430
rect 82280 8380 83360 8430
rect 82280 8370 82290 8380
rect 82210 8360 82290 8370
rect 82210 7980 82280 8360
rect 82210 7740 82230 7980
rect 82270 7740 82280 7980
rect 83290 7980 83360 8380
rect 82740 7960 82820 7970
rect 82430 7920 82630 7926
rect 82740 7920 82750 7960
rect 82320 7890 82400 7910
rect 82320 7830 82330 7890
rect 82390 7876 82400 7890
rect 82430 7886 82442 7920
rect 82618 7900 82750 7920
rect 82810 7920 82820 7960
rect 82928 7920 83128 7926
rect 82810 7900 82940 7920
rect 82618 7890 82940 7900
rect 82618 7886 82630 7890
rect 82430 7880 82630 7886
rect 82928 7886 82940 7890
rect 83116 7886 83128 7920
rect 82928 7880 83128 7886
rect 83160 7890 83240 7910
rect 82392 7842 82400 7876
rect 82390 7830 82400 7842
rect 82320 7810 82400 7830
rect 82430 7832 82630 7838
rect 82430 7798 82442 7832
rect 82618 7830 82630 7832
rect 82928 7832 83128 7838
rect 82928 7830 82940 7832
rect 82618 7800 82940 7830
rect 82618 7798 82630 7800
rect 82430 7792 82630 7798
rect 82210 7680 82280 7740
rect 82210 7420 82230 7680
rect 82270 7420 82280 7680
rect 82740 7790 82820 7800
rect 82928 7798 82940 7800
rect 83116 7798 83128 7832
rect 83160 7830 83170 7890
rect 83230 7830 83240 7890
rect 83160 7810 83240 7830
rect 82928 7792 83128 7798
rect 82740 7730 82750 7790
rect 82810 7730 82820 7790
rect 82740 7680 82820 7730
rect 82740 7620 82750 7680
rect 82810 7620 82820 7680
rect 82430 7610 82630 7616
rect 82740 7610 82820 7620
rect 83290 7740 83300 7980
rect 83340 7740 83360 7980
rect 83290 7660 83360 7740
rect 82928 7610 83128 7616
rect 82320 7580 82400 7600
rect 82320 7520 82330 7580
rect 82390 7566 82400 7580
rect 82430 7576 82442 7610
rect 82618 7580 82940 7610
rect 82618 7576 82630 7580
rect 82430 7570 82630 7576
rect 82928 7576 82940 7580
rect 83116 7576 83128 7610
rect 82928 7570 83128 7576
rect 83160 7580 83240 7600
rect 82392 7532 82400 7566
rect 82390 7520 82400 7532
rect 82320 7500 82400 7520
rect 82430 7522 82630 7528
rect 82430 7488 82442 7522
rect 82618 7520 82630 7522
rect 82928 7522 83128 7528
rect 82928 7520 82940 7522
rect 82618 7510 82940 7520
rect 82618 7490 82750 7510
rect 82618 7488 82630 7490
rect 82430 7482 82630 7488
rect 82740 7450 82750 7490
rect 82810 7490 82940 7510
rect 82810 7450 82820 7490
rect 82928 7488 82940 7490
rect 83116 7488 83128 7522
rect 83160 7520 83170 7580
rect 83230 7520 83240 7580
rect 83160 7500 83240 7520
rect 82928 7482 83128 7488
rect 82740 7440 82820 7450
rect 82210 6730 82280 7420
rect 83290 7420 83300 7660
rect 83340 7420 83360 7660
rect 83290 7010 83360 7420
rect 83270 6970 83360 6980
rect 83270 6910 83280 6970
rect 83350 6910 83360 6970
rect 83270 6900 83360 6910
rect 83290 6840 83360 6900
rect 83280 6830 83360 6840
rect 83280 6770 83290 6830
rect 83350 6770 83360 6830
rect 83280 6760 83360 6770
rect 82210 6720 83360 6730
rect 82210 6660 82220 6720
rect 82280 6670 83360 6720
rect 82280 6660 82290 6670
rect 82210 6650 82290 6660
rect 82210 6270 82280 6650
rect 82210 6030 82230 6270
rect 82270 6030 82280 6270
rect 83290 6270 83360 6670
rect 82740 6250 82820 6260
rect 82430 6210 82630 6216
rect 82740 6210 82750 6250
rect 82320 6180 82400 6200
rect 82320 6120 82330 6180
rect 82390 6166 82400 6180
rect 82430 6176 82442 6210
rect 82618 6190 82750 6210
rect 82810 6210 82820 6250
rect 82928 6210 83128 6216
rect 82810 6190 82940 6210
rect 82618 6180 82940 6190
rect 82618 6176 82630 6180
rect 82430 6170 82630 6176
rect 82928 6176 82940 6180
rect 83116 6176 83128 6210
rect 82928 6170 83128 6176
rect 83160 6180 83240 6200
rect 82392 6132 82400 6166
rect 82390 6120 82400 6132
rect 82320 6100 82400 6120
rect 82430 6122 82630 6128
rect 82430 6088 82442 6122
rect 82618 6120 82630 6122
rect 82928 6122 83128 6128
rect 82928 6120 82940 6122
rect 82618 6090 82940 6120
rect 82618 6088 82630 6090
rect 82430 6082 82630 6088
rect 82210 5970 82280 6030
rect 82210 5710 82230 5970
rect 82270 5710 82280 5970
rect 82740 6080 82820 6090
rect 82928 6088 82940 6090
rect 83116 6088 83128 6122
rect 83160 6120 83170 6180
rect 83230 6120 83240 6180
rect 83160 6100 83240 6120
rect 82928 6082 83128 6088
rect 82740 6020 82750 6080
rect 82810 6020 82820 6080
rect 82740 5970 82820 6020
rect 82740 5910 82750 5970
rect 82810 5910 82820 5970
rect 82430 5900 82630 5906
rect 82740 5900 82820 5910
rect 83290 6030 83300 6270
rect 83340 6030 83360 6270
rect 83290 5950 83360 6030
rect 82928 5900 83128 5906
rect 82320 5870 82400 5890
rect 82320 5810 82330 5870
rect 82390 5856 82400 5870
rect 82430 5866 82442 5900
rect 82618 5870 82940 5900
rect 82618 5866 82630 5870
rect 82430 5860 82630 5866
rect 82928 5866 82940 5870
rect 83116 5866 83128 5900
rect 82928 5860 83128 5866
rect 83160 5870 83240 5890
rect 82392 5822 82400 5856
rect 82390 5810 82400 5822
rect 82320 5790 82400 5810
rect 82430 5812 82630 5818
rect 82430 5778 82442 5812
rect 82618 5810 82630 5812
rect 82928 5812 83128 5818
rect 82928 5810 82940 5812
rect 82618 5800 82940 5810
rect 82618 5780 82750 5800
rect 82618 5778 82630 5780
rect 82430 5772 82630 5778
rect 82740 5740 82750 5780
rect 82810 5780 82940 5800
rect 82810 5740 82820 5780
rect 82928 5778 82940 5780
rect 83116 5778 83128 5812
rect 83160 5810 83170 5870
rect 83230 5810 83240 5870
rect 83160 5790 83240 5810
rect 82928 5772 83128 5778
rect 82740 5730 82820 5740
rect 82210 5020 82280 5710
rect 83290 5710 83300 5950
rect 83340 5710 83360 5950
rect 83290 5300 83360 5710
rect 83270 5260 83360 5270
rect 83270 5200 83280 5260
rect 83350 5200 83360 5260
rect 83270 5190 83360 5200
rect 83290 5130 83360 5190
rect 83280 5120 83360 5130
rect 83280 5060 83290 5120
rect 83350 5060 83360 5120
rect 83280 5050 83360 5060
rect 82210 5010 83360 5020
rect 82210 4950 82220 5010
rect 82280 4960 83360 5010
rect 82280 4950 82290 4960
rect 82210 4940 82290 4950
rect 82210 4560 82280 4940
rect 82210 4320 82230 4560
rect 82270 4320 82280 4560
rect 83290 4560 83360 4960
rect 82740 4540 82820 4550
rect 82430 4500 82630 4506
rect 82740 4500 82750 4540
rect 82320 4470 82400 4490
rect 82320 4410 82330 4470
rect 82390 4456 82400 4470
rect 82430 4466 82442 4500
rect 82618 4480 82750 4500
rect 82810 4500 82820 4540
rect 82928 4500 83128 4506
rect 82810 4480 82940 4500
rect 82618 4470 82940 4480
rect 82618 4466 82630 4470
rect 82430 4460 82630 4466
rect 82928 4466 82940 4470
rect 83116 4466 83128 4500
rect 82928 4460 83128 4466
rect 83160 4470 83240 4490
rect 82392 4422 82400 4456
rect 82390 4410 82400 4422
rect 82320 4390 82400 4410
rect 82430 4412 82630 4418
rect 82430 4378 82442 4412
rect 82618 4410 82630 4412
rect 82928 4412 83128 4418
rect 82928 4410 82940 4412
rect 82618 4380 82940 4410
rect 82618 4378 82630 4380
rect 82430 4372 82630 4378
rect 82210 4260 82280 4320
rect 82210 4000 82230 4260
rect 82270 4000 82280 4260
rect 82740 4370 82820 4380
rect 82928 4378 82940 4380
rect 83116 4378 83128 4412
rect 83160 4410 83170 4470
rect 83230 4410 83240 4470
rect 83160 4390 83240 4410
rect 82928 4372 83128 4378
rect 82740 4310 82750 4370
rect 82810 4310 82820 4370
rect 82740 4260 82820 4310
rect 82740 4200 82750 4260
rect 82810 4200 82820 4260
rect 82430 4190 82630 4196
rect 82740 4190 82820 4200
rect 83290 4320 83300 4560
rect 83340 4320 83360 4560
rect 83290 4240 83360 4320
rect 82928 4190 83128 4196
rect 82320 4160 82400 4180
rect 82320 4100 82330 4160
rect 82390 4146 82400 4160
rect 82430 4156 82442 4190
rect 82618 4160 82940 4190
rect 82618 4156 82630 4160
rect 82430 4150 82630 4156
rect 82928 4156 82940 4160
rect 83116 4156 83128 4190
rect 82928 4150 83128 4156
rect 83160 4160 83240 4180
rect 82392 4112 82400 4146
rect 82390 4100 82400 4112
rect 82320 4080 82400 4100
rect 82430 4102 82630 4108
rect 82430 4068 82442 4102
rect 82618 4100 82630 4102
rect 82928 4102 83128 4108
rect 82928 4100 82940 4102
rect 82618 4090 82940 4100
rect 82618 4070 82750 4090
rect 82618 4068 82630 4070
rect 82430 4062 82630 4068
rect 82740 4030 82750 4070
rect 82810 4070 82940 4090
rect 82810 4030 82820 4070
rect 82928 4068 82940 4070
rect 83116 4068 83128 4102
rect 83160 4100 83170 4160
rect 83230 4100 83240 4160
rect 83160 4080 83240 4100
rect 82928 4062 83128 4068
rect 82740 4020 82820 4030
rect 82210 3310 82280 4000
rect 83290 4000 83300 4240
rect 83340 4000 83360 4240
rect 83290 3590 83360 4000
rect 83270 3550 83360 3560
rect 83270 3490 83280 3550
rect 83350 3490 83360 3550
rect 83270 3480 83360 3490
rect 83290 3420 83360 3480
rect 83280 3410 83360 3420
rect 83280 3350 83290 3410
rect 83350 3350 83360 3410
rect 83280 3340 83360 3350
rect 82210 3300 83360 3310
rect 82210 3240 82220 3300
rect 82280 3250 83360 3300
rect 82280 3240 82290 3250
rect 82210 3230 82290 3240
rect 82210 2850 82280 3230
rect 82210 2610 82230 2850
rect 82270 2610 82280 2850
rect 83290 2850 83360 3250
rect 82740 2830 82820 2840
rect 82430 2790 82630 2796
rect 82740 2790 82750 2830
rect 82320 2760 82400 2780
rect 82320 2700 82330 2760
rect 82390 2746 82400 2760
rect 82430 2756 82442 2790
rect 82618 2770 82750 2790
rect 82810 2790 82820 2830
rect 82928 2790 83128 2796
rect 82810 2770 82940 2790
rect 82618 2760 82940 2770
rect 82618 2756 82630 2760
rect 82430 2750 82630 2756
rect 82928 2756 82940 2760
rect 83116 2756 83128 2790
rect 82928 2750 83128 2756
rect 83160 2760 83240 2780
rect 82392 2712 82400 2746
rect 82390 2700 82400 2712
rect 82320 2680 82400 2700
rect 82430 2702 82630 2708
rect 82430 2668 82442 2702
rect 82618 2700 82630 2702
rect 82928 2702 83128 2708
rect 82928 2700 82940 2702
rect 82618 2670 82940 2700
rect 82618 2668 82630 2670
rect 82430 2662 82630 2668
rect 82210 2550 82280 2610
rect 82210 2290 82230 2550
rect 82270 2290 82280 2550
rect 82740 2660 82820 2670
rect 82928 2668 82940 2670
rect 83116 2668 83128 2702
rect 83160 2700 83170 2760
rect 83230 2700 83240 2760
rect 83160 2680 83240 2700
rect 82928 2662 83128 2668
rect 82740 2600 82750 2660
rect 82810 2600 82820 2660
rect 82740 2550 82820 2600
rect 82740 2490 82750 2550
rect 82810 2490 82820 2550
rect 82430 2480 82630 2486
rect 82740 2480 82820 2490
rect 83290 2610 83300 2850
rect 83340 2610 83360 2850
rect 83290 2530 83360 2610
rect 82928 2480 83128 2486
rect 82320 2450 82400 2470
rect 82320 2390 82330 2450
rect 82390 2436 82400 2450
rect 82430 2446 82442 2480
rect 82618 2450 82940 2480
rect 82618 2446 82630 2450
rect 82430 2440 82630 2446
rect 82928 2446 82940 2450
rect 83116 2446 83128 2480
rect 82928 2440 83128 2446
rect 83160 2450 83240 2470
rect 82392 2402 82400 2436
rect 82390 2390 82400 2402
rect 82320 2370 82400 2390
rect 82430 2392 82630 2398
rect 82430 2358 82442 2392
rect 82618 2390 82630 2392
rect 82928 2392 83128 2398
rect 82928 2390 82940 2392
rect 82618 2380 82940 2390
rect 82618 2360 82750 2380
rect 82618 2358 82630 2360
rect 82430 2352 82630 2358
rect 82740 2320 82750 2360
rect 82810 2360 82940 2380
rect 82810 2320 82820 2360
rect 82928 2358 82940 2360
rect 83116 2358 83128 2392
rect 83160 2390 83170 2450
rect 83230 2390 83240 2450
rect 83160 2370 83240 2390
rect 82928 2352 83128 2358
rect 82740 2310 82820 2320
rect 82210 1600 82280 2290
rect 83290 2290 83300 2530
rect 83340 2290 83360 2530
rect 83290 1880 83360 2290
rect 83270 1840 83360 1850
rect 83270 1780 83280 1840
rect 83350 1780 83360 1840
rect 83270 1770 83360 1780
rect 83290 1710 83360 1770
rect 83280 1700 83360 1710
rect 83280 1640 83290 1700
rect 83350 1640 83360 1700
rect 83280 1630 83360 1640
rect 82210 1590 83360 1600
rect 82210 1530 82220 1590
rect 82280 1540 83360 1590
rect 82280 1530 82290 1540
rect 82210 1520 82290 1530
rect 82210 1140 82280 1520
rect 82210 900 82230 1140
rect 82270 900 82280 1140
rect 83290 1140 83360 1540
rect 82740 1120 82820 1130
rect 82430 1080 82630 1086
rect 82740 1080 82750 1120
rect 82320 1050 82400 1070
rect 82320 990 82330 1050
rect 82390 1036 82400 1050
rect 82430 1046 82442 1080
rect 82618 1060 82750 1080
rect 82810 1080 82820 1120
rect 82928 1080 83128 1086
rect 82810 1060 82940 1080
rect 82618 1050 82940 1060
rect 82618 1046 82630 1050
rect 82430 1040 82630 1046
rect 82928 1046 82940 1050
rect 83116 1046 83128 1080
rect 82928 1040 83128 1046
rect 83160 1050 83240 1070
rect 82392 1002 82400 1036
rect 82390 990 82400 1002
rect 82320 970 82400 990
rect 82430 992 82630 998
rect 82430 958 82442 992
rect 82618 990 82630 992
rect 82928 992 83128 998
rect 82928 990 82940 992
rect 82618 960 82940 990
rect 82618 958 82630 960
rect 82430 952 82630 958
rect 82210 840 82280 900
rect 82210 580 82230 840
rect 82270 580 82280 840
rect 82740 950 82820 960
rect 82928 958 82940 960
rect 83116 958 83128 992
rect 83160 990 83170 1050
rect 83230 990 83240 1050
rect 83160 970 83240 990
rect 82928 952 83128 958
rect 82740 890 82750 950
rect 82810 890 82820 950
rect 82740 840 82820 890
rect 82740 780 82750 840
rect 82810 780 82820 840
rect 82430 770 82630 776
rect 82740 770 82820 780
rect 83290 900 83300 1140
rect 83340 900 83360 1140
rect 83290 820 83360 900
rect 82928 770 83128 776
rect 82320 740 82400 760
rect 82320 680 82330 740
rect 82390 726 82400 740
rect 82430 736 82442 770
rect 82618 740 82940 770
rect 82618 736 82630 740
rect 82430 730 82630 736
rect 82928 736 82940 740
rect 83116 736 83128 770
rect 82928 730 83128 736
rect 83160 740 83240 760
rect 82392 692 82400 726
rect 82390 680 82400 692
rect 82320 660 82400 680
rect 82430 682 82630 688
rect 82430 648 82442 682
rect 82618 680 82630 682
rect 82928 682 83128 688
rect 82928 680 82940 682
rect 82618 670 82940 680
rect 82618 650 82750 670
rect 82618 648 82630 650
rect 82430 642 82630 648
rect 82740 610 82750 650
rect 82810 650 82940 670
rect 82810 610 82820 650
rect 82928 648 82940 650
rect 83116 648 83128 682
rect 83160 680 83170 740
rect 83230 680 83240 740
rect 83160 660 83240 680
rect 82928 642 83128 648
rect 82740 600 82820 610
rect 82210 150 82280 580
rect 83290 580 83300 820
rect 83340 580 83360 820
rect 83290 170 83360 580
rect 82210 140 82290 150
rect 83390 140 83420 29070
rect 83480 140 83510 29070
rect 83540 140 83570 29070
rect 83660 140 83690 29070
rect 83780 140 83810 29070
rect 83900 140 83930 29070
rect 84020 140 84050 29070
rect 84140 140 84170 29070
rect 84260 140 84290 29070
rect 82210 80 82220 140
rect 82280 80 82290 140
rect 82210 70 82290 80
rect 83270 130 83360 140
rect 83270 70 83280 130
rect 83350 70 83360 130
rect 82210 -110 82280 70
rect 83270 60 83360 70
rect 83290 0 83360 60
rect 83280 -10 83360 0
rect 83280 -70 83290 -10
rect 83350 -70 83360 -10
rect 83280 -80 83360 -70
rect 82210 -120 83360 -110
rect 82210 -180 82220 -120
rect 82280 -170 83360 -120
rect 82280 -180 82290 -170
rect 82210 -190 82290 -180
rect 82210 -570 82280 -190
rect 82210 -810 82230 -570
rect 82270 -810 82280 -570
rect 83290 -570 83360 -170
rect 82740 -590 82820 -580
rect 82430 -630 82630 -624
rect 82740 -630 82750 -590
rect 82320 -660 82400 -640
rect 82320 -720 82330 -660
rect 82390 -674 82400 -660
rect 82430 -664 82442 -630
rect 82618 -650 82750 -630
rect 82810 -630 82820 -590
rect 82928 -630 83128 -624
rect 82810 -650 82940 -630
rect 82618 -660 82940 -650
rect 82618 -664 82630 -660
rect 82430 -670 82630 -664
rect 82928 -664 82940 -660
rect 83116 -664 83128 -630
rect 82928 -670 83128 -664
rect 83160 -660 83240 -640
rect 82392 -708 82400 -674
rect 82390 -720 82400 -708
rect 82320 -740 82400 -720
rect 82430 -718 82630 -712
rect 82430 -752 82442 -718
rect 82618 -720 82630 -718
rect 82928 -718 83128 -712
rect 82928 -720 82940 -718
rect 82618 -750 82940 -720
rect 82618 -752 82630 -750
rect 82430 -758 82630 -752
rect 82210 -870 82280 -810
rect 82210 -1130 82230 -870
rect 82270 -1130 82280 -870
rect 82740 -760 82820 -750
rect 82928 -752 82940 -750
rect 83116 -752 83128 -718
rect 83160 -720 83170 -660
rect 83230 -720 83240 -660
rect 83160 -740 83240 -720
rect 82928 -758 83128 -752
rect 82740 -820 82750 -760
rect 82810 -820 82820 -760
rect 82740 -870 82820 -820
rect 82740 -930 82750 -870
rect 82810 -930 82820 -870
rect 82430 -940 82630 -934
rect 82740 -940 82820 -930
rect 83290 -810 83300 -570
rect 83340 -810 83360 -570
rect 83290 -890 83360 -810
rect 82928 -940 83128 -934
rect 82320 -970 82400 -950
rect 82320 -1030 82330 -970
rect 82390 -984 82400 -970
rect 82430 -974 82442 -940
rect 82618 -970 82940 -940
rect 82618 -974 82630 -970
rect 82430 -980 82630 -974
rect 82928 -974 82940 -970
rect 83116 -974 83128 -940
rect 82928 -980 83128 -974
rect 83160 -970 83240 -950
rect 82392 -1018 82400 -984
rect 82390 -1030 82400 -1018
rect 82320 -1050 82400 -1030
rect 82430 -1028 82630 -1022
rect 82430 -1062 82442 -1028
rect 82618 -1030 82630 -1028
rect 82928 -1028 83128 -1022
rect 82928 -1030 82940 -1028
rect 82618 -1040 82940 -1030
rect 82618 -1060 82750 -1040
rect 82618 -1062 82630 -1060
rect 82430 -1068 82630 -1062
rect 82740 -1100 82750 -1060
rect 82810 -1060 82940 -1040
rect 82810 -1100 82820 -1060
rect 82928 -1062 82940 -1060
rect 83116 -1062 83128 -1028
rect 83160 -1030 83170 -970
rect 83230 -1030 83240 -970
rect 83160 -1050 83240 -1030
rect 82928 -1068 83128 -1062
rect 82740 -1110 82820 -1100
rect 82210 -1710 82280 -1130
rect 83290 -1130 83300 -890
rect 83340 -1130 83360 -890
rect 83290 -1540 83360 -1130
rect 83270 -1580 83360 -1570
rect 83270 -1640 83280 -1580
rect 83350 -1640 83360 -1580
rect 83270 -1650 83360 -1640
rect 83290 -1710 83360 -1650
rect 83390 -1710 83420 -110
rect 83480 -1710 83510 -110
rect 83540 -1710 83570 -110
rect 83660 -1710 83690 -110
rect 83780 -1710 83810 -110
rect 83900 -1710 83930 -110
rect 84020 -1710 84050 -110
rect 84140 -1710 84170 -110
rect 84260 -1710 84290 -110
<< via1 >>
rect 4160 32590 4220 32650
rect 9150 32590 9210 32650
rect 14140 32590 14200 32650
rect 19130 32590 19190 32650
rect 24120 32590 24180 32650
rect 29110 32590 29170 32650
rect 34100 32590 34160 32650
rect 39090 32590 39150 32650
rect 44080 32590 44140 32650
rect 49070 32590 49130 32650
rect 54060 32590 54120 32650
rect 59050 32590 59110 32650
rect 64040 32590 64100 32650
rect 69030 32590 69090 32650
rect 74020 32590 74080 32650
rect 79010 32590 79070 32650
rect 4100 32450 4160 32510
rect 9090 32450 9150 32510
rect 14080 32450 14140 32510
rect 19070 32450 19130 32510
rect 24060 32450 24120 32510
rect 29050 32450 29110 32510
rect 34040 32450 34100 32510
rect 39030 32450 39090 32510
rect 44020 32450 44080 32510
rect 49010 32450 49070 32510
rect 54000 32450 54060 32510
rect 58990 32450 59050 32510
rect 63980 32450 64040 32510
rect 68970 32450 69030 32510
rect 73960 32450 74020 32510
rect 78950 32450 79010 32510
rect 14320 32310 14380 32370
rect 19310 32310 19370 32370
rect 24300 32310 24360 32370
rect 29290 32310 29350 32370
rect 34280 32310 34340 32370
rect 39270 32310 39330 32370
rect 44260 32310 44320 32370
rect 49250 32310 49310 32370
rect 54240 32310 54300 32370
rect 59230 32310 59290 32370
rect 64220 32310 64280 32370
rect 69210 32310 69270 32370
rect 14260 32170 14320 32230
rect 19250 32170 19310 32230
rect 24240 32170 24300 32230
rect 29230 32170 29290 32230
rect 34220 32170 34280 32230
rect 39210 32170 39270 32230
rect 44200 32170 44260 32230
rect 49190 32170 49250 32230
rect 54180 32170 54240 32230
rect 59170 32170 59230 32230
rect 64160 32170 64220 32230
rect 69150 32170 69210 32230
rect 24660 32030 24720 32090
rect 29650 32030 29710 32090
rect 34460 32030 34520 32090
rect 39450 32030 39510 32090
rect 44440 32030 44500 32090
rect 49430 32030 49490 32090
rect 54600 32030 54660 32090
rect 59590 32030 59650 32090
rect 24600 31890 24660 31950
rect 29590 31890 29650 31950
rect 34400 31890 34460 31950
rect 39390 31890 39450 31950
rect 44380 31890 44440 31950
rect 49370 31890 49430 31950
rect 54540 31890 54600 31950
rect 59530 31890 59590 31950
rect 24480 31750 24540 31810
rect 29470 31750 29530 31810
rect 34640 31750 34700 31810
rect 39630 31750 39690 31810
rect 44620 31750 44680 31810
rect 49610 31750 49670 31810
rect 54420 31750 54480 31810
rect 59410 31750 59470 31810
rect 24420 31610 24480 31670
rect 29410 31610 29470 31670
rect 34580 31610 34640 31670
rect 39570 31610 39630 31670
rect 44560 31610 44620 31670
rect 49550 31610 49610 31670
rect 54360 31610 54420 31670
rect 59350 31610 59410 31670
rect 35000 31470 35060 31530
rect 39810 31470 39870 31530
rect 44800 31470 44860 31530
rect 49970 31470 50030 31530
rect 34940 31330 35000 31390
rect 39750 31330 39810 31390
rect 44740 31330 44800 31390
rect 49910 31330 49970 31390
rect 34820 31190 34880 31250
rect 49790 31190 49850 31250
rect 34760 31050 34820 31110
rect 49730 31050 49790 31110
rect 39990 30910 40050 30970
rect 45160 30910 45220 30970
rect 39930 30770 39990 30830
rect 45100 30770 45160 30830
rect 45010 30630 45070 30690
rect 44920 30490 44980 30550
rect 40170 30350 40230 30410
rect 40100 30210 40160 30270
rect -5100 30120 -5040 30180
rect -5510 30060 -5450 30120
rect 3870 30060 3930 30120
rect 8860 30060 8920 30120
rect 13850 30060 13910 30120
rect 18840 30060 18900 30120
rect 23830 30060 23890 30120
rect 28820 30060 28880 30120
rect 33810 30060 33870 30120
rect 38800 30060 38860 30120
rect 43790 30060 43850 30120
rect 48780 30060 48840 30120
rect 53770 30060 53830 30120
rect 58760 30060 58820 30120
rect 63750 30060 63810 30120
rect 68740 30060 68800 30120
rect 73730 30060 73790 30120
rect 78720 30060 78780 30120
rect -5240 29930 -5180 29990
rect -5360 29790 -5300 29850
rect 2350 29530 2410 29590
rect -2070 29080 -2010 29140
rect 2650 29080 2710 29140
rect 3720 29080 3780 29140
rect 2650 28890 2710 28950
rect 2760 28396 2820 28410
rect 3180 28420 3240 28480
rect 2760 28362 2788 28396
rect 2788 28362 2820 28396
rect 2760 28350 2820 28362
rect 3600 28396 3660 28410
rect 3600 28362 3605 28396
rect 3605 28362 3639 28396
rect 3639 28362 3660 28396
rect 3600 28350 3660 28362
rect 3180 28250 3240 28310
rect 3180 28140 3240 28200
rect 2760 28086 2820 28100
rect 2760 28052 2788 28086
rect 2788 28052 2820 28086
rect 2760 28040 2820 28052
rect 3180 27970 3240 28030
rect 3600 28086 3660 28100
rect 3600 28052 3605 28086
rect 3605 28052 3639 28086
rect 3639 28052 3660 28086
rect 3600 28040 3660 28052
rect 4170 29530 4230 29590
rect 7340 29530 7400 29590
rect 3880 29080 3940 29140
rect 7640 29080 7700 29140
rect 8710 29080 8770 29140
rect 7640 28890 7700 28950
rect 7750 28396 7810 28410
rect 8170 28420 8230 28480
rect 7750 28362 7778 28396
rect 7778 28362 7810 28396
rect 7750 28350 7810 28362
rect 8590 28396 8650 28410
rect 8590 28362 8595 28396
rect 8595 28362 8629 28396
rect 8629 28362 8650 28396
rect 8590 28350 8650 28362
rect 8170 28250 8230 28310
rect 8170 28140 8230 28200
rect 7750 28086 7810 28100
rect 7750 28052 7778 28086
rect 7778 28052 7810 28086
rect 7750 28040 7810 28052
rect 8170 27970 8230 28030
rect 8590 28086 8650 28100
rect 8590 28052 8595 28086
rect 8595 28052 8629 28086
rect 8629 28052 8650 28086
rect 8590 28040 8650 28052
rect 9160 29530 9220 29590
rect 8870 29080 8930 29140
rect 12150 29470 12210 29530
rect 12330 29530 12390 29590
rect 12630 29080 12690 29140
rect 13700 29080 13760 29140
rect 12630 28890 12690 28950
rect 12740 28396 12800 28410
rect 13160 28420 13220 28480
rect 12740 28362 12768 28396
rect 12768 28362 12800 28396
rect 12740 28350 12800 28362
rect 13580 28396 13640 28410
rect 13580 28362 13585 28396
rect 13585 28362 13619 28396
rect 13619 28362 13640 28396
rect 13580 28350 13640 28362
rect 13160 28250 13220 28310
rect 13160 28140 13220 28200
rect 12740 28086 12800 28100
rect 12740 28052 12768 28086
rect 12768 28052 12800 28086
rect 12740 28040 12800 28052
rect 13160 27970 13220 28030
rect 13580 28086 13640 28100
rect 13580 28052 13585 28086
rect 13585 28052 13619 28086
rect 13619 28052 13640 28086
rect 13580 28040 13640 28052
rect 14150 29530 14210 29590
rect 13860 29080 13920 29140
rect 14330 29470 14390 29530
rect 17140 29470 17200 29530
rect 17320 29530 17380 29590
rect 17620 29080 17680 29140
rect 18690 29080 18750 29140
rect 17620 28890 17680 28950
rect 17730 28396 17790 28410
rect 18150 28420 18210 28480
rect 17730 28362 17758 28396
rect 17758 28362 17790 28396
rect 17730 28350 17790 28362
rect 18570 28396 18630 28410
rect 18570 28362 18575 28396
rect 18575 28362 18609 28396
rect 18609 28362 18630 28396
rect 18570 28350 18630 28362
rect 18150 28250 18210 28310
rect 18150 28140 18210 28200
rect 17730 28086 17790 28100
rect 17730 28052 17758 28086
rect 17758 28052 17790 28086
rect 17730 28040 17790 28052
rect 18150 27970 18210 28030
rect 18570 28086 18630 28100
rect 18570 28052 18575 28086
rect 18575 28052 18609 28086
rect 18609 28052 18630 28086
rect 18570 28040 18630 28052
rect 19140 29530 19200 29590
rect 18850 29080 18910 29140
rect 19320 29470 19380 29530
rect 21770 29350 21830 29410
rect 21950 29410 22010 29470
rect 22130 29470 22190 29530
rect 22310 29530 22370 29590
rect 22610 29080 22670 29140
rect 23680 29080 23740 29140
rect 22610 28890 22670 28950
rect 22720 28396 22780 28410
rect 23140 28420 23200 28480
rect 22720 28362 22748 28396
rect 22748 28362 22780 28396
rect 22720 28350 22780 28362
rect 23560 28396 23620 28410
rect 23560 28362 23565 28396
rect 23565 28362 23599 28396
rect 23599 28362 23620 28396
rect 23560 28350 23620 28362
rect 23140 28250 23200 28310
rect 23140 28140 23200 28200
rect 22720 28086 22780 28100
rect 22720 28052 22748 28086
rect 22748 28052 22780 28086
rect 22720 28040 22780 28052
rect 23140 27970 23200 28030
rect 23560 28086 23620 28100
rect 23560 28052 23565 28086
rect 23565 28052 23599 28086
rect 23599 28052 23620 28086
rect 23560 28040 23620 28052
rect 24130 29530 24190 29590
rect 23840 29080 23900 29140
rect 24310 29470 24370 29530
rect 24490 29410 24550 29470
rect 24670 29350 24730 29410
rect 26760 29350 26820 29410
rect 26940 29410 27000 29470
rect 27120 29470 27180 29530
rect 27300 29530 27360 29590
rect 27600 29080 27660 29140
rect 28670 29080 28730 29140
rect 27600 28890 27660 28950
rect 27710 28396 27770 28410
rect 28130 28420 28190 28480
rect 27710 28362 27738 28396
rect 27738 28362 27770 28396
rect 27710 28350 27770 28362
rect 28550 28396 28610 28410
rect 28550 28362 28555 28396
rect 28555 28362 28589 28396
rect 28589 28362 28610 28396
rect 28550 28350 28610 28362
rect 28130 28250 28190 28310
rect 28130 28140 28190 28200
rect 27710 28086 27770 28100
rect 27710 28052 27738 28086
rect 27738 28052 27770 28086
rect 27710 28040 27770 28052
rect 28130 27970 28190 28030
rect 28550 28086 28610 28100
rect 28550 28052 28555 28086
rect 28555 28052 28589 28086
rect 28589 28052 28610 28086
rect 28550 28040 28610 28052
rect 29120 29530 29180 29590
rect 28830 29080 28890 29140
rect 29300 29470 29360 29530
rect 29480 29410 29540 29470
rect 29660 29350 29720 29410
rect 31390 29230 31450 29290
rect 31570 29290 31630 29350
rect 31750 29350 31810 29410
rect 31930 29410 31990 29470
rect 32110 29470 32170 29530
rect 32290 29530 32350 29590
rect 32590 29080 32650 29140
rect 33660 29080 33720 29140
rect 32590 28890 32650 28950
rect 32700 28396 32760 28410
rect 33120 28420 33180 28480
rect 32700 28362 32728 28396
rect 32728 28362 32760 28396
rect 32700 28350 32760 28362
rect 33540 28396 33600 28410
rect 33540 28362 33545 28396
rect 33545 28362 33579 28396
rect 33579 28362 33600 28396
rect 33540 28350 33600 28362
rect 33120 28250 33180 28310
rect 33120 28140 33180 28200
rect 32700 28086 32760 28100
rect 32700 28052 32728 28086
rect 32728 28052 32760 28086
rect 32700 28040 32760 28052
rect 33120 27970 33180 28030
rect 33540 28086 33600 28100
rect 33540 28052 33545 28086
rect 33545 28052 33579 28086
rect 33579 28052 33600 28086
rect 33540 28040 33600 28052
rect 34110 29530 34170 29590
rect 33820 29080 33880 29140
rect 34290 29470 34350 29530
rect 34470 29410 34530 29470
rect 34650 29350 34710 29410
rect 34830 29290 34890 29350
rect 35010 29230 35070 29290
rect 36200 29170 36260 29230
rect 36380 29230 36440 29290
rect 36560 29290 36620 29350
rect 36740 29350 36800 29410
rect 36920 29410 36980 29470
rect 37100 29470 37160 29530
rect 37280 29530 37340 29590
rect 37580 29080 37640 29140
rect 38650 29080 38710 29140
rect 37580 28890 37640 28950
rect 37690 28396 37750 28410
rect 38110 28420 38170 28480
rect 37690 28362 37718 28396
rect 37718 28362 37750 28396
rect 37690 28350 37750 28362
rect 38530 28396 38590 28410
rect 38530 28362 38535 28396
rect 38535 28362 38569 28396
rect 38569 28362 38590 28396
rect 38530 28350 38590 28362
rect 38110 28250 38170 28310
rect 38110 28140 38170 28200
rect 37690 28086 37750 28100
rect 37690 28052 37718 28086
rect 37718 28052 37750 28086
rect 37690 28040 37750 28052
rect 38110 27970 38170 28030
rect 38530 28086 38590 28100
rect 38530 28052 38535 28086
rect 38535 28052 38569 28086
rect 38569 28052 38590 28086
rect 38530 28040 38590 28052
rect 39100 29530 39160 29590
rect 38810 29080 38870 29140
rect 39280 29470 39340 29530
rect 39460 29410 39520 29470
rect 39640 29350 39700 29410
rect 39820 29290 39880 29350
rect 40000 29230 40060 29290
rect 40180 29170 40240 29230
rect 41190 29170 41250 29230
rect 41370 29230 41430 29290
rect 41550 29290 41610 29350
rect 41730 29350 41790 29410
rect 41910 29410 41970 29470
rect 42090 29470 42150 29530
rect 42270 29530 42330 29590
rect 42570 29080 42630 29140
rect 43640 29080 43700 29140
rect 42570 28890 42630 28950
rect 42680 28396 42740 28410
rect 43100 28420 43160 28480
rect 42680 28362 42708 28396
rect 42708 28362 42740 28396
rect 42680 28350 42740 28362
rect 43520 28396 43580 28410
rect 43520 28362 43525 28396
rect 43525 28362 43559 28396
rect 43559 28362 43580 28396
rect 43520 28350 43580 28362
rect 43100 28250 43160 28310
rect 43100 28140 43160 28200
rect 42680 28086 42740 28100
rect 42680 28052 42708 28086
rect 42708 28052 42740 28086
rect 42680 28040 42740 28052
rect 43100 27970 43160 28030
rect 43520 28086 43580 28100
rect 43520 28052 43525 28086
rect 43525 28052 43559 28086
rect 43559 28052 43580 28086
rect 43520 28040 43580 28052
rect 44090 29530 44150 29590
rect 43800 29080 43860 29140
rect 44270 29470 44330 29530
rect 44450 29410 44510 29470
rect 44630 29350 44690 29410
rect 44810 29290 44870 29350
rect 44990 29230 45050 29290
rect 45170 29170 45230 29230
rect 46360 29230 46420 29290
rect 46540 29290 46600 29350
rect 46720 29350 46780 29410
rect 46900 29410 46960 29470
rect 47080 29470 47140 29530
rect 47260 29530 47320 29590
rect 47560 29080 47620 29140
rect 48630 29080 48690 29140
rect 47560 28890 47620 28950
rect 47670 28396 47730 28410
rect 48090 28420 48150 28480
rect 47670 28362 47698 28396
rect 47698 28362 47730 28396
rect 47670 28350 47730 28362
rect 48510 28396 48570 28410
rect 48510 28362 48515 28396
rect 48515 28362 48549 28396
rect 48549 28362 48570 28396
rect 48510 28350 48570 28362
rect 48090 28250 48150 28310
rect 48090 28140 48150 28200
rect 47670 28086 47730 28100
rect 47670 28052 47698 28086
rect 47698 28052 47730 28086
rect 47670 28040 47730 28052
rect 48090 27970 48150 28030
rect 48510 28086 48570 28100
rect 48510 28052 48515 28086
rect 48515 28052 48549 28086
rect 48549 28052 48570 28086
rect 48510 28040 48570 28052
rect 49080 29530 49140 29590
rect 48790 29080 48850 29140
rect 49260 29470 49320 29530
rect 49440 29410 49500 29470
rect 49620 29350 49680 29410
rect 49800 29290 49860 29350
rect 51710 29350 51770 29410
rect 51890 29410 51950 29470
rect 52070 29470 52130 29530
rect 52250 29530 52310 29590
rect 49980 29230 50040 29290
rect 52550 29080 52610 29140
rect 53620 29080 53680 29140
rect 52550 28890 52610 28950
rect 52660 28396 52720 28410
rect 53080 28420 53140 28480
rect 52660 28362 52688 28396
rect 52688 28362 52720 28396
rect 52660 28350 52720 28362
rect 53500 28396 53560 28410
rect 53500 28362 53505 28396
rect 53505 28362 53539 28396
rect 53539 28362 53560 28396
rect 53500 28350 53560 28362
rect 53080 28250 53140 28310
rect 53080 28140 53140 28200
rect 52660 28086 52720 28100
rect 52660 28052 52688 28086
rect 52688 28052 52720 28086
rect 52660 28040 52720 28052
rect 53080 27970 53140 28030
rect 53500 28086 53560 28100
rect 53500 28052 53505 28086
rect 53505 28052 53539 28086
rect 53539 28052 53560 28086
rect 53500 28040 53560 28052
rect 54070 29530 54130 29590
rect 53780 29080 53840 29140
rect 54250 29470 54310 29530
rect 54430 29410 54490 29470
rect 54610 29350 54670 29410
rect 56700 29350 56760 29410
rect 56880 29410 56940 29470
rect 57060 29470 57120 29530
rect 57240 29530 57300 29590
rect 57540 29080 57600 29140
rect 58610 29080 58670 29140
rect 57540 28890 57600 28950
rect 57650 28396 57710 28410
rect 58070 28420 58130 28480
rect 57650 28362 57678 28396
rect 57678 28362 57710 28396
rect 57650 28350 57710 28362
rect 58490 28396 58550 28410
rect 58490 28362 58495 28396
rect 58495 28362 58529 28396
rect 58529 28362 58550 28396
rect 58490 28350 58550 28362
rect 58070 28250 58130 28310
rect 58070 28140 58130 28200
rect 57650 28086 57710 28100
rect 57650 28052 57678 28086
rect 57678 28052 57710 28086
rect 57650 28040 57710 28052
rect 58070 27970 58130 28030
rect 58490 28086 58550 28100
rect 58490 28052 58495 28086
rect 58495 28052 58529 28086
rect 58529 28052 58550 28086
rect 58490 28040 58550 28052
rect 59060 29530 59120 29590
rect 58770 29080 58830 29140
rect 59240 29470 59300 29530
rect 59420 29410 59480 29470
rect 62050 29470 62110 29530
rect 62230 29530 62290 29590
rect 59600 29350 59660 29410
rect 62530 29080 62590 29140
rect 63600 29080 63660 29140
rect 62530 28890 62590 28950
rect 62640 28396 62700 28410
rect 63060 28420 63120 28480
rect 62640 28362 62668 28396
rect 62668 28362 62700 28396
rect 62640 28350 62700 28362
rect 63480 28396 63540 28410
rect 63480 28362 63485 28396
rect 63485 28362 63519 28396
rect 63519 28362 63540 28396
rect 63480 28350 63540 28362
rect 63060 28250 63120 28310
rect 63060 28140 63120 28200
rect 62640 28086 62700 28100
rect 62640 28052 62668 28086
rect 62668 28052 62700 28086
rect 62640 28040 62700 28052
rect 63060 27970 63120 28030
rect 63480 28086 63540 28100
rect 63480 28052 63485 28086
rect 63485 28052 63519 28086
rect 63519 28052 63540 28086
rect 63480 28040 63540 28052
rect 64050 29530 64110 29590
rect 63760 29080 63820 29140
rect 64230 29470 64290 29530
rect 67040 29470 67100 29530
rect 67220 29530 67280 29590
rect 67520 29080 67580 29140
rect 68590 29080 68650 29140
rect 67520 28890 67580 28950
rect 67630 28396 67690 28410
rect 68050 28420 68110 28480
rect 67630 28362 67658 28396
rect 67658 28362 67690 28396
rect 67630 28350 67690 28362
rect 68470 28396 68530 28410
rect 68470 28362 68475 28396
rect 68475 28362 68509 28396
rect 68509 28362 68530 28396
rect 68470 28350 68530 28362
rect 68050 28250 68110 28310
rect 68050 28140 68110 28200
rect 67630 28086 67690 28100
rect 67630 28052 67658 28086
rect 67658 28052 67690 28086
rect 67630 28040 67690 28052
rect 68050 27970 68110 28030
rect 68470 28086 68530 28100
rect 68470 28052 68475 28086
rect 68475 28052 68509 28086
rect 68509 28052 68530 28086
rect 68470 28040 68530 28052
rect 69040 29530 69100 29590
rect 68750 29080 68810 29140
rect 69220 29470 69280 29530
rect 72210 29530 72270 29590
rect 72510 29080 72570 29140
rect 73580 29080 73640 29140
rect 72510 28890 72570 28950
rect 72620 28396 72680 28410
rect 73040 28420 73100 28480
rect 72620 28362 72648 28396
rect 72648 28362 72680 28396
rect 72620 28350 72680 28362
rect 73460 28396 73520 28410
rect 73460 28362 73465 28396
rect 73465 28362 73499 28396
rect 73499 28362 73520 28396
rect 73460 28350 73520 28362
rect 73040 28250 73100 28310
rect 73040 28140 73100 28200
rect 72620 28086 72680 28100
rect 72620 28052 72648 28086
rect 72648 28052 72680 28086
rect 72620 28040 72680 28052
rect 73040 27970 73100 28030
rect 73460 28086 73520 28100
rect 73460 28052 73465 28086
rect 73465 28052 73499 28086
rect 73499 28052 73520 28086
rect 73460 28040 73520 28052
rect 74030 29530 74090 29590
rect 77200 29530 77260 29590
rect 73740 29080 73800 29140
rect 77500 29080 77560 29140
rect 78570 29080 78630 29140
rect 77500 28890 77560 28950
rect 77610 28396 77670 28410
rect 78030 28420 78090 28480
rect 77610 28362 77638 28396
rect 77638 28362 77670 28396
rect 77610 28350 77670 28362
rect 78450 28396 78510 28410
rect 78450 28362 78455 28396
rect 78455 28362 78489 28396
rect 78489 28362 78510 28396
rect 78450 28350 78510 28362
rect 78030 28250 78090 28310
rect 78030 28140 78090 28200
rect 77610 28086 77670 28100
rect 77610 28052 77638 28086
rect 77638 28052 77670 28086
rect 77610 28040 77670 28052
rect 78030 27970 78090 28030
rect 78450 28086 78510 28100
rect 78450 28052 78455 28086
rect 78455 28052 78489 28086
rect 78489 28052 78510 28086
rect 78450 28040 78510 28052
rect 79020 29530 79080 29590
rect 78730 29080 78790 29140
rect 82220 29080 82280 29140
rect -1000 23870 -940 23930
rect -2070 23760 -2010 23820
rect -1960 23266 -1900 23280
rect -1540 23290 -1480 23350
rect -1960 23232 -1932 23266
rect -1932 23232 -1900 23266
rect -1960 23220 -1900 23232
rect -1120 23266 -1060 23280
rect -1120 23232 -1115 23266
rect -1115 23232 -1081 23266
rect -1081 23232 -1060 23266
rect -1120 23220 -1060 23232
rect -1540 23120 -1480 23180
rect -1540 23010 -1480 23070
rect -1960 22956 -1900 22970
rect -1960 22922 -1932 22956
rect -1932 22922 -1900 22956
rect -1960 22910 -1900 22922
rect -1540 22840 -1480 22900
rect -1120 22956 -1060 22970
rect -1120 22922 -1115 22956
rect -1115 22922 -1081 22956
rect -1081 22922 -1060 22956
rect -1120 22910 -1060 22922
rect -1010 22300 -940 22360
rect -1000 22160 -940 22220
rect -2070 22050 -2010 22110
rect -1960 21556 -1900 21570
rect -1540 21580 -1480 21640
rect -1960 21522 -1932 21556
rect -1932 21522 -1900 21556
rect -1960 21510 -1900 21522
rect -1120 21556 -1060 21570
rect -1120 21522 -1115 21556
rect -1115 21522 -1081 21556
rect -1081 21522 -1060 21556
rect -1120 21510 -1060 21522
rect -1540 21410 -1480 21470
rect -1540 21300 -1480 21360
rect -1960 21246 -1900 21260
rect -1960 21212 -1932 21246
rect -1932 21212 -1900 21246
rect -1960 21200 -1900 21212
rect -1540 21130 -1480 21190
rect -1120 21246 -1060 21260
rect -1120 21212 -1115 21246
rect -1115 21212 -1081 21246
rect -1081 21212 -1060 21246
rect -1120 21200 -1060 21212
rect -1010 20590 -940 20650
rect -1000 20450 -940 20510
rect -2070 20340 -2010 20400
rect -1960 19846 -1900 19860
rect -1540 19870 -1480 19930
rect -1960 19812 -1932 19846
rect -1932 19812 -1900 19846
rect -1960 19800 -1900 19812
rect -1120 19846 -1060 19860
rect -1120 19812 -1115 19846
rect -1115 19812 -1081 19846
rect -1081 19812 -1060 19846
rect -1120 19800 -1060 19812
rect -1540 19700 -1480 19760
rect -1540 19590 -1480 19650
rect -1960 19536 -1900 19550
rect -1960 19502 -1932 19536
rect -1932 19502 -1900 19536
rect -1960 19490 -1900 19502
rect -1540 19420 -1480 19480
rect -1120 19536 -1060 19550
rect -1120 19502 -1115 19536
rect -1115 19502 -1081 19536
rect -1081 19502 -1060 19536
rect -1120 19490 -1060 19502
rect -1010 18880 -940 18940
rect -1000 18740 -940 18800
rect -2070 18630 -2010 18690
rect -1960 18136 -1900 18150
rect -1540 18160 -1480 18220
rect -1960 18102 -1932 18136
rect -1932 18102 -1900 18136
rect -1960 18090 -1900 18102
rect -1120 18136 -1060 18150
rect -1120 18102 -1115 18136
rect -1115 18102 -1081 18136
rect -1081 18102 -1060 18136
rect -1120 18090 -1060 18102
rect -1540 17990 -1480 18050
rect -1540 17880 -1480 17940
rect -1960 17826 -1900 17840
rect -1960 17792 -1932 17826
rect -1932 17792 -1900 17826
rect -1960 17780 -1900 17792
rect -1540 17710 -1480 17770
rect -1120 17826 -1060 17840
rect -1120 17792 -1115 17826
rect -1115 17792 -1081 17826
rect -1081 17792 -1060 17826
rect -1120 17780 -1060 17792
rect -1010 17170 -940 17230
rect -1000 17030 -940 17090
rect -2070 16920 -2010 16980
rect -1960 16426 -1900 16440
rect -1540 16450 -1480 16510
rect -1960 16392 -1932 16426
rect -1932 16392 -1900 16426
rect -1960 16380 -1900 16392
rect -1120 16426 -1060 16440
rect -1120 16392 -1115 16426
rect -1115 16392 -1081 16426
rect -1081 16392 -1060 16426
rect -1120 16380 -1060 16392
rect -1540 16280 -1480 16340
rect -1540 16170 -1480 16230
rect -1960 16116 -1900 16130
rect -1960 16082 -1932 16116
rect -1932 16082 -1900 16116
rect -1960 16070 -1900 16082
rect -1540 16000 -1480 16060
rect -1120 16116 -1060 16130
rect -1120 16082 -1115 16116
rect -1115 16082 -1081 16116
rect -1081 16082 -1060 16116
rect -1120 16070 -1060 16082
rect -1010 15460 -940 15520
rect -1000 15320 -940 15380
rect -2070 15210 -2010 15270
rect -1960 14716 -1900 14730
rect -1540 14740 -1480 14800
rect -1960 14682 -1932 14716
rect -1932 14682 -1900 14716
rect -1960 14670 -1900 14682
rect -1120 14716 -1060 14730
rect -1120 14682 -1115 14716
rect -1115 14682 -1081 14716
rect -1081 14682 -1060 14716
rect -1120 14670 -1060 14682
rect -1540 14570 -1480 14630
rect -1540 14460 -1480 14520
rect -1960 14406 -1900 14420
rect -1960 14372 -1932 14406
rect -1932 14372 -1900 14406
rect -1960 14360 -1900 14372
rect -1540 14290 -1480 14350
rect -1120 14406 -1060 14420
rect -1120 14372 -1115 14406
rect -1115 14372 -1081 14406
rect -1081 14372 -1060 14406
rect -1120 14360 -1060 14372
rect -1010 13750 -940 13810
rect -1000 13610 -940 13670
rect -2070 13500 -2010 13560
rect -1960 13006 -1900 13020
rect -1540 13030 -1480 13090
rect -1960 12972 -1932 13006
rect -1932 12972 -1900 13006
rect -1960 12960 -1900 12972
rect -1120 13006 -1060 13020
rect -1120 12972 -1115 13006
rect -1115 12972 -1081 13006
rect -1081 12972 -1060 13006
rect -1120 12960 -1060 12972
rect -1540 12860 -1480 12920
rect -1540 12750 -1480 12810
rect -1960 12696 -1900 12710
rect -1960 12662 -1932 12696
rect -1932 12662 -1900 12696
rect -1960 12650 -1900 12662
rect -1540 12580 -1480 12640
rect -1120 12696 -1060 12710
rect -1120 12662 -1115 12696
rect -1115 12662 -1081 12696
rect -1081 12662 -1060 12696
rect -1120 12650 -1060 12662
rect -1010 12040 -940 12100
rect -1000 11900 -940 11960
rect -2070 11790 -2010 11850
rect -1960 11296 -1900 11310
rect -1540 11320 -1480 11380
rect -1960 11262 -1932 11296
rect -1932 11262 -1900 11296
rect -1960 11250 -1900 11262
rect -1120 11296 -1060 11310
rect -1120 11262 -1115 11296
rect -1115 11262 -1081 11296
rect -1081 11262 -1060 11296
rect -1120 11250 -1060 11262
rect -1540 11150 -1480 11210
rect -1540 11040 -1480 11100
rect -1960 10986 -1900 11000
rect -1960 10952 -1932 10986
rect -1932 10952 -1900 10986
rect -1960 10940 -1900 10952
rect -1540 10870 -1480 10930
rect -1120 10986 -1060 11000
rect -1120 10952 -1115 10986
rect -1115 10952 -1081 10986
rect -1081 10952 -1060 10986
rect -1120 10940 -1060 10952
rect -1010 10330 -940 10390
rect -1000 10190 -940 10250
rect -2070 10080 -2010 10140
rect -1960 9586 -1900 9600
rect -1540 9610 -1480 9670
rect -1960 9552 -1932 9586
rect -1932 9552 -1900 9586
rect -1960 9540 -1900 9552
rect -1120 9586 -1060 9600
rect -1120 9552 -1115 9586
rect -1115 9552 -1081 9586
rect -1081 9552 -1060 9586
rect -1120 9540 -1060 9552
rect -1540 9440 -1480 9500
rect -1540 9330 -1480 9390
rect -1960 9276 -1900 9290
rect -1960 9242 -1932 9276
rect -1932 9242 -1900 9276
rect -1960 9230 -1900 9242
rect -1540 9160 -1480 9220
rect -1120 9276 -1060 9290
rect -1120 9242 -1115 9276
rect -1115 9242 -1081 9276
rect -1081 9242 -1060 9276
rect -1120 9230 -1060 9242
rect -1010 8620 -940 8680
rect -1000 8480 -940 8540
rect -2070 8370 -2010 8430
rect -1960 7876 -1900 7890
rect -1540 7900 -1480 7960
rect -1960 7842 -1932 7876
rect -1932 7842 -1900 7876
rect -1960 7830 -1900 7842
rect -1120 7876 -1060 7890
rect -1120 7842 -1115 7876
rect -1115 7842 -1081 7876
rect -1081 7842 -1060 7876
rect -1120 7830 -1060 7842
rect -1540 7730 -1480 7790
rect -1540 7620 -1480 7680
rect -1960 7566 -1900 7580
rect -1960 7532 -1932 7566
rect -1932 7532 -1900 7566
rect -1960 7520 -1900 7532
rect -1540 7450 -1480 7510
rect -1120 7566 -1060 7580
rect -1120 7532 -1115 7566
rect -1115 7532 -1081 7566
rect -1081 7532 -1060 7566
rect -1120 7520 -1060 7532
rect -1010 6910 -940 6970
rect -1000 6770 -940 6830
rect -2070 6660 -2010 6720
rect -1960 6166 -1900 6180
rect -1540 6190 -1480 6250
rect -1960 6132 -1932 6166
rect -1932 6132 -1900 6166
rect -1960 6120 -1900 6132
rect -1120 6166 -1060 6180
rect -1120 6132 -1115 6166
rect -1115 6132 -1081 6166
rect -1081 6132 -1060 6166
rect -1120 6120 -1060 6132
rect -1540 6020 -1480 6080
rect -1540 5910 -1480 5970
rect -1960 5856 -1900 5870
rect -1960 5822 -1932 5856
rect -1932 5822 -1900 5856
rect -1960 5810 -1900 5822
rect -1540 5740 -1480 5800
rect -1120 5856 -1060 5870
rect -1120 5822 -1115 5856
rect -1115 5822 -1081 5856
rect -1081 5822 -1060 5856
rect -1120 5810 -1060 5822
rect -1010 5200 -940 5260
rect -1000 5060 -940 5120
rect -2070 4950 -2010 5010
rect -1960 4456 -1900 4470
rect -1540 4480 -1480 4540
rect -1960 4422 -1932 4456
rect -1932 4422 -1900 4456
rect -1960 4410 -1900 4422
rect -1120 4456 -1060 4470
rect -1120 4422 -1115 4456
rect -1115 4422 -1081 4456
rect -1081 4422 -1060 4456
rect -1120 4410 -1060 4422
rect -1540 4310 -1480 4370
rect -1540 4200 -1480 4260
rect -1960 4146 -1900 4160
rect -1960 4112 -1932 4146
rect -1932 4112 -1900 4146
rect -1960 4100 -1900 4112
rect -1540 4030 -1480 4090
rect -1120 4146 -1060 4160
rect -1120 4112 -1115 4146
rect -1115 4112 -1081 4146
rect -1081 4112 -1060 4146
rect -1120 4100 -1060 4112
rect -1010 3490 -940 3550
rect -1000 3350 -940 3410
rect -2070 3240 -2010 3300
rect -1960 2746 -1900 2760
rect -1540 2770 -1480 2830
rect -1960 2712 -1932 2746
rect -1932 2712 -1900 2746
rect -1960 2700 -1900 2712
rect -1120 2746 -1060 2760
rect -1120 2712 -1115 2746
rect -1115 2712 -1081 2746
rect -1081 2712 -1060 2746
rect -1120 2700 -1060 2712
rect -1540 2600 -1480 2660
rect -1540 2490 -1480 2550
rect -1960 2436 -1900 2450
rect -1960 2402 -1932 2436
rect -1932 2402 -1900 2436
rect -1960 2390 -1900 2402
rect -1540 2320 -1480 2380
rect -1120 2436 -1060 2450
rect -1120 2402 -1115 2436
rect -1115 2402 -1081 2436
rect -1081 2402 -1060 2436
rect -1120 2390 -1060 2402
rect -1010 1780 -940 1840
rect -1000 1640 -940 1700
rect -2070 1530 -2010 1590
rect -1960 1036 -1900 1050
rect -1540 1060 -1480 1120
rect -1960 1002 -1932 1036
rect -1932 1002 -1900 1036
rect -1960 990 -1900 1002
rect -1120 1036 -1060 1050
rect -1120 1002 -1115 1036
rect -1115 1002 -1081 1036
rect -1081 1002 -1060 1036
rect -1120 990 -1060 1002
rect -1540 890 -1480 950
rect -1540 780 -1480 840
rect -1960 726 -1900 740
rect -1960 692 -1932 726
rect -1932 692 -1900 726
rect -1960 680 -1900 692
rect -1540 610 -1480 670
rect -1120 726 -1060 740
rect -1120 692 -1115 726
rect -1115 692 -1081 726
rect -1081 692 -1060 726
rect -1120 680 -1060 692
rect -2070 80 -2010 140
rect -1010 70 -940 130
rect -1000 -70 -940 -10
rect -2070 -180 -2010 -120
rect -1960 -674 -1900 -660
rect -1540 -650 -1480 -590
rect -1960 -708 -1932 -674
rect -1932 -708 -1900 -674
rect -1960 -720 -1900 -708
rect -1120 -674 -1060 -660
rect -1120 -708 -1115 -674
rect -1115 -708 -1081 -674
rect -1081 -708 -1060 -674
rect -1120 -720 -1060 -708
rect -1540 -820 -1480 -760
rect -1540 -930 -1480 -870
rect -1960 -984 -1900 -970
rect -1960 -1018 -1932 -984
rect -1932 -1018 -1900 -984
rect -1960 -1030 -1900 -1018
rect -1540 -1100 -1480 -1040
rect -1120 -984 -1060 -970
rect -1120 -1018 -1115 -984
rect -1115 -1018 -1081 -984
rect -1081 -1018 -1060 -984
rect -1120 -1030 -1060 -1018
rect -1010 -1640 -940 -1580
rect 2650 80 2710 140
rect 2650 -180 2710 -120
rect 2760 -674 2820 -660
rect 3180 -650 3240 -590
rect 2760 -708 2788 -674
rect 2788 -708 2820 -674
rect 2760 -720 2820 -708
rect 3600 -674 3660 -660
rect 3600 -708 3605 -674
rect 3605 -708 3639 -674
rect 3639 -708 3660 -674
rect 3600 -720 3660 -708
rect 3180 -820 3240 -760
rect 3180 -930 3240 -870
rect 2760 -984 2820 -970
rect 2760 -1018 2788 -984
rect 2788 -1018 2820 -984
rect 2760 -1030 2820 -1018
rect 3180 -1100 3240 -1040
rect 3600 -984 3660 -970
rect 3600 -1018 3605 -984
rect 3605 -1018 3639 -984
rect 3639 -1018 3660 -984
rect 3600 -1030 3660 -1018
rect 3720 -1700 3780 -1640
rect 7640 80 7700 140
rect 7640 -180 7700 -120
rect 7750 -674 7810 -660
rect 8170 -650 8230 -590
rect 7750 -708 7778 -674
rect 7778 -708 7810 -674
rect 7750 -720 7810 -708
rect 8590 -674 8650 -660
rect 8590 -708 8595 -674
rect 8595 -708 8629 -674
rect 8629 -708 8650 -674
rect 8590 -720 8650 -708
rect 8170 -820 8230 -760
rect 8170 -930 8230 -870
rect 7750 -984 7810 -970
rect 7750 -1018 7778 -984
rect 7778 -1018 7810 -984
rect 7750 -1030 7810 -1018
rect 8170 -1100 8230 -1040
rect 8590 -984 8650 -970
rect 8590 -1018 8595 -984
rect 8595 -1018 8629 -984
rect 8629 -1018 8650 -984
rect 8590 -1030 8650 -1018
rect 8710 -1700 8770 -1640
rect 12630 80 12690 140
rect 12630 -180 12690 -120
rect 12740 -674 12800 -660
rect 13160 -650 13220 -590
rect 12740 -708 12768 -674
rect 12768 -708 12800 -674
rect 12740 -720 12800 -708
rect 13580 -674 13640 -660
rect 13580 -708 13585 -674
rect 13585 -708 13619 -674
rect 13619 -708 13640 -674
rect 13580 -720 13640 -708
rect 13160 -820 13220 -760
rect 13160 -930 13220 -870
rect 12740 -984 12800 -970
rect 12740 -1018 12768 -984
rect 12768 -1018 12800 -984
rect 12740 -1030 12800 -1018
rect 13160 -1100 13220 -1040
rect 13580 -984 13640 -970
rect 13580 -1018 13585 -984
rect 13585 -1018 13619 -984
rect 13619 -1018 13640 -984
rect 13580 -1030 13640 -1018
rect 13700 -1700 13760 -1640
rect 17620 80 17680 140
rect 17620 -180 17680 -120
rect 17730 -674 17790 -660
rect 18150 -650 18210 -590
rect 17730 -708 17758 -674
rect 17758 -708 17790 -674
rect 17730 -720 17790 -708
rect 18570 -674 18630 -660
rect 18570 -708 18575 -674
rect 18575 -708 18609 -674
rect 18609 -708 18630 -674
rect 18570 -720 18630 -708
rect 18150 -820 18210 -760
rect 18150 -930 18210 -870
rect 17730 -984 17790 -970
rect 17730 -1018 17758 -984
rect 17758 -1018 17790 -984
rect 17730 -1030 17790 -1018
rect 18150 -1100 18210 -1040
rect 18570 -984 18630 -970
rect 18570 -1018 18575 -984
rect 18575 -1018 18609 -984
rect 18609 -1018 18630 -984
rect 18570 -1030 18630 -1018
rect 18690 -1700 18750 -1640
rect 22610 80 22670 140
rect 22610 -180 22670 -120
rect 22720 -674 22780 -660
rect 23140 -650 23200 -590
rect 22720 -708 22748 -674
rect 22748 -708 22780 -674
rect 22720 -720 22780 -708
rect 23560 -674 23620 -660
rect 23560 -708 23565 -674
rect 23565 -708 23599 -674
rect 23599 -708 23620 -674
rect 23560 -720 23620 -708
rect 23140 -820 23200 -760
rect 23140 -930 23200 -870
rect 22720 -984 22780 -970
rect 22720 -1018 22748 -984
rect 22748 -1018 22780 -984
rect 22720 -1030 22780 -1018
rect 23140 -1100 23200 -1040
rect 23560 -984 23620 -970
rect 23560 -1018 23565 -984
rect 23565 -1018 23599 -984
rect 23599 -1018 23620 -984
rect 23560 -1030 23620 -1018
rect 23680 -1700 23740 -1640
rect 27600 80 27660 140
rect 27600 -180 27660 -120
rect 27710 -674 27770 -660
rect 28130 -650 28190 -590
rect 27710 -708 27738 -674
rect 27738 -708 27770 -674
rect 27710 -720 27770 -708
rect 28550 -674 28610 -660
rect 28550 -708 28555 -674
rect 28555 -708 28589 -674
rect 28589 -708 28610 -674
rect 28550 -720 28610 -708
rect 28130 -820 28190 -760
rect 28130 -930 28190 -870
rect 27710 -984 27770 -970
rect 27710 -1018 27738 -984
rect 27738 -1018 27770 -984
rect 27710 -1030 27770 -1018
rect 28130 -1100 28190 -1040
rect 28550 -984 28610 -970
rect 28550 -1018 28555 -984
rect 28555 -1018 28589 -984
rect 28589 -1018 28610 -984
rect 28550 -1030 28610 -1018
rect 28670 -1700 28730 -1640
rect 32590 80 32650 140
rect 32590 -180 32650 -120
rect 32700 -674 32760 -660
rect 33120 -650 33180 -590
rect 32700 -708 32728 -674
rect 32728 -708 32760 -674
rect 32700 -720 32760 -708
rect 33540 -674 33600 -660
rect 33540 -708 33545 -674
rect 33545 -708 33579 -674
rect 33579 -708 33600 -674
rect 33540 -720 33600 -708
rect 33120 -820 33180 -760
rect 33120 -930 33180 -870
rect 32700 -984 32760 -970
rect 32700 -1018 32728 -984
rect 32728 -1018 32760 -984
rect 32700 -1030 32760 -1018
rect 33120 -1100 33180 -1040
rect 33540 -984 33600 -970
rect 33540 -1018 33545 -984
rect 33545 -1018 33579 -984
rect 33579 -1018 33600 -984
rect 33540 -1030 33600 -1018
rect 33660 -1700 33720 -1640
rect 37580 80 37640 140
rect 37580 -180 37640 -120
rect 37690 -674 37750 -660
rect 38110 -650 38170 -590
rect 37690 -708 37718 -674
rect 37718 -708 37750 -674
rect 37690 -720 37750 -708
rect 38530 -674 38590 -660
rect 38530 -708 38535 -674
rect 38535 -708 38569 -674
rect 38569 -708 38590 -674
rect 38530 -720 38590 -708
rect 38110 -820 38170 -760
rect 38110 -930 38170 -870
rect 37690 -984 37750 -970
rect 37690 -1018 37718 -984
rect 37718 -1018 37750 -984
rect 37690 -1030 37750 -1018
rect 38110 -1100 38170 -1040
rect 38530 -984 38590 -970
rect 38530 -1018 38535 -984
rect 38535 -1018 38569 -984
rect 38569 -1018 38590 -984
rect 38530 -1030 38590 -1018
rect 38650 -1700 38710 -1640
rect 42570 80 42630 140
rect 42570 -180 42630 -120
rect 42680 -674 42740 -660
rect 43100 -650 43160 -590
rect 42680 -708 42708 -674
rect 42708 -708 42740 -674
rect 42680 -720 42740 -708
rect 43520 -674 43580 -660
rect 43520 -708 43525 -674
rect 43525 -708 43559 -674
rect 43559 -708 43580 -674
rect 43520 -720 43580 -708
rect 43100 -820 43160 -760
rect 43100 -930 43160 -870
rect 42680 -984 42740 -970
rect 42680 -1018 42708 -984
rect 42708 -1018 42740 -984
rect 42680 -1030 42740 -1018
rect 43100 -1100 43160 -1040
rect 43520 -984 43580 -970
rect 43520 -1018 43525 -984
rect 43525 -1018 43559 -984
rect 43559 -1018 43580 -984
rect 43520 -1030 43580 -1018
rect 43640 -1700 43700 -1640
rect 47560 80 47620 140
rect 47560 -180 47620 -120
rect 47670 -674 47730 -660
rect 48090 -650 48150 -590
rect 47670 -708 47698 -674
rect 47698 -708 47730 -674
rect 47670 -720 47730 -708
rect 48510 -674 48570 -660
rect 48510 -708 48515 -674
rect 48515 -708 48549 -674
rect 48549 -708 48570 -674
rect 48510 -720 48570 -708
rect 48090 -820 48150 -760
rect 48090 -930 48150 -870
rect 47670 -984 47730 -970
rect 47670 -1018 47698 -984
rect 47698 -1018 47730 -984
rect 47670 -1030 47730 -1018
rect 48090 -1100 48150 -1040
rect 48510 -984 48570 -970
rect 48510 -1018 48515 -984
rect 48515 -1018 48549 -984
rect 48549 -1018 48570 -984
rect 48510 -1030 48570 -1018
rect 48630 -1700 48690 -1640
rect 52550 80 52610 140
rect 52550 -180 52610 -120
rect 52660 -674 52720 -660
rect 53080 -650 53140 -590
rect 52660 -708 52688 -674
rect 52688 -708 52720 -674
rect 52660 -720 52720 -708
rect 53500 -674 53560 -660
rect 53500 -708 53505 -674
rect 53505 -708 53539 -674
rect 53539 -708 53560 -674
rect 53500 -720 53560 -708
rect 53080 -820 53140 -760
rect 53080 -930 53140 -870
rect 52660 -984 52720 -970
rect 52660 -1018 52688 -984
rect 52688 -1018 52720 -984
rect 52660 -1030 52720 -1018
rect 53080 -1100 53140 -1040
rect 53500 -984 53560 -970
rect 53500 -1018 53505 -984
rect 53505 -1018 53539 -984
rect 53539 -1018 53560 -984
rect 53500 -1030 53560 -1018
rect 53620 -1700 53680 -1640
rect 57540 80 57600 140
rect 57540 -180 57600 -120
rect 57650 -674 57710 -660
rect 58070 -650 58130 -590
rect 57650 -708 57678 -674
rect 57678 -708 57710 -674
rect 57650 -720 57710 -708
rect 58490 -674 58550 -660
rect 58490 -708 58495 -674
rect 58495 -708 58529 -674
rect 58529 -708 58550 -674
rect 58490 -720 58550 -708
rect 58070 -820 58130 -760
rect 58070 -930 58130 -870
rect 57650 -984 57710 -970
rect 57650 -1018 57678 -984
rect 57678 -1018 57710 -984
rect 57650 -1030 57710 -1018
rect 58070 -1100 58130 -1040
rect 58490 -984 58550 -970
rect 58490 -1018 58495 -984
rect 58495 -1018 58529 -984
rect 58529 -1018 58550 -984
rect 58490 -1030 58550 -1018
rect 58610 -1700 58670 -1640
rect 62530 80 62590 140
rect 62530 -180 62590 -120
rect 62640 -674 62700 -660
rect 63060 -650 63120 -590
rect 62640 -708 62668 -674
rect 62668 -708 62700 -674
rect 62640 -720 62700 -708
rect 63480 -674 63540 -660
rect 63480 -708 63485 -674
rect 63485 -708 63519 -674
rect 63519 -708 63540 -674
rect 63480 -720 63540 -708
rect 63060 -820 63120 -760
rect 63060 -930 63120 -870
rect 62640 -984 62700 -970
rect 62640 -1018 62668 -984
rect 62668 -1018 62700 -984
rect 62640 -1030 62700 -1018
rect 63060 -1100 63120 -1040
rect 63480 -984 63540 -970
rect 63480 -1018 63485 -984
rect 63485 -1018 63519 -984
rect 63519 -1018 63540 -984
rect 63480 -1030 63540 -1018
rect 63600 -1700 63660 -1640
rect 67520 80 67580 140
rect 67520 -180 67580 -120
rect 67630 -674 67690 -660
rect 68050 -650 68110 -590
rect 67630 -708 67658 -674
rect 67658 -708 67690 -674
rect 67630 -720 67690 -708
rect 68470 -674 68530 -660
rect 68470 -708 68475 -674
rect 68475 -708 68509 -674
rect 68509 -708 68530 -674
rect 68470 -720 68530 -708
rect 68050 -820 68110 -760
rect 68050 -930 68110 -870
rect 67630 -984 67690 -970
rect 67630 -1018 67658 -984
rect 67658 -1018 67690 -984
rect 67630 -1030 67690 -1018
rect 68050 -1100 68110 -1040
rect 68470 -984 68530 -970
rect 68470 -1018 68475 -984
rect 68475 -1018 68509 -984
rect 68509 -1018 68530 -984
rect 68470 -1030 68530 -1018
rect 68590 -1700 68650 -1640
rect 72510 80 72570 140
rect 72510 -180 72570 -120
rect 72620 -674 72680 -660
rect 73040 -650 73100 -590
rect 72620 -708 72648 -674
rect 72648 -708 72680 -674
rect 72620 -720 72680 -708
rect 73460 -674 73520 -660
rect 73460 -708 73465 -674
rect 73465 -708 73499 -674
rect 73499 -708 73520 -674
rect 73460 -720 73520 -708
rect 73040 -820 73100 -760
rect 73040 -930 73100 -870
rect 72620 -984 72680 -970
rect 72620 -1018 72648 -984
rect 72648 -1018 72680 -984
rect 72620 -1030 72680 -1018
rect 73040 -1100 73100 -1040
rect 73460 -984 73520 -970
rect 73460 -1018 73465 -984
rect 73465 -1018 73499 -984
rect 73499 -1018 73520 -984
rect 73460 -1030 73520 -1018
rect 73580 -1700 73640 -1640
rect 77500 80 77560 140
rect 77500 -180 77560 -120
rect 77610 -674 77670 -660
rect 78030 -650 78090 -590
rect 77610 -708 77638 -674
rect 77638 -708 77670 -674
rect 77610 -720 77670 -708
rect 78450 -674 78510 -660
rect 78450 -708 78455 -674
rect 78455 -708 78489 -674
rect 78489 -708 78510 -674
rect 78450 -720 78510 -708
rect 78030 -820 78090 -760
rect 78030 -930 78090 -870
rect 77610 -984 77670 -970
rect 77610 -1018 77638 -984
rect 77638 -1018 77670 -984
rect 77610 -1030 77670 -1018
rect 78030 -1100 78090 -1040
rect 78450 -984 78510 -970
rect 78450 -1018 78455 -984
rect 78455 -1018 78489 -984
rect 78489 -1018 78510 -984
rect 78450 -1030 78510 -1018
rect 78570 -1700 78630 -1640
rect 83290 29000 83350 29060
rect 82220 28890 82280 28950
rect 82330 28396 82390 28410
rect 82750 28420 82810 28480
rect 82330 28362 82358 28396
rect 82358 28362 82390 28396
rect 82330 28350 82390 28362
rect 83170 28396 83230 28410
rect 83170 28362 83175 28396
rect 83175 28362 83209 28396
rect 83209 28362 83230 28396
rect 83170 28350 83230 28362
rect 82750 28250 82810 28310
rect 82750 28140 82810 28200
rect 82330 28086 82390 28100
rect 82330 28052 82358 28086
rect 82358 28052 82390 28086
rect 82330 28040 82390 28052
rect 82750 27970 82810 28030
rect 83170 28086 83230 28100
rect 83170 28052 83175 28086
rect 83175 28052 83209 28086
rect 83209 28052 83230 28086
rect 83170 28040 83230 28052
rect 83280 27430 83350 27490
rect 83290 27290 83350 27350
rect 82220 27180 82280 27240
rect 82330 26686 82390 26700
rect 82750 26710 82810 26770
rect 82330 26652 82358 26686
rect 82358 26652 82390 26686
rect 82330 26640 82390 26652
rect 83170 26686 83230 26700
rect 83170 26652 83175 26686
rect 83175 26652 83209 26686
rect 83209 26652 83230 26686
rect 83170 26640 83230 26652
rect 82750 26540 82810 26600
rect 82750 26430 82810 26490
rect 82330 26376 82390 26390
rect 82330 26342 82358 26376
rect 82358 26342 82390 26376
rect 82330 26330 82390 26342
rect 82750 26260 82810 26320
rect 83170 26376 83230 26390
rect 83170 26342 83175 26376
rect 83175 26342 83209 26376
rect 83209 26342 83230 26376
rect 83170 26330 83230 26342
rect 83280 25720 83350 25780
rect 83290 25580 83350 25640
rect 82220 25470 82280 25530
rect 82330 24976 82390 24990
rect 82750 25000 82810 25060
rect 82330 24942 82358 24976
rect 82358 24942 82390 24976
rect 82330 24930 82390 24942
rect 83170 24976 83230 24990
rect 83170 24942 83175 24976
rect 83175 24942 83209 24976
rect 83209 24942 83230 24976
rect 83170 24930 83230 24942
rect 82750 24830 82810 24890
rect 82750 24720 82810 24780
rect 82330 24666 82390 24680
rect 82330 24632 82358 24666
rect 82358 24632 82390 24666
rect 82330 24620 82390 24632
rect 82750 24550 82810 24610
rect 83170 24666 83230 24680
rect 83170 24632 83175 24666
rect 83175 24632 83209 24666
rect 83209 24632 83230 24666
rect 83170 24620 83230 24632
rect 83280 24010 83350 24070
rect 83290 23870 83350 23930
rect 82220 23760 82280 23820
rect 82330 23266 82390 23280
rect 82750 23290 82810 23350
rect 82330 23232 82358 23266
rect 82358 23232 82390 23266
rect 82330 23220 82390 23232
rect 83170 23266 83230 23280
rect 83170 23232 83175 23266
rect 83175 23232 83209 23266
rect 83209 23232 83230 23266
rect 83170 23220 83230 23232
rect 82750 23120 82810 23180
rect 82750 23010 82810 23070
rect 82330 22956 82390 22970
rect 82330 22922 82358 22956
rect 82358 22922 82390 22956
rect 82330 22910 82390 22922
rect 82750 22840 82810 22900
rect 83170 22956 83230 22970
rect 83170 22922 83175 22956
rect 83175 22922 83209 22956
rect 83209 22922 83230 22956
rect 83170 22910 83230 22922
rect 83280 22300 83350 22360
rect 83290 22160 83350 22220
rect 82220 22050 82280 22110
rect 82330 21556 82390 21570
rect 82750 21580 82810 21640
rect 82330 21522 82358 21556
rect 82358 21522 82390 21556
rect 82330 21510 82390 21522
rect 83170 21556 83230 21570
rect 83170 21522 83175 21556
rect 83175 21522 83209 21556
rect 83209 21522 83230 21556
rect 83170 21510 83230 21522
rect 82750 21410 82810 21470
rect 82750 21300 82810 21360
rect 82330 21246 82390 21260
rect 82330 21212 82358 21246
rect 82358 21212 82390 21246
rect 82330 21200 82390 21212
rect 82750 21130 82810 21190
rect 83170 21246 83230 21260
rect 83170 21212 83175 21246
rect 83175 21212 83209 21246
rect 83209 21212 83230 21246
rect 83170 21200 83230 21212
rect 83280 20590 83350 20650
rect 83290 20450 83350 20510
rect 82220 20340 82280 20400
rect 82330 19846 82390 19860
rect 82750 19870 82810 19930
rect 82330 19812 82358 19846
rect 82358 19812 82390 19846
rect 82330 19800 82390 19812
rect 83170 19846 83230 19860
rect 83170 19812 83175 19846
rect 83175 19812 83209 19846
rect 83209 19812 83230 19846
rect 83170 19800 83230 19812
rect 82750 19700 82810 19760
rect 82750 19590 82810 19650
rect 82330 19536 82390 19550
rect 82330 19502 82358 19536
rect 82358 19502 82390 19536
rect 82330 19490 82390 19502
rect 82750 19420 82810 19480
rect 83170 19536 83230 19550
rect 83170 19502 83175 19536
rect 83175 19502 83209 19536
rect 83209 19502 83230 19536
rect 83170 19490 83230 19502
rect 83280 18880 83350 18940
rect 83290 18740 83350 18800
rect 82220 18630 82280 18690
rect 82330 18136 82390 18150
rect 82750 18160 82810 18220
rect 82330 18102 82358 18136
rect 82358 18102 82390 18136
rect 82330 18090 82390 18102
rect 83170 18136 83230 18150
rect 83170 18102 83175 18136
rect 83175 18102 83209 18136
rect 83209 18102 83230 18136
rect 83170 18090 83230 18102
rect 82750 17990 82810 18050
rect 82750 17880 82810 17940
rect 82330 17826 82390 17840
rect 82330 17792 82358 17826
rect 82358 17792 82390 17826
rect 82330 17780 82390 17792
rect 82750 17710 82810 17770
rect 83170 17826 83230 17840
rect 83170 17792 83175 17826
rect 83175 17792 83209 17826
rect 83209 17792 83230 17826
rect 83170 17780 83230 17792
rect 83280 17170 83350 17230
rect 83290 17030 83350 17090
rect 82220 16920 82280 16980
rect 82330 16426 82390 16440
rect 82750 16450 82810 16510
rect 82330 16392 82358 16426
rect 82358 16392 82390 16426
rect 82330 16380 82390 16392
rect 83170 16426 83230 16440
rect 83170 16392 83175 16426
rect 83175 16392 83209 16426
rect 83209 16392 83230 16426
rect 83170 16380 83230 16392
rect 82750 16280 82810 16340
rect 82750 16170 82810 16230
rect 82330 16116 82390 16130
rect 82330 16082 82358 16116
rect 82358 16082 82390 16116
rect 82330 16070 82390 16082
rect 82750 16000 82810 16060
rect 83170 16116 83230 16130
rect 83170 16082 83175 16116
rect 83175 16082 83209 16116
rect 83209 16082 83230 16116
rect 83170 16070 83230 16082
rect 83280 15460 83350 15520
rect 83290 15320 83350 15380
rect 82220 15210 82280 15270
rect 82330 14716 82390 14730
rect 82750 14740 82810 14800
rect 82330 14682 82358 14716
rect 82358 14682 82390 14716
rect 82330 14670 82390 14682
rect 83170 14716 83230 14730
rect 83170 14682 83175 14716
rect 83175 14682 83209 14716
rect 83209 14682 83230 14716
rect 83170 14670 83230 14682
rect 82750 14570 82810 14630
rect 82750 14460 82810 14520
rect 82330 14406 82390 14420
rect 82330 14372 82358 14406
rect 82358 14372 82390 14406
rect 82330 14360 82390 14372
rect 82750 14290 82810 14350
rect 83170 14406 83230 14420
rect 83170 14372 83175 14406
rect 83175 14372 83209 14406
rect 83209 14372 83230 14406
rect 83170 14360 83230 14372
rect 83280 13750 83350 13810
rect 83290 13610 83350 13670
rect 82220 13500 82280 13560
rect 82330 13006 82390 13020
rect 82750 13030 82810 13090
rect 82330 12972 82358 13006
rect 82358 12972 82390 13006
rect 82330 12960 82390 12972
rect 83170 13006 83230 13020
rect 83170 12972 83175 13006
rect 83175 12972 83209 13006
rect 83209 12972 83230 13006
rect 83170 12960 83230 12972
rect 82750 12860 82810 12920
rect 82750 12750 82810 12810
rect 82330 12696 82390 12710
rect 82330 12662 82358 12696
rect 82358 12662 82390 12696
rect 82330 12650 82390 12662
rect 82750 12580 82810 12640
rect 83170 12696 83230 12710
rect 83170 12662 83175 12696
rect 83175 12662 83209 12696
rect 83209 12662 83230 12696
rect 83170 12650 83230 12662
rect 83280 12040 83350 12100
rect 83290 11900 83350 11960
rect 82220 11790 82280 11850
rect 82330 11296 82390 11310
rect 82750 11320 82810 11380
rect 82330 11262 82358 11296
rect 82358 11262 82390 11296
rect 82330 11250 82390 11262
rect 83170 11296 83230 11310
rect 83170 11262 83175 11296
rect 83175 11262 83209 11296
rect 83209 11262 83230 11296
rect 83170 11250 83230 11262
rect 82750 11150 82810 11210
rect 82750 11040 82810 11100
rect 82330 10986 82390 11000
rect 82330 10952 82358 10986
rect 82358 10952 82390 10986
rect 82330 10940 82390 10952
rect 82750 10870 82810 10930
rect 83170 10986 83230 11000
rect 83170 10952 83175 10986
rect 83175 10952 83209 10986
rect 83209 10952 83230 10986
rect 83170 10940 83230 10952
rect 83280 10330 83350 10390
rect 83290 10190 83350 10250
rect 82220 10080 82280 10140
rect 82330 9586 82390 9600
rect 82750 9610 82810 9670
rect 82330 9552 82358 9586
rect 82358 9552 82390 9586
rect 82330 9540 82390 9552
rect 83170 9586 83230 9600
rect 83170 9552 83175 9586
rect 83175 9552 83209 9586
rect 83209 9552 83230 9586
rect 83170 9540 83230 9552
rect 82750 9440 82810 9500
rect 82750 9330 82810 9390
rect 82330 9276 82390 9290
rect 82330 9242 82358 9276
rect 82358 9242 82390 9276
rect 82330 9230 82390 9242
rect 82750 9160 82810 9220
rect 83170 9276 83230 9290
rect 83170 9242 83175 9276
rect 83175 9242 83209 9276
rect 83209 9242 83230 9276
rect 83170 9230 83230 9242
rect 83280 8620 83350 8680
rect 83290 8480 83350 8540
rect 82220 8370 82280 8430
rect 82330 7876 82390 7890
rect 82750 7900 82810 7960
rect 82330 7842 82358 7876
rect 82358 7842 82390 7876
rect 82330 7830 82390 7842
rect 83170 7876 83230 7890
rect 83170 7842 83175 7876
rect 83175 7842 83209 7876
rect 83209 7842 83230 7876
rect 83170 7830 83230 7842
rect 82750 7730 82810 7790
rect 82750 7620 82810 7680
rect 82330 7566 82390 7580
rect 82330 7532 82358 7566
rect 82358 7532 82390 7566
rect 82330 7520 82390 7532
rect 82750 7450 82810 7510
rect 83170 7566 83230 7580
rect 83170 7532 83175 7566
rect 83175 7532 83209 7566
rect 83209 7532 83230 7566
rect 83170 7520 83230 7532
rect 83280 6910 83350 6970
rect 83290 6770 83350 6830
rect 82220 6660 82280 6720
rect 82330 6166 82390 6180
rect 82750 6190 82810 6250
rect 82330 6132 82358 6166
rect 82358 6132 82390 6166
rect 82330 6120 82390 6132
rect 83170 6166 83230 6180
rect 83170 6132 83175 6166
rect 83175 6132 83209 6166
rect 83209 6132 83230 6166
rect 83170 6120 83230 6132
rect 82750 6020 82810 6080
rect 82750 5910 82810 5970
rect 82330 5856 82390 5870
rect 82330 5822 82358 5856
rect 82358 5822 82390 5856
rect 82330 5810 82390 5822
rect 82750 5740 82810 5800
rect 83170 5856 83230 5870
rect 83170 5822 83175 5856
rect 83175 5822 83209 5856
rect 83209 5822 83230 5856
rect 83170 5810 83230 5822
rect 83280 5200 83350 5260
rect 83290 5060 83350 5120
rect 82220 4950 82280 5010
rect 82330 4456 82390 4470
rect 82750 4480 82810 4540
rect 82330 4422 82358 4456
rect 82358 4422 82390 4456
rect 82330 4410 82390 4422
rect 83170 4456 83230 4470
rect 83170 4422 83175 4456
rect 83175 4422 83209 4456
rect 83209 4422 83230 4456
rect 83170 4410 83230 4422
rect 82750 4310 82810 4370
rect 82750 4200 82810 4260
rect 82330 4146 82390 4160
rect 82330 4112 82358 4146
rect 82358 4112 82390 4146
rect 82330 4100 82390 4112
rect 82750 4030 82810 4090
rect 83170 4146 83230 4160
rect 83170 4112 83175 4146
rect 83175 4112 83209 4146
rect 83209 4112 83230 4146
rect 83170 4100 83230 4112
rect 83280 3490 83350 3550
rect 83290 3350 83350 3410
rect 82220 3240 82280 3300
rect 82330 2746 82390 2760
rect 82750 2770 82810 2830
rect 82330 2712 82358 2746
rect 82358 2712 82390 2746
rect 82330 2700 82390 2712
rect 83170 2746 83230 2760
rect 83170 2712 83175 2746
rect 83175 2712 83209 2746
rect 83209 2712 83230 2746
rect 83170 2700 83230 2712
rect 82750 2600 82810 2660
rect 82750 2490 82810 2550
rect 82330 2436 82390 2450
rect 82330 2402 82358 2436
rect 82358 2402 82390 2436
rect 82330 2390 82390 2402
rect 82750 2320 82810 2380
rect 83170 2436 83230 2450
rect 83170 2402 83175 2436
rect 83175 2402 83209 2436
rect 83209 2402 83230 2436
rect 83170 2390 83230 2402
rect 83280 1780 83350 1840
rect 83290 1640 83350 1700
rect 82220 1530 82280 1590
rect 82330 1036 82390 1050
rect 82750 1060 82810 1120
rect 82330 1002 82358 1036
rect 82358 1002 82390 1036
rect 82330 990 82390 1002
rect 83170 1036 83230 1050
rect 83170 1002 83175 1036
rect 83175 1002 83209 1036
rect 83209 1002 83230 1036
rect 83170 990 83230 1002
rect 82750 890 82810 950
rect 82750 780 82810 840
rect 82330 726 82390 740
rect 82330 692 82358 726
rect 82358 692 82390 726
rect 82330 680 82390 692
rect 82750 610 82810 670
rect 83170 726 83230 740
rect 83170 692 83175 726
rect 83175 692 83209 726
rect 83209 692 83230 726
rect 83170 680 83230 692
rect 82220 80 82280 140
rect 83280 70 83350 130
rect 83290 -70 83350 -10
rect 82220 -180 82280 -120
rect 82330 -674 82390 -660
rect 82750 -650 82810 -590
rect 82330 -708 82358 -674
rect 82358 -708 82390 -674
rect 82330 -720 82390 -708
rect 83170 -674 83230 -660
rect 83170 -708 83175 -674
rect 83175 -708 83209 -674
rect 83209 -708 83230 -674
rect 83170 -720 83230 -708
rect 82750 -820 82810 -760
rect 82750 -930 82810 -870
rect 82330 -984 82390 -970
rect 82330 -1018 82358 -984
rect 82358 -1018 82390 -984
rect 82330 -1030 82390 -1018
rect 82750 -1100 82810 -1040
rect 83170 -984 83230 -970
rect 83170 -1018 83175 -984
rect 83175 -1018 83209 -984
rect 83209 -1018 83230 -984
rect 83170 -1030 83230 -1018
rect 83280 -1640 83350 -1580
<< metal2 >>
rect 2350 32660 2430 32670
rect 2350 32600 2360 32660
rect 2420 32600 2430 32660
rect 7340 32660 7420 32670
rect 2350 32590 2430 32600
rect 4150 32590 4160 32650
rect 4220 32590 4230 32650
rect -5530 30120 -5430 30140
rect -5530 30060 -5510 30120
rect -5450 30060 -5430 30120
rect -5530 30040 -5430 30060
rect -5110 30120 -5100 30180
rect -5040 30120 -5030 30180
rect -5110 30000 -5080 30120
rect -5250 29990 -5170 30000
rect -5250 29930 -5240 29990
rect -5180 29930 -5170 29990
rect -5250 29920 -5170 29930
rect -5110 29990 -5030 30000
rect -5110 29930 -5100 29990
rect -5040 29930 -5030 29990
rect -5110 29920 -5030 29930
rect -2080 29990 -2000 30000
rect -2080 29930 -2070 29990
rect -2010 29930 -2000 29990
rect -2080 29920 -2000 29930
rect -5370 29850 -5290 29860
rect -5370 29790 -5360 29850
rect -5300 29790 -5290 29850
rect -5370 29780 -5290 29790
rect -2080 29140 -2010 29920
rect 2350 29600 2380 32590
rect 2410 32520 2490 32530
rect 2410 32460 2420 32520
rect 2480 32460 2490 32520
rect 2410 32450 2490 32460
rect 4090 32450 4100 32510
rect 4160 32450 4170 32510
rect 2350 29590 2410 29600
rect 2350 29520 2410 29530
rect 2440 29550 2470 32450
rect 3710 30130 3790 30140
rect 3710 30070 3720 30130
rect 3780 30070 3790 30130
rect 3710 30060 3790 30070
rect 3860 30060 3870 30120
rect 3930 30060 3940 30120
rect 2640 29990 2720 30000
rect 2640 29930 2650 29990
rect 2710 29930 2720 29990
rect 2640 29920 2720 29930
rect 2440 29520 2610 29550
rect -2080 29080 -2070 29140
rect -2010 29080 -2000 29140
rect -2080 29070 -2000 29080
rect 1860 27360 1890 29070
rect 1980 27360 2010 29070
rect 2100 27360 2130 29070
rect 2220 27360 2250 29070
rect 2340 27360 2370 29070
rect 2460 27360 2490 29070
rect 2580 27360 2610 29520
rect 2640 29140 2710 29920
rect 3720 29150 3790 30060
rect 3910 29150 3940 30060
rect 4110 29550 4140 32450
rect 4200 29600 4230 32590
rect 3710 29140 3790 29150
rect 2640 29080 2650 29140
rect 2710 29080 2720 29140
rect 2640 29070 2720 29080
rect 3710 29080 3720 29140
rect 3780 29080 3790 29140
rect 3710 29060 3790 29080
rect 3880 29140 3940 29150
rect 3880 29070 3940 29080
rect 3970 29520 4140 29550
rect 4170 29590 4230 29600
rect 4170 29520 4230 29530
rect 7340 32600 7350 32660
rect 7410 32600 7420 32660
rect 12330 32660 12410 32670
rect 7340 32590 7420 32600
rect 9140 32590 9150 32650
rect 9210 32590 9220 32650
rect 7340 29600 7370 32590
rect 7400 32520 7480 32530
rect 7400 32460 7410 32520
rect 7470 32460 7480 32520
rect 7400 32450 7480 32460
rect 9080 32450 9090 32510
rect 9150 32450 9160 32510
rect 7340 29590 7400 29600
rect 7340 29520 7400 29530
rect 7430 29550 7460 32450
rect 8700 30130 8780 30140
rect 8700 30070 8710 30130
rect 8770 30070 8780 30130
rect 8700 30060 8780 30070
rect 8850 30060 8860 30120
rect 8920 30060 8930 30120
rect 7630 29990 7710 30000
rect 7630 29930 7640 29990
rect 7700 29930 7710 29990
rect 7630 29920 7710 29930
rect 7430 29520 7600 29550
rect 3710 29000 3720 29060
rect 3780 29000 3790 29060
rect 3710 28990 3790 29000
rect 2640 28950 2720 28960
rect 2640 28890 2650 28950
rect 2710 28890 2720 28950
rect 2640 28880 2720 28890
rect 3170 28480 3790 28490
rect 3170 28420 3180 28480
rect 3240 28460 3790 28480
rect 3240 28420 3250 28460
rect 2750 28410 2830 28420
rect 3170 28410 3250 28420
rect 3590 28410 3670 28420
rect 2750 28390 2760 28410
rect 2640 28360 2760 28390
rect 2750 28350 2760 28360
rect 2820 28350 2830 28410
rect 2750 28340 2830 28350
rect 3590 28350 3600 28410
rect 3660 28390 3670 28410
rect 3660 28360 3790 28390
rect 3660 28350 3670 28360
rect 3590 28340 3670 28350
rect 3160 28310 3260 28330
rect 3160 28240 3180 28310
rect 3250 28240 3260 28310
rect 3160 28200 3260 28240
rect 3160 28130 3180 28200
rect 3250 28130 3260 28200
rect 3160 28120 3260 28130
rect 2750 28100 2830 28110
rect 2750 28080 2760 28100
rect 2640 28050 2760 28080
rect 2750 28040 2760 28050
rect 2820 28040 2830 28100
rect 3590 28100 3670 28110
rect 3590 28040 3600 28100
rect 3660 28080 3670 28100
rect 3660 28050 3790 28080
rect 3660 28040 3670 28050
rect 2750 28030 2830 28040
rect 3170 28030 3250 28040
rect 3590 28030 3670 28040
rect 3170 27970 3180 28030
rect 3240 27990 3250 28030
rect 3240 27970 3790 27990
rect 3170 27960 3790 27970
rect 3780 27420 3790 27440
rect 3970 27360 4000 29520
rect 4090 27360 4120 29070
rect 4210 27360 4240 29070
rect 4330 27360 4360 29070
rect 4450 27360 4480 29070
rect 4570 27360 4600 29070
rect 4690 27360 4720 29070
rect 6850 27360 6880 29070
rect 6970 27360 7000 29070
rect 7090 27360 7120 29070
rect 7210 27360 7240 29070
rect 7330 27360 7360 29070
rect 7450 27360 7480 29070
rect 7570 27360 7600 29520
rect 7630 29140 7700 29920
rect 8710 29150 8780 30060
rect 8900 29150 8930 30060
rect 9100 29550 9130 32450
rect 9190 29600 9220 32590
rect 12330 32600 12340 32660
rect 12400 32600 12410 32660
rect 17320 32660 17400 32670
rect 12330 32590 12410 32600
rect 14130 32590 14140 32650
rect 14200 32590 14210 32650
rect 8700 29140 8780 29150
rect 7630 29080 7640 29140
rect 7700 29080 7710 29140
rect 7630 29070 7710 29080
rect 8700 29080 8710 29140
rect 8770 29080 8780 29140
rect 8700 29060 8780 29080
rect 8870 29140 8930 29150
rect 8870 29070 8930 29080
rect 8960 29520 9130 29550
rect 9160 29590 9220 29600
rect 9160 29520 9220 29530
rect 12150 32380 12230 32390
rect 12150 32320 12160 32380
rect 12220 32320 12230 32380
rect 12150 32310 12230 32320
rect 12150 29540 12180 32310
rect 12210 32240 12290 32250
rect 12210 32180 12220 32240
rect 12280 32180 12290 32240
rect 12210 32170 12290 32180
rect 12150 29530 12210 29540
rect 8700 29000 8710 29060
rect 8770 29000 8780 29060
rect 8700 28990 8780 29000
rect 7630 28950 7710 28960
rect 7630 28890 7640 28950
rect 7700 28890 7710 28950
rect 7630 28880 7710 28890
rect 8160 28480 8780 28490
rect 8160 28420 8170 28480
rect 8230 28460 8780 28480
rect 8230 28420 8240 28460
rect 7740 28410 7820 28420
rect 8160 28410 8240 28420
rect 8580 28410 8660 28420
rect 7740 28390 7750 28410
rect 7630 28360 7750 28390
rect 7740 28350 7750 28360
rect 7810 28350 7820 28410
rect 7740 28340 7820 28350
rect 8580 28350 8590 28410
rect 8650 28390 8660 28410
rect 8650 28360 8780 28390
rect 8650 28350 8660 28360
rect 8580 28340 8660 28350
rect 8150 28310 8250 28330
rect 8150 28240 8170 28310
rect 8240 28240 8250 28310
rect 8150 28200 8250 28240
rect 8150 28130 8170 28200
rect 8240 28130 8250 28200
rect 8150 28120 8250 28130
rect 7740 28100 7820 28110
rect 7740 28080 7750 28100
rect 7630 28050 7750 28080
rect 7740 28040 7750 28050
rect 7810 28040 7820 28100
rect 8580 28100 8660 28110
rect 8580 28040 8590 28100
rect 8650 28080 8660 28100
rect 8650 28050 8780 28080
rect 8650 28040 8660 28050
rect 7740 28030 7820 28040
rect 8160 28030 8240 28040
rect 8580 28030 8660 28040
rect 8160 27970 8170 28030
rect 8230 27990 8240 28030
rect 8230 27970 8780 27990
rect 8160 27960 8780 27970
rect 8770 27420 8780 27440
rect 8960 27360 8990 29520
rect 12150 29460 12210 29470
rect 12240 29490 12270 32170
rect 12330 29600 12360 32590
rect 12390 32520 12470 32530
rect 12390 32460 12400 32520
rect 12460 32460 12470 32520
rect 12390 32450 12470 32460
rect 14070 32450 14080 32510
rect 14140 32450 14150 32510
rect 12330 29590 12390 29600
rect 12330 29520 12390 29530
rect 12420 29550 12450 32450
rect 13690 30130 13770 30140
rect 13690 30070 13700 30130
rect 13760 30070 13770 30130
rect 13690 30060 13770 30070
rect 13840 30060 13850 30120
rect 13910 30060 13920 30120
rect 12620 29990 12700 30000
rect 12620 29930 12630 29990
rect 12690 29930 12700 29990
rect 12620 29920 12700 29930
rect 12420 29520 12590 29550
rect 12240 29460 12470 29490
rect 9080 27360 9110 29070
rect 9200 27360 9230 29070
rect 9320 27360 9350 29070
rect 9440 27360 9470 29070
rect 9560 27360 9590 29070
rect 9680 27360 9710 29070
rect 11840 27360 11870 29070
rect 11960 27360 11990 29070
rect 12080 27360 12110 29070
rect 12200 27360 12230 29070
rect 12320 27360 12350 29070
rect 12440 27360 12470 29460
rect 12560 27360 12590 29520
rect 12620 29140 12690 29920
rect 13700 29150 13770 30060
rect 13890 29150 13920 30060
rect 14090 29550 14120 32450
rect 14180 29600 14210 32590
rect 17320 32600 17330 32660
rect 17390 32600 17400 32660
rect 22310 32660 22390 32670
rect 17320 32590 17400 32600
rect 19120 32590 19130 32650
rect 19190 32590 19200 32650
rect 17140 32380 17220 32390
rect 14310 32310 14320 32370
rect 14380 32310 14390 32370
rect 14250 32170 14260 32230
rect 14320 32170 14330 32230
rect 13690 29140 13770 29150
rect 12620 29080 12630 29140
rect 12690 29080 12700 29140
rect 12620 29070 12700 29080
rect 13690 29080 13700 29140
rect 13760 29080 13770 29140
rect 13690 29060 13770 29080
rect 13860 29140 13920 29150
rect 13860 29070 13920 29080
rect 13950 29520 14120 29550
rect 14150 29590 14210 29600
rect 14150 29520 14210 29530
rect 13690 29000 13700 29060
rect 13760 29000 13770 29060
rect 13690 28990 13770 29000
rect 12620 28950 12700 28960
rect 12620 28890 12630 28950
rect 12690 28890 12700 28950
rect 12620 28880 12700 28890
rect 13150 28480 13770 28490
rect 13150 28420 13160 28480
rect 13220 28460 13770 28480
rect 13220 28420 13230 28460
rect 12730 28410 12810 28420
rect 13150 28410 13230 28420
rect 13570 28410 13650 28420
rect 12730 28390 12740 28410
rect 12620 28360 12740 28390
rect 12730 28350 12740 28360
rect 12800 28350 12810 28410
rect 12730 28340 12810 28350
rect 13570 28350 13580 28410
rect 13640 28390 13650 28410
rect 13640 28360 13770 28390
rect 13640 28350 13650 28360
rect 13570 28340 13650 28350
rect 13140 28310 13240 28330
rect 13140 28240 13160 28310
rect 13230 28240 13240 28310
rect 13140 28200 13240 28240
rect 13140 28130 13160 28200
rect 13230 28130 13240 28200
rect 13140 28120 13240 28130
rect 12730 28100 12810 28110
rect 12730 28080 12740 28100
rect 12620 28050 12740 28080
rect 12730 28040 12740 28050
rect 12800 28040 12810 28100
rect 13570 28100 13650 28110
rect 13570 28040 13580 28100
rect 13640 28080 13650 28100
rect 13640 28050 13770 28080
rect 13640 28040 13650 28050
rect 12730 28030 12810 28040
rect 13150 28030 13230 28040
rect 13570 28030 13650 28040
rect 13150 27970 13160 28030
rect 13220 27990 13230 28030
rect 13220 27970 13770 27990
rect 13150 27960 13770 27970
rect 13760 27420 13770 27440
rect 13950 27360 13980 29520
rect 14270 29490 14300 32170
rect 14360 29540 14390 32310
rect 14070 29460 14300 29490
rect 14330 29530 14390 29540
rect 14330 29460 14390 29470
rect 17140 32320 17150 32380
rect 17210 32320 17220 32380
rect 17140 32310 17220 32320
rect 17140 29540 17170 32310
rect 17200 32240 17280 32250
rect 17200 32180 17210 32240
rect 17270 32180 17280 32240
rect 17200 32170 17280 32180
rect 17140 29530 17200 29540
rect 17140 29460 17200 29470
rect 17230 29490 17260 32170
rect 17320 29600 17350 32590
rect 17380 32520 17460 32530
rect 17380 32460 17390 32520
rect 17450 32460 17460 32520
rect 17380 32450 17460 32460
rect 19060 32450 19070 32510
rect 19130 32450 19140 32510
rect 17320 29590 17380 29600
rect 17320 29520 17380 29530
rect 17410 29550 17440 32450
rect 18680 30130 18760 30140
rect 18680 30070 18690 30130
rect 18750 30070 18760 30130
rect 18680 30060 18760 30070
rect 18830 30060 18840 30120
rect 18900 30060 18910 30120
rect 17610 29990 17690 30000
rect 17610 29930 17620 29990
rect 17680 29930 17690 29990
rect 17610 29920 17690 29930
rect 17410 29520 17580 29550
rect 17230 29460 17460 29490
rect 14070 27360 14100 29460
rect 14190 27360 14220 29070
rect 14310 27360 14340 29070
rect 14430 27360 14460 29070
rect 14550 27360 14580 29070
rect 14670 27360 14700 29070
rect 16830 27360 16860 29070
rect 16950 27360 16980 29070
rect 17070 27360 17100 29070
rect 17190 27360 17220 29070
rect 17310 27360 17340 29070
rect 17430 27360 17460 29460
rect 17550 27360 17580 29520
rect 17610 29140 17680 29920
rect 18690 29150 18760 30060
rect 18880 29150 18910 30060
rect 19080 29550 19110 32450
rect 19170 29600 19200 32590
rect 22310 32600 22320 32660
rect 22380 32600 22390 32660
rect 27300 32660 27380 32670
rect 22310 32590 22390 32600
rect 24110 32590 24120 32650
rect 24180 32590 24190 32650
rect 22130 32380 22210 32390
rect 19300 32310 19310 32370
rect 19370 32310 19380 32370
rect 19240 32170 19250 32230
rect 19310 32170 19320 32230
rect 18680 29140 18760 29150
rect 17610 29080 17620 29140
rect 17680 29080 17690 29140
rect 17610 29070 17690 29080
rect 18680 29080 18690 29140
rect 18750 29080 18760 29140
rect 18680 29060 18760 29080
rect 18850 29140 18910 29150
rect 18850 29070 18910 29080
rect 18940 29520 19110 29550
rect 19140 29590 19200 29600
rect 19140 29520 19200 29530
rect 18680 29000 18690 29060
rect 18750 29000 18760 29060
rect 18680 28990 18760 29000
rect 17610 28950 17690 28960
rect 17610 28890 17620 28950
rect 17680 28890 17690 28950
rect 17610 28880 17690 28890
rect 18140 28480 18760 28490
rect 18140 28420 18150 28480
rect 18210 28460 18760 28480
rect 18210 28420 18220 28460
rect 17720 28410 17800 28420
rect 18140 28410 18220 28420
rect 18560 28410 18640 28420
rect 17720 28390 17730 28410
rect 17610 28360 17730 28390
rect 17720 28350 17730 28360
rect 17790 28350 17800 28410
rect 17720 28340 17800 28350
rect 18560 28350 18570 28410
rect 18630 28390 18640 28410
rect 18630 28360 18760 28390
rect 18630 28350 18640 28360
rect 18560 28340 18640 28350
rect 18130 28310 18230 28330
rect 18130 28240 18150 28310
rect 18220 28240 18230 28310
rect 18130 28200 18230 28240
rect 18130 28130 18150 28200
rect 18220 28130 18230 28200
rect 18130 28120 18230 28130
rect 17720 28100 17800 28110
rect 17720 28080 17730 28100
rect 17610 28050 17730 28080
rect 17720 28040 17730 28050
rect 17790 28040 17800 28100
rect 18560 28100 18640 28110
rect 18560 28040 18570 28100
rect 18630 28080 18640 28100
rect 18630 28050 18760 28080
rect 18630 28040 18640 28050
rect 17720 28030 17800 28040
rect 18140 28030 18220 28040
rect 18560 28030 18640 28040
rect 18140 27970 18150 28030
rect 18210 27990 18220 28030
rect 18210 27970 18760 27990
rect 18140 27960 18760 27970
rect 18750 27420 18760 27440
rect 18940 27360 18970 29520
rect 19260 29490 19290 32170
rect 19350 29540 19380 32310
rect 22130 32320 22140 32380
rect 22200 32320 22210 32380
rect 22130 32310 22210 32320
rect 19060 29460 19290 29490
rect 19320 29530 19380 29540
rect 19320 29460 19380 29470
rect 21770 32100 21850 32110
rect 21770 32040 21780 32100
rect 21840 32040 21850 32100
rect 21770 32030 21850 32040
rect 19060 27360 19090 29460
rect 21770 29420 21800 32030
rect 21830 31960 21910 31970
rect 21830 31900 21840 31960
rect 21900 31900 21910 31960
rect 21830 31890 21910 31900
rect 21770 29410 21830 29420
rect 21770 29340 21830 29350
rect 21860 29370 21890 31890
rect 21950 31820 22030 31830
rect 21950 31760 21960 31820
rect 22020 31760 22030 31820
rect 21950 31750 22030 31760
rect 21950 29480 21980 31750
rect 22010 31680 22090 31690
rect 22010 31620 22020 31680
rect 22080 31620 22090 31680
rect 22010 31610 22090 31620
rect 21950 29470 22010 29480
rect 21950 29400 22010 29410
rect 22040 29430 22070 31610
rect 22130 29540 22160 32310
rect 22190 32240 22270 32250
rect 22190 32180 22200 32240
rect 22260 32180 22270 32240
rect 22190 32170 22270 32180
rect 22130 29530 22190 29540
rect 22130 29460 22190 29470
rect 22220 29490 22250 32170
rect 22310 29600 22340 32590
rect 22370 32520 22450 32530
rect 22370 32460 22380 32520
rect 22440 32460 22450 32520
rect 22370 32450 22450 32460
rect 24050 32450 24060 32510
rect 24120 32450 24130 32510
rect 22310 29590 22370 29600
rect 22310 29520 22370 29530
rect 22400 29550 22430 32450
rect 23670 30130 23750 30140
rect 23670 30070 23680 30130
rect 23740 30070 23750 30130
rect 23670 30060 23750 30070
rect 23820 30060 23830 30120
rect 23890 30060 23900 30120
rect 22600 29990 22680 30000
rect 22600 29930 22610 29990
rect 22670 29930 22680 29990
rect 22600 29920 22680 29930
rect 22400 29520 22570 29550
rect 22220 29460 22450 29490
rect 22040 29400 22330 29430
rect 21860 29340 22210 29370
rect 19180 27360 19210 29070
rect 19300 27360 19330 29070
rect 19420 27360 19450 29070
rect 19540 27360 19570 29070
rect 19660 27360 19690 29070
rect 21820 27360 21850 29070
rect 21940 27360 21970 29070
rect 22060 27360 22090 29070
rect 22180 27360 22210 29340
rect 22300 27360 22330 29400
rect 22420 27360 22450 29460
rect 22540 27360 22570 29520
rect 22600 29140 22670 29920
rect 23680 29150 23750 30060
rect 23870 29150 23900 30060
rect 24070 29550 24100 32450
rect 24160 29600 24190 32590
rect 27300 32600 27310 32660
rect 27370 32600 27380 32660
rect 32290 32660 32370 32670
rect 27300 32590 27380 32600
rect 29100 32590 29110 32650
rect 29170 32590 29180 32650
rect 27120 32380 27200 32390
rect 24290 32310 24300 32370
rect 24360 32310 24370 32370
rect 24230 32170 24240 32230
rect 24300 32170 24310 32230
rect 23670 29140 23750 29150
rect 22600 29080 22610 29140
rect 22670 29080 22680 29140
rect 22600 29070 22680 29080
rect 23670 29080 23680 29140
rect 23740 29080 23750 29140
rect 23670 29060 23750 29080
rect 23840 29140 23900 29150
rect 23840 29070 23900 29080
rect 23930 29520 24100 29550
rect 24130 29590 24190 29600
rect 24130 29520 24190 29530
rect 23670 29000 23680 29060
rect 23740 29000 23750 29060
rect 23670 28990 23750 29000
rect 22600 28950 22680 28960
rect 22600 28890 22610 28950
rect 22670 28890 22680 28950
rect 22600 28880 22680 28890
rect 23130 28480 23750 28490
rect 23130 28420 23140 28480
rect 23200 28460 23750 28480
rect 23200 28420 23210 28460
rect 22710 28410 22790 28420
rect 23130 28410 23210 28420
rect 23550 28410 23630 28420
rect 22710 28390 22720 28410
rect 22600 28360 22720 28390
rect 22710 28350 22720 28360
rect 22780 28350 22790 28410
rect 22710 28340 22790 28350
rect 23550 28350 23560 28410
rect 23620 28390 23630 28410
rect 23620 28360 23750 28390
rect 23620 28350 23630 28360
rect 23550 28340 23630 28350
rect 23120 28310 23220 28330
rect 23120 28240 23140 28310
rect 23210 28240 23220 28310
rect 23120 28200 23220 28240
rect 23120 28130 23140 28200
rect 23210 28130 23220 28200
rect 23120 28120 23220 28130
rect 22710 28100 22790 28110
rect 22710 28080 22720 28100
rect 22600 28050 22720 28080
rect 22710 28040 22720 28050
rect 22780 28040 22790 28100
rect 23550 28100 23630 28110
rect 23550 28040 23560 28100
rect 23620 28080 23630 28100
rect 23620 28050 23750 28080
rect 23620 28040 23630 28050
rect 22710 28030 22790 28040
rect 23130 28030 23210 28040
rect 23550 28030 23630 28040
rect 23130 27970 23140 28030
rect 23200 27990 23210 28030
rect 23200 27970 23750 27990
rect 23130 27960 23750 27970
rect 23740 27420 23750 27440
rect 23930 27360 23960 29520
rect 24250 29490 24280 32170
rect 24340 29540 24370 32310
rect 27120 32320 27130 32380
rect 27190 32320 27200 32380
rect 27120 32310 27200 32320
rect 26760 32100 26840 32110
rect 24650 32030 24660 32090
rect 24720 32030 24730 32090
rect 24590 31890 24600 31950
rect 24660 31890 24670 31950
rect 24470 31750 24480 31810
rect 24540 31750 24550 31810
rect 24410 31610 24420 31670
rect 24480 31610 24490 31670
rect 24050 29460 24280 29490
rect 24310 29530 24370 29540
rect 24310 29460 24370 29470
rect 24050 27360 24080 29460
rect 24430 29430 24460 31610
rect 24520 29480 24550 31750
rect 24170 29400 24460 29430
rect 24490 29470 24550 29480
rect 24490 29400 24550 29410
rect 24170 27360 24200 29400
rect 24610 29370 24640 31890
rect 24700 29420 24730 32030
rect 24290 29340 24640 29370
rect 24670 29410 24730 29420
rect 24670 29340 24730 29350
rect 26760 32040 26770 32100
rect 26830 32040 26840 32100
rect 26760 32030 26840 32040
rect 26760 29420 26790 32030
rect 26820 31960 26900 31970
rect 26820 31900 26830 31960
rect 26890 31900 26900 31960
rect 26820 31890 26900 31900
rect 26760 29410 26820 29420
rect 26760 29340 26820 29350
rect 26850 29370 26880 31890
rect 26940 31820 27020 31830
rect 26940 31760 26950 31820
rect 27010 31760 27020 31820
rect 26940 31750 27020 31760
rect 26940 29480 26970 31750
rect 27000 31680 27080 31690
rect 27000 31620 27010 31680
rect 27070 31620 27080 31680
rect 27000 31610 27080 31620
rect 26940 29470 27000 29480
rect 26940 29400 27000 29410
rect 27030 29430 27060 31610
rect 27120 29540 27150 32310
rect 27180 32240 27260 32250
rect 27180 32180 27190 32240
rect 27250 32180 27260 32240
rect 27180 32170 27260 32180
rect 27120 29530 27180 29540
rect 27120 29460 27180 29470
rect 27210 29490 27240 32170
rect 27300 29600 27330 32590
rect 27360 32520 27440 32530
rect 27360 32460 27370 32520
rect 27430 32460 27440 32520
rect 27360 32450 27440 32460
rect 29040 32450 29050 32510
rect 29110 32450 29120 32510
rect 27300 29590 27360 29600
rect 27300 29520 27360 29530
rect 27390 29550 27420 32450
rect 28660 30130 28740 30140
rect 28660 30070 28670 30130
rect 28730 30070 28740 30130
rect 28660 30060 28740 30070
rect 28810 30060 28820 30120
rect 28880 30060 28890 30120
rect 27590 29990 27670 30000
rect 27590 29930 27600 29990
rect 27660 29930 27670 29990
rect 27590 29920 27670 29930
rect 27390 29520 27560 29550
rect 27210 29460 27440 29490
rect 27030 29400 27320 29430
rect 26850 29340 27200 29370
rect 24290 27360 24320 29340
rect 24410 27360 24440 29070
rect 24530 27360 24560 29070
rect 24650 27360 24680 29070
rect 26810 27360 26840 29070
rect 26930 27360 26960 29070
rect 27050 27360 27080 29070
rect 27170 27360 27200 29340
rect 27290 27360 27320 29400
rect 27410 27360 27440 29460
rect 27530 27360 27560 29520
rect 27590 29140 27660 29920
rect 28670 29150 28740 30060
rect 28860 29150 28890 30060
rect 29060 29550 29090 32450
rect 29150 29600 29180 32590
rect 32290 32600 32300 32660
rect 32360 32600 32370 32660
rect 37280 32660 37360 32670
rect 32290 32590 32370 32600
rect 34090 32590 34100 32650
rect 34160 32590 34170 32650
rect 32110 32380 32190 32390
rect 29280 32310 29290 32370
rect 29350 32310 29360 32370
rect 29220 32170 29230 32230
rect 29290 32170 29300 32230
rect 28660 29140 28740 29150
rect 27590 29080 27600 29140
rect 27660 29080 27670 29140
rect 27590 29070 27670 29080
rect 28660 29080 28670 29140
rect 28730 29080 28740 29140
rect 28660 29060 28740 29080
rect 28830 29140 28890 29150
rect 28830 29070 28890 29080
rect 28920 29520 29090 29550
rect 29120 29590 29180 29600
rect 29120 29520 29180 29530
rect 28660 29000 28670 29060
rect 28730 29000 28740 29060
rect 28660 28990 28740 29000
rect 27590 28950 27670 28960
rect 27590 28890 27600 28950
rect 27660 28890 27670 28950
rect 27590 28880 27670 28890
rect 28120 28480 28740 28490
rect 28120 28420 28130 28480
rect 28190 28460 28740 28480
rect 28190 28420 28200 28460
rect 27700 28410 27780 28420
rect 28120 28410 28200 28420
rect 28540 28410 28620 28420
rect 27700 28390 27710 28410
rect 27590 28360 27710 28390
rect 27700 28350 27710 28360
rect 27770 28350 27780 28410
rect 27700 28340 27780 28350
rect 28540 28350 28550 28410
rect 28610 28390 28620 28410
rect 28610 28360 28740 28390
rect 28610 28350 28620 28360
rect 28540 28340 28620 28350
rect 28110 28310 28210 28330
rect 28110 28240 28130 28310
rect 28200 28240 28210 28310
rect 28110 28200 28210 28240
rect 28110 28130 28130 28200
rect 28200 28130 28210 28200
rect 28110 28120 28210 28130
rect 27700 28100 27780 28110
rect 27700 28080 27710 28100
rect 27590 28050 27710 28080
rect 27700 28040 27710 28050
rect 27770 28040 27780 28100
rect 28540 28100 28620 28110
rect 28540 28040 28550 28100
rect 28610 28080 28620 28100
rect 28610 28050 28740 28080
rect 28610 28040 28620 28050
rect 27700 28030 27780 28040
rect 28120 28030 28200 28040
rect 28540 28030 28620 28040
rect 28120 27970 28130 28030
rect 28190 27990 28200 28030
rect 28190 27970 28740 27990
rect 28120 27960 28740 27970
rect 28730 27420 28740 27440
rect 28920 27360 28950 29520
rect 29240 29490 29270 32170
rect 29330 29540 29360 32310
rect 32110 32320 32120 32380
rect 32180 32320 32190 32380
rect 32110 32310 32190 32320
rect 31930 32100 32010 32110
rect 29640 32030 29650 32090
rect 29710 32030 29720 32090
rect 29580 31890 29590 31950
rect 29650 31890 29660 31950
rect 29460 31750 29470 31810
rect 29530 31750 29540 31810
rect 29400 31610 29410 31670
rect 29470 31610 29480 31670
rect 29040 29460 29270 29490
rect 29300 29530 29360 29540
rect 29300 29460 29360 29470
rect 29040 27360 29070 29460
rect 29420 29430 29450 31610
rect 29510 29480 29540 31750
rect 29160 29400 29450 29430
rect 29480 29470 29540 29480
rect 29480 29400 29540 29410
rect 29160 27360 29190 29400
rect 29600 29370 29630 31890
rect 29690 29420 29720 32030
rect 31930 32040 31940 32100
rect 32000 32040 32010 32100
rect 31930 32030 32010 32040
rect 31750 31820 31830 31830
rect 31750 31760 31760 31820
rect 31820 31760 31830 31820
rect 31750 31750 31830 31760
rect 29280 29340 29630 29370
rect 29660 29410 29720 29420
rect 29660 29340 29720 29350
rect 31390 31540 31470 31550
rect 31390 31480 31400 31540
rect 31460 31480 31470 31540
rect 31390 31470 31470 31480
rect 29280 27360 29310 29340
rect 31390 29300 31420 31470
rect 31450 31400 31530 31410
rect 31450 31340 31460 31400
rect 31520 31340 31530 31400
rect 31450 31330 31530 31340
rect 31390 29290 31450 29300
rect 31390 29220 31450 29230
rect 31480 29250 31510 31330
rect 31570 31260 31650 31270
rect 31570 31200 31580 31260
rect 31640 31200 31650 31260
rect 31570 31190 31650 31200
rect 31570 29360 31600 31190
rect 31630 31120 31710 31130
rect 31630 31060 31640 31120
rect 31700 31060 31710 31120
rect 31630 31050 31710 31060
rect 31570 29350 31630 29360
rect 31570 29280 31630 29290
rect 31660 29310 31690 31050
rect 31750 29420 31780 31750
rect 31810 31680 31890 31690
rect 31810 31620 31820 31680
rect 31880 31620 31890 31680
rect 31810 31610 31890 31620
rect 31750 29410 31810 29420
rect 31750 29340 31810 29350
rect 31840 29370 31870 31610
rect 31930 29480 31960 32030
rect 31990 31960 32070 31970
rect 31990 31900 32000 31960
rect 32060 31900 32070 31960
rect 31990 31890 32070 31900
rect 31930 29470 31990 29480
rect 31930 29400 31990 29410
rect 32020 29430 32050 31890
rect 32110 29540 32140 32310
rect 32170 32240 32250 32250
rect 32170 32180 32180 32240
rect 32240 32180 32250 32240
rect 32170 32170 32250 32180
rect 32110 29530 32170 29540
rect 32110 29460 32170 29470
rect 32200 29490 32230 32170
rect 32290 29600 32320 32590
rect 32350 32520 32430 32530
rect 32350 32460 32360 32520
rect 32420 32460 32430 32520
rect 32350 32450 32430 32460
rect 34030 32450 34040 32510
rect 34100 32450 34110 32510
rect 32290 29590 32350 29600
rect 32290 29520 32350 29530
rect 32380 29550 32410 32450
rect 33650 30130 33730 30140
rect 33650 30070 33660 30130
rect 33720 30070 33730 30130
rect 33650 30060 33730 30070
rect 33800 30060 33810 30120
rect 33870 30060 33880 30120
rect 32580 29990 32660 30000
rect 32580 29930 32590 29990
rect 32650 29930 32660 29990
rect 32580 29920 32660 29930
rect 32380 29520 32550 29550
rect 32200 29460 32430 29490
rect 32020 29400 32310 29430
rect 31840 29340 32190 29370
rect 31660 29280 32070 29310
rect 31480 29220 31950 29250
rect 29400 27360 29430 29070
rect 29520 27360 29550 29070
rect 29640 27360 29670 29070
rect 31800 27360 31830 29070
rect 31920 27360 31950 29220
rect 32040 27360 32070 29280
rect 32160 27360 32190 29340
rect 32280 27360 32310 29400
rect 32400 27360 32430 29460
rect 32520 27360 32550 29520
rect 32580 29140 32650 29920
rect 33660 29150 33730 30060
rect 33850 29150 33880 30060
rect 34050 29550 34080 32450
rect 34140 29600 34170 32590
rect 37280 32600 37290 32660
rect 37350 32600 37360 32660
rect 42270 32660 42350 32670
rect 37280 32590 37360 32600
rect 39080 32590 39090 32650
rect 39150 32590 39160 32650
rect 37100 32380 37180 32390
rect 34270 32310 34280 32370
rect 34340 32310 34350 32370
rect 34210 32170 34220 32230
rect 34280 32170 34290 32230
rect 33650 29140 33730 29150
rect 32580 29080 32590 29140
rect 32650 29080 32660 29140
rect 32580 29070 32660 29080
rect 33650 29080 33660 29140
rect 33720 29080 33730 29140
rect 33650 29060 33730 29080
rect 33820 29140 33880 29150
rect 33820 29070 33880 29080
rect 33910 29520 34080 29550
rect 34110 29590 34170 29600
rect 34110 29520 34170 29530
rect 33650 29000 33660 29060
rect 33720 29000 33730 29060
rect 33650 28990 33730 29000
rect 32580 28950 32660 28960
rect 32580 28890 32590 28950
rect 32650 28890 32660 28950
rect 32580 28880 32660 28890
rect 33110 28480 33730 28490
rect 33110 28420 33120 28480
rect 33180 28460 33730 28480
rect 33180 28420 33190 28460
rect 32690 28410 32770 28420
rect 33110 28410 33190 28420
rect 33530 28410 33610 28420
rect 32690 28390 32700 28410
rect 32580 28360 32700 28390
rect 32690 28350 32700 28360
rect 32760 28350 32770 28410
rect 32690 28340 32770 28350
rect 33530 28350 33540 28410
rect 33600 28390 33610 28410
rect 33600 28360 33730 28390
rect 33600 28350 33610 28360
rect 33530 28340 33610 28350
rect 33100 28310 33200 28330
rect 33100 28240 33120 28310
rect 33190 28240 33200 28310
rect 33100 28200 33200 28240
rect 33100 28130 33120 28200
rect 33190 28130 33200 28200
rect 33100 28120 33200 28130
rect 32690 28100 32770 28110
rect 32690 28080 32700 28100
rect 32580 28050 32700 28080
rect 32690 28040 32700 28050
rect 32760 28040 32770 28100
rect 33530 28100 33610 28110
rect 33530 28040 33540 28100
rect 33600 28080 33610 28100
rect 33600 28050 33730 28080
rect 33600 28040 33610 28050
rect 32690 28030 32770 28040
rect 33110 28030 33190 28040
rect 33530 28030 33610 28040
rect 33110 27970 33120 28030
rect 33180 27990 33190 28030
rect 33180 27970 33730 27990
rect 33110 27960 33730 27970
rect 33720 27420 33730 27440
rect 33910 27360 33940 29520
rect 34230 29490 34260 32170
rect 34320 29540 34350 32310
rect 37100 32320 37110 32380
rect 37170 32320 37180 32380
rect 37100 32310 37180 32320
rect 36920 32100 37000 32110
rect 34450 32030 34460 32090
rect 34520 32030 34530 32090
rect 34390 31890 34400 31950
rect 34460 31890 34470 31950
rect 34030 29460 34260 29490
rect 34290 29530 34350 29540
rect 34290 29460 34350 29470
rect 34030 27360 34060 29460
rect 34410 29430 34440 31890
rect 34500 29480 34530 32030
rect 36920 32040 36930 32100
rect 36990 32040 37000 32100
rect 36920 32030 37000 32040
rect 36740 31820 36820 31830
rect 34630 31750 34640 31810
rect 34700 31750 34710 31810
rect 34570 31610 34580 31670
rect 34640 31610 34650 31670
rect 34150 29400 34440 29430
rect 34470 29470 34530 29480
rect 34470 29400 34530 29410
rect 34150 27360 34180 29400
rect 34590 29370 34620 31610
rect 34680 29420 34710 31750
rect 36740 31760 36750 31820
rect 36810 31760 36820 31820
rect 36740 31750 36820 31760
rect 36560 31540 36640 31550
rect 34990 31470 35000 31530
rect 35060 31470 35070 31530
rect 34930 31330 34940 31390
rect 35000 31330 35010 31390
rect 34810 31190 34820 31250
rect 34880 31190 34890 31250
rect 34750 31050 34760 31110
rect 34820 31050 34830 31110
rect 34270 29340 34620 29370
rect 34650 29410 34710 29420
rect 34650 29340 34710 29350
rect 34270 27360 34300 29340
rect 34770 29310 34800 31050
rect 34860 29360 34890 31190
rect 34390 29280 34800 29310
rect 34830 29350 34890 29360
rect 34830 29280 34890 29290
rect 34390 27360 34420 29280
rect 34950 29250 34980 31330
rect 35040 29300 35070 31470
rect 36560 31480 36570 31540
rect 36630 31480 36640 31540
rect 36560 31470 36640 31480
rect 36380 30980 36460 30990
rect 36380 30920 36390 30980
rect 36450 30920 36460 30980
rect 36380 30910 36460 30920
rect 34510 29220 34980 29250
rect 35010 29290 35070 29300
rect 35010 29220 35070 29230
rect 36200 30420 36280 30430
rect 36200 30360 36210 30420
rect 36270 30360 36280 30420
rect 36200 30350 36280 30360
rect 36200 29240 36230 30350
rect 36260 30280 36340 30290
rect 36260 30220 36270 30280
rect 36330 30220 36340 30280
rect 36260 30210 36340 30220
rect 36200 29230 36260 29240
rect 34510 27360 34540 29220
rect 36200 29160 36260 29170
rect 36290 29190 36320 30210
rect 36380 29300 36410 30910
rect 36440 30840 36520 30850
rect 36440 30780 36450 30840
rect 36510 30780 36520 30840
rect 36440 30770 36520 30780
rect 36380 29290 36440 29300
rect 36380 29220 36440 29230
rect 36470 29250 36500 30770
rect 36560 29360 36590 31470
rect 36620 31400 36700 31410
rect 36620 31340 36630 31400
rect 36690 31340 36700 31400
rect 36620 31330 36700 31340
rect 36560 29350 36620 29360
rect 36560 29280 36620 29290
rect 36650 29310 36680 31330
rect 36740 29420 36770 31750
rect 36800 31680 36880 31690
rect 36800 31620 36810 31680
rect 36870 31620 36880 31680
rect 36800 31610 36880 31620
rect 36740 29410 36800 29420
rect 36740 29340 36800 29350
rect 36830 29370 36860 31610
rect 36920 29480 36950 32030
rect 36980 31960 37060 31970
rect 36980 31900 36990 31960
rect 37050 31900 37060 31960
rect 36980 31890 37060 31900
rect 36920 29470 36980 29480
rect 36920 29400 36980 29410
rect 37010 29430 37040 31890
rect 37100 29540 37130 32310
rect 37160 32240 37240 32250
rect 37160 32180 37170 32240
rect 37230 32180 37240 32240
rect 37160 32170 37240 32180
rect 37100 29530 37160 29540
rect 37100 29460 37160 29470
rect 37190 29490 37220 32170
rect 37280 29600 37310 32590
rect 37340 32520 37420 32530
rect 37340 32460 37350 32520
rect 37410 32460 37420 32520
rect 37340 32450 37420 32460
rect 39020 32450 39030 32510
rect 39090 32450 39100 32510
rect 37280 29590 37340 29600
rect 37280 29520 37340 29530
rect 37370 29550 37400 32450
rect 38640 30130 38720 30140
rect 38640 30070 38650 30130
rect 38710 30070 38720 30130
rect 38640 30060 38720 30070
rect 38790 30060 38800 30120
rect 38860 30060 38870 30120
rect 37570 29990 37650 30000
rect 37570 29930 37580 29990
rect 37640 29930 37650 29990
rect 37570 29920 37650 29930
rect 37370 29520 37540 29550
rect 37190 29460 37420 29490
rect 37010 29400 37300 29430
rect 36830 29340 37180 29370
rect 36650 29280 37060 29310
rect 36470 29220 36940 29250
rect 36290 29160 36820 29190
rect 34630 27360 34660 29070
rect 36790 27360 36820 29160
rect 36910 27360 36940 29220
rect 37030 27360 37060 29280
rect 37150 27360 37180 29340
rect 37270 27360 37300 29400
rect 37390 27360 37420 29460
rect 37510 27360 37540 29520
rect 37570 29140 37640 29920
rect 38650 29150 38720 30060
rect 38840 29150 38870 30060
rect 39040 29550 39070 32450
rect 39130 29600 39160 32590
rect 42270 32600 42280 32660
rect 42340 32600 42350 32660
rect 47260 32660 47340 32670
rect 42270 32590 42350 32600
rect 44070 32590 44080 32650
rect 44140 32590 44150 32650
rect 42090 32380 42170 32390
rect 39260 32310 39270 32370
rect 39330 32310 39340 32370
rect 39200 32170 39210 32230
rect 39270 32170 39280 32230
rect 38640 29140 38720 29150
rect 37570 29080 37580 29140
rect 37640 29080 37650 29140
rect 37570 29070 37650 29080
rect 38640 29080 38650 29140
rect 38710 29080 38720 29140
rect 38640 29060 38720 29080
rect 38810 29140 38870 29150
rect 38810 29070 38870 29080
rect 38900 29520 39070 29550
rect 39100 29590 39160 29600
rect 39100 29520 39160 29530
rect 38640 29000 38650 29060
rect 38710 29000 38720 29060
rect 38640 28990 38720 29000
rect 37570 28950 37650 28960
rect 37570 28890 37580 28950
rect 37640 28890 37650 28950
rect 37570 28880 37650 28890
rect 38100 28480 38720 28490
rect 38100 28420 38110 28480
rect 38170 28460 38720 28480
rect 38170 28420 38180 28460
rect 37680 28410 37760 28420
rect 38100 28410 38180 28420
rect 38520 28410 38600 28420
rect 37680 28390 37690 28410
rect 37570 28360 37690 28390
rect 37680 28350 37690 28360
rect 37750 28350 37760 28410
rect 37680 28340 37760 28350
rect 38520 28350 38530 28410
rect 38590 28390 38600 28410
rect 38590 28360 38720 28390
rect 38590 28350 38600 28360
rect 38520 28340 38600 28350
rect 38090 28310 38190 28330
rect 38090 28240 38110 28310
rect 38180 28240 38190 28310
rect 38090 28200 38190 28240
rect 38090 28130 38110 28200
rect 38180 28130 38190 28200
rect 38090 28120 38190 28130
rect 37680 28100 37760 28110
rect 37680 28080 37690 28100
rect 37570 28050 37690 28080
rect 37680 28040 37690 28050
rect 37750 28040 37760 28100
rect 38520 28100 38600 28110
rect 38520 28040 38530 28100
rect 38590 28080 38600 28100
rect 38590 28050 38720 28080
rect 38590 28040 38600 28050
rect 37680 28030 37760 28040
rect 38100 28030 38180 28040
rect 38520 28030 38600 28040
rect 38100 27970 38110 28030
rect 38170 27990 38180 28030
rect 38170 27970 38720 27990
rect 38100 27960 38720 27970
rect 38710 27420 38720 27440
rect 38900 27360 38930 29520
rect 39220 29490 39250 32170
rect 39310 29540 39340 32310
rect 42090 32320 42100 32380
rect 42160 32320 42170 32380
rect 42090 32310 42170 32320
rect 41910 32100 41990 32110
rect 39440 32030 39450 32090
rect 39510 32030 39520 32090
rect 39380 31890 39390 31950
rect 39450 31890 39460 31950
rect 39020 29460 39250 29490
rect 39280 29530 39340 29540
rect 39280 29460 39340 29470
rect 39020 27360 39050 29460
rect 39400 29430 39430 31890
rect 39490 29480 39520 32030
rect 41910 32040 41920 32100
rect 41980 32040 41990 32100
rect 41910 32030 41990 32040
rect 41730 31820 41810 31830
rect 39620 31750 39630 31810
rect 39690 31750 39700 31810
rect 39560 31610 39570 31670
rect 39630 31610 39640 31670
rect 39140 29400 39430 29430
rect 39460 29470 39520 29480
rect 39460 29400 39520 29410
rect 39140 27360 39170 29400
rect 39580 29370 39610 31610
rect 39670 29420 39700 31750
rect 41730 31760 41740 31820
rect 41800 31760 41810 31820
rect 41730 31750 41810 31760
rect 41550 31540 41630 31550
rect 39800 31470 39810 31530
rect 39870 31470 39880 31530
rect 39740 31330 39750 31390
rect 39810 31330 39820 31390
rect 39260 29340 39610 29370
rect 39640 29410 39700 29420
rect 39640 29340 39700 29350
rect 39260 27360 39290 29340
rect 39760 29310 39790 31330
rect 39850 29360 39880 31470
rect 41550 31480 41560 31540
rect 41620 31480 41630 31540
rect 41550 31470 41630 31480
rect 41190 30980 41270 30990
rect 39980 30910 39990 30970
rect 40050 30910 40060 30970
rect 39920 30770 39930 30830
rect 39990 30770 40000 30830
rect 39380 29280 39790 29310
rect 39820 29350 39880 29360
rect 39820 29280 39880 29290
rect 39380 27360 39410 29280
rect 39940 29250 39970 30770
rect 40030 29300 40060 30910
rect 41190 30920 41200 30980
rect 41260 30920 41270 30980
rect 41190 30910 41270 30920
rect 40160 30350 40170 30410
rect 40230 30350 40240 30410
rect 40090 30210 40100 30270
rect 40160 30210 40170 30270
rect 39500 29220 39970 29250
rect 40000 29290 40060 29300
rect 40000 29220 40060 29230
rect 39500 27360 39530 29220
rect 40120 29190 40150 30210
rect 40210 29240 40240 30350
rect 39620 29160 40150 29190
rect 40180 29230 40240 29240
rect 40180 29160 40240 29170
rect 41190 29240 41220 30910
rect 41250 30840 41330 30850
rect 41250 30780 41260 30840
rect 41320 30780 41330 30840
rect 41250 30770 41330 30780
rect 41190 29230 41250 29240
rect 41190 29160 41250 29170
rect 41280 29190 41310 30770
rect 41340 30700 41420 30710
rect 41340 30640 41350 30700
rect 41410 30640 41420 30700
rect 41340 30630 41420 30640
rect 41370 29300 41400 30630
rect 41430 30560 41510 30570
rect 41430 30500 41440 30560
rect 41500 30500 41510 30560
rect 41430 30490 41510 30500
rect 41370 29290 41430 29300
rect 41370 29220 41430 29230
rect 41460 29250 41490 30490
rect 41550 29360 41580 31470
rect 41610 31400 41690 31410
rect 41610 31340 41620 31400
rect 41680 31340 41690 31400
rect 41610 31330 41690 31340
rect 41550 29350 41610 29360
rect 41550 29280 41610 29290
rect 41640 29310 41670 31330
rect 41730 29420 41760 31750
rect 41790 31680 41870 31690
rect 41790 31620 41800 31680
rect 41860 31620 41870 31680
rect 41790 31610 41870 31620
rect 41730 29410 41790 29420
rect 41730 29340 41790 29350
rect 41820 29370 41850 31610
rect 41910 29480 41940 32030
rect 41970 31960 42050 31970
rect 41970 31900 41980 31960
rect 42040 31900 42050 31960
rect 41970 31890 42050 31900
rect 41910 29470 41970 29480
rect 41910 29400 41970 29410
rect 42000 29430 42030 31890
rect 42090 29540 42120 32310
rect 42150 32240 42230 32250
rect 42150 32180 42160 32240
rect 42220 32180 42230 32240
rect 42150 32170 42230 32180
rect 42090 29530 42150 29540
rect 42090 29460 42150 29470
rect 42180 29490 42210 32170
rect 42270 29600 42300 32590
rect 42330 32520 42410 32530
rect 42330 32460 42340 32520
rect 42400 32460 42410 32520
rect 42330 32450 42410 32460
rect 44010 32450 44020 32510
rect 44080 32450 44090 32510
rect 42270 29590 42330 29600
rect 42270 29520 42330 29530
rect 42360 29550 42390 32450
rect 43630 30130 43710 30140
rect 43630 30070 43640 30130
rect 43700 30070 43710 30130
rect 43630 30060 43710 30070
rect 43780 30060 43790 30120
rect 43850 30060 43860 30120
rect 42560 29990 42640 30000
rect 42560 29930 42570 29990
rect 42630 29930 42640 29990
rect 42560 29920 42640 29930
rect 42360 29520 42530 29550
rect 42180 29460 42410 29490
rect 42000 29400 42290 29430
rect 41820 29340 42170 29370
rect 41640 29280 42050 29310
rect 41460 29220 41930 29250
rect 41280 29160 41810 29190
rect 39620 27360 39650 29160
rect 41780 27360 41810 29160
rect 41900 27360 41930 29220
rect 42020 27360 42050 29280
rect 42140 27360 42170 29340
rect 42260 27360 42290 29400
rect 42380 27360 42410 29460
rect 42500 27360 42530 29520
rect 42560 29140 42630 29920
rect 43640 29150 43710 30060
rect 43830 29150 43860 30060
rect 44030 29550 44060 32450
rect 44120 29600 44150 32590
rect 47260 32600 47270 32660
rect 47330 32600 47340 32660
rect 52250 32660 52330 32670
rect 47260 32590 47340 32600
rect 49060 32590 49070 32650
rect 49130 32590 49140 32650
rect 47080 32380 47160 32390
rect 44250 32310 44260 32370
rect 44320 32310 44330 32370
rect 44190 32170 44200 32230
rect 44260 32170 44270 32230
rect 43630 29140 43710 29150
rect 42560 29080 42570 29140
rect 42630 29080 42640 29140
rect 42560 29070 42640 29080
rect 43630 29080 43640 29140
rect 43700 29080 43710 29140
rect 43630 29060 43710 29080
rect 43800 29140 43860 29150
rect 43800 29070 43860 29080
rect 43890 29520 44060 29550
rect 44090 29590 44150 29600
rect 44090 29520 44150 29530
rect 43630 29000 43640 29060
rect 43700 29000 43710 29060
rect 43630 28990 43710 29000
rect 42560 28950 42640 28960
rect 42560 28890 42570 28950
rect 42630 28890 42640 28950
rect 42560 28880 42640 28890
rect 43090 28480 43710 28490
rect 43090 28420 43100 28480
rect 43160 28460 43710 28480
rect 43160 28420 43170 28460
rect 42670 28410 42750 28420
rect 43090 28410 43170 28420
rect 43510 28410 43590 28420
rect 42670 28390 42680 28410
rect 42560 28360 42680 28390
rect 42670 28350 42680 28360
rect 42740 28350 42750 28410
rect 42670 28340 42750 28350
rect 43510 28350 43520 28410
rect 43580 28390 43590 28410
rect 43580 28360 43710 28390
rect 43580 28350 43590 28360
rect 43510 28340 43590 28350
rect 43080 28310 43180 28330
rect 43080 28240 43100 28310
rect 43170 28240 43180 28310
rect 43080 28200 43180 28240
rect 43080 28130 43100 28200
rect 43170 28130 43180 28200
rect 43080 28120 43180 28130
rect 42670 28100 42750 28110
rect 42670 28080 42680 28100
rect 42560 28050 42680 28080
rect 42670 28040 42680 28050
rect 42740 28040 42750 28100
rect 43510 28100 43590 28110
rect 43510 28040 43520 28100
rect 43580 28080 43590 28100
rect 43580 28050 43710 28080
rect 43580 28040 43590 28050
rect 42670 28030 42750 28040
rect 43090 28030 43170 28040
rect 43510 28030 43590 28040
rect 43090 27970 43100 28030
rect 43160 27990 43170 28030
rect 43160 27970 43710 27990
rect 43090 27960 43710 27970
rect 43700 27420 43710 27440
rect 43890 27360 43920 29520
rect 44210 29490 44240 32170
rect 44300 29540 44330 32310
rect 47080 32320 47090 32380
rect 47150 32320 47160 32380
rect 47080 32310 47160 32320
rect 46900 32100 46980 32110
rect 44430 32030 44440 32090
rect 44500 32030 44510 32090
rect 44370 31890 44380 31950
rect 44440 31890 44450 31950
rect 44010 29460 44240 29490
rect 44270 29530 44330 29540
rect 44270 29460 44330 29470
rect 44010 27360 44040 29460
rect 44390 29430 44420 31890
rect 44480 29480 44510 32030
rect 46900 32040 46910 32100
rect 46970 32040 46980 32100
rect 46900 32030 46980 32040
rect 46720 31820 46800 31830
rect 44610 31750 44620 31810
rect 44680 31750 44690 31810
rect 44550 31610 44560 31670
rect 44620 31610 44630 31670
rect 44130 29400 44420 29430
rect 44450 29470 44510 29480
rect 44450 29400 44510 29410
rect 44130 27360 44160 29400
rect 44570 29370 44600 31610
rect 44660 29420 44690 31750
rect 46720 31760 46730 31820
rect 46790 31760 46800 31820
rect 46720 31750 46800 31760
rect 46360 31540 46440 31550
rect 44790 31470 44800 31530
rect 44860 31470 44870 31530
rect 44730 31330 44740 31390
rect 44800 31330 44810 31390
rect 44250 29340 44600 29370
rect 44630 29410 44690 29420
rect 44630 29340 44690 29350
rect 44250 27360 44280 29340
rect 44750 29310 44780 31330
rect 44840 29360 44870 31470
rect 46360 31480 46370 31540
rect 46430 31480 46440 31540
rect 46360 31470 46440 31480
rect 45150 30910 45160 30970
rect 45220 30910 45230 30970
rect 45090 30770 45100 30830
rect 45160 30770 45170 30830
rect 45000 30630 45010 30690
rect 45070 30630 45080 30690
rect 44910 30490 44920 30550
rect 44980 30490 44990 30550
rect 44370 29280 44780 29310
rect 44810 29350 44870 29360
rect 44810 29280 44870 29290
rect 44370 27330 44400 29280
rect 44930 29250 44960 30490
rect 45020 29300 45050 30630
rect 44490 29220 44960 29250
rect 44990 29290 45050 29300
rect 44990 29220 45050 29230
rect 44490 27360 44520 29220
rect 45110 29190 45140 30770
rect 45200 29240 45230 30910
rect 44610 29160 45140 29190
rect 45170 29230 45230 29240
rect 46360 29300 46390 31470
rect 46420 31400 46500 31410
rect 46420 31340 46430 31400
rect 46490 31340 46500 31400
rect 46420 31330 46500 31340
rect 46360 29290 46420 29300
rect 46360 29220 46420 29230
rect 46450 29250 46480 31330
rect 46540 31260 46620 31270
rect 46540 31200 46550 31260
rect 46610 31200 46620 31260
rect 46540 31190 46620 31200
rect 46540 29360 46570 31190
rect 46600 31120 46680 31130
rect 46600 31060 46610 31120
rect 46670 31060 46680 31120
rect 46600 31050 46680 31060
rect 46540 29350 46600 29360
rect 46540 29280 46600 29290
rect 46630 29310 46660 31050
rect 46720 29420 46750 31750
rect 46780 31680 46860 31690
rect 46780 31620 46790 31680
rect 46850 31620 46860 31680
rect 46780 31610 46860 31620
rect 46720 29410 46780 29420
rect 46720 29340 46780 29350
rect 46810 29370 46840 31610
rect 46900 29480 46930 32030
rect 46960 31960 47040 31970
rect 46960 31900 46970 31960
rect 47030 31900 47040 31960
rect 46960 31890 47040 31900
rect 46900 29470 46960 29480
rect 46900 29400 46960 29410
rect 46990 29430 47020 31890
rect 47080 29540 47110 32310
rect 47140 32240 47220 32250
rect 47140 32180 47150 32240
rect 47210 32180 47220 32240
rect 47140 32170 47220 32180
rect 47080 29530 47140 29540
rect 47080 29460 47140 29470
rect 47170 29490 47200 32170
rect 47260 29600 47290 32590
rect 47320 32520 47400 32530
rect 47320 32460 47330 32520
rect 47390 32460 47400 32520
rect 47320 32450 47400 32460
rect 49000 32450 49010 32510
rect 49070 32450 49080 32510
rect 47260 29590 47320 29600
rect 47260 29520 47320 29530
rect 47350 29550 47380 32450
rect 48620 30130 48700 30140
rect 48620 30070 48630 30130
rect 48690 30070 48700 30130
rect 48620 30060 48700 30070
rect 48770 30060 48780 30120
rect 48840 30060 48850 30120
rect 47550 29990 47630 30000
rect 47550 29930 47560 29990
rect 47620 29930 47630 29990
rect 47550 29920 47630 29930
rect 47350 29520 47520 29550
rect 47170 29460 47400 29490
rect 46990 29400 47280 29430
rect 46810 29340 47160 29370
rect 46630 29280 47040 29310
rect 46450 29220 46920 29250
rect 45170 29160 45230 29170
rect 44610 27360 44640 29160
rect 46770 27360 46800 29070
rect 46890 27360 46920 29220
rect 47010 27360 47040 29280
rect 47130 27360 47160 29340
rect 47250 27360 47280 29400
rect 47370 27360 47400 29460
rect 47490 27360 47520 29520
rect 47550 29140 47620 29920
rect 48630 29150 48700 30060
rect 48820 29150 48850 30060
rect 49020 29550 49050 32450
rect 49110 29600 49140 32590
rect 52250 32600 52260 32660
rect 52320 32600 52330 32660
rect 57240 32660 57320 32670
rect 52250 32590 52330 32600
rect 54050 32590 54060 32650
rect 54120 32590 54130 32650
rect 52070 32380 52150 32390
rect 49240 32310 49250 32370
rect 49310 32310 49320 32370
rect 49180 32170 49190 32230
rect 49250 32170 49260 32230
rect 48620 29140 48700 29150
rect 47550 29080 47560 29140
rect 47620 29080 47630 29140
rect 47550 29070 47630 29080
rect 48620 29080 48630 29140
rect 48690 29080 48700 29140
rect 48620 29060 48700 29080
rect 48790 29140 48850 29150
rect 48790 29070 48850 29080
rect 48880 29520 49050 29550
rect 49080 29590 49140 29600
rect 49080 29520 49140 29530
rect 48620 29000 48630 29060
rect 48690 29000 48700 29060
rect 48620 28990 48700 29000
rect 47550 28950 47630 28960
rect 47550 28890 47560 28950
rect 47620 28890 47630 28950
rect 47550 28880 47630 28890
rect 48080 28480 48700 28490
rect 48080 28420 48090 28480
rect 48150 28460 48700 28480
rect 48150 28420 48160 28460
rect 47660 28410 47740 28420
rect 48080 28410 48160 28420
rect 48500 28410 48580 28420
rect 47660 28390 47670 28410
rect 47550 28360 47670 28390
rect 47660 28350 47670 28360
rect 47730 28350 47740 28410
rect 47660 28340 47740 28350
rect 48500 28350 48510 28410
rect 48570 28390 48580 28410
rect 48570 28360 48700 28390
rect 48570 28350 48580 28360
rect 48500 28340 48580 28350
rect 48070 28310 48170 28330
rect 48070 28240 48090 28310
rect 48160 28240 48170 28310
rect 48070 28200 48170 28240
rect 48070 28130 48090 28200
rect 48160 28130 48170 28200
rect 48070 28120 48170 28130
rect 47660 28100 47740 28110
rect 47660 28080 47670 28100
rect 47550 28050 47670 28080
rect 47660 28040 47670 28050
rect 47730 28040 47740 28100
rect 48500 28100 48580 28110
rect 48500 28040 48510 28100
rect 48570 28080 48580 28100
rect 48570 28050 48700 28080
rect 48570 28040 48580 28050
rect 47660 28030 47740 28040
rect 48080 28030 48160 28040
rect 48500 28030 48580 28040
rect 48080 27970 48090 28030
rect 48150 27990 48160 28030
rect 48150 27970 48700 27990
rect 48080 27960 48700 27970
rect 48690 27420 48700 27440
rect 48880 27360 48910 29520
rect 49200 29490 49230 32170
rect 49290 29540 49320 32310
rect 52070 32320 52080 32380
rect 52140 32320 52150 32380
rect 52070 32310 52150 32320
rect 51710 32100 51790 32110
rect 49420 32030 49430 32090
rect 49490 32030 49500 32090
rect 49360 31890 49370 31950
rect 49430 31890 49440 31950
rect 49000 29460 49230 29490
rect 49260 29530 49320 29540
rect 49260 29460 49320 29470
rect 49000 27360 49030 29460
rect 49380 29430 49410 31890
rect 49470 29480 49500 32030
rect 51710 32040 51720 32100
rect 51780 32040 51790 32100
rect 51710 32030 51790 32040
rect 49600 31750 49610 31810
rect 49670 31750 49680 31810
rect 49540 31610 49550 31670
rect 49610 31610 49620 31670
rect 49120 29400 49410 29430
rect 49440 29470 49500 29480
rect 49440 29400 49500 29410
rect 49120 27360 49150 29400
rect 49560 29370 49590 31610
rect 49650 29420 49680 31750
rect 49960 31470 49970 31530
rect 50030 31470 50040 31530
rect 49900 31330 49910 31390
rect 49970 31330 49980 31390
rect 49780 31190 49790 31250
rect 49850 31190 49860 31250
rect 49720 31050 49730 31110
rect 49790 31050 49800 31110
rect 49240 29340 49590 29370
rect 49620 29410 49680 29420
rect 49620 29340 49680 29350
rect 49240 27360 49270 29340
rect 49740 29310 49770 31050
rect 49830 29360 49860 31190
rect 49360 29280 49770 29310
rect 49800 29350 49860 29360
rect 49800 29280 49860 29290
rect 49360 27360 49390 29280
rect 49920 29250 49950 31330
rect 50010 29300 50040 31470
rect 51710 29420 51740 32030
rect 51770 31960 51850 31970
rect 51770 31900 51780 31960
rect 51840 31900 51850 31960
rect 51770 31890 51850 31900
rect 51710 29410 51770 29420
rect 51710 29340 51770 29350
rect 51800 29370 51830 31890
rect 51890 31820 51970 31830
rect 51890 31760 51900 31820
rect 51960 31760 51970 31820
rect 51890 31750 51970 31760
rect 51890 29480 51920 31750
rect 51950 31680 52030 31690
rect 51950 31620 51960 31680
rect 52020 31620 52030 31680
rect 51950 31610 52030 31620
rect 51890 29470 51950 29480
rect 51890 29400 51950 29410
rect 51980 29430 52010 31610
rect 52070 29540 52100 32310
rect 52130 32240 52210 32250
rect 52130 32180 52140 32240
rect 52200 32180 52210 32240
rect 52130 32170 52210 32180
rect 52070 29530 52130 29540
rect 52070 29460 52130 29470
rect 52160 29490 52190 32170
rect 52250 29600 52280 32590
rect 52310 32520 52390 32530
rect 52310 32460 52320 32520
rect 52380 32460 52390 32520
rect 52310 32450 52390 32460
rect 53990 32450 54000 32510
rect 54060 32450 54070 32510
rect 52250 29590 52310 29600
rect 52250 29520 52310 29530
rect 52340 29550 52370 32450
rect 53610 30130 53690 30140
rect 53610 30070 53620 30130
rect 53680 30070 53690 30130
rect 53610 30060 53690 30070
rect 53760 30060 53770 30120
rect 53830 30060 53840 30120
rect 52540 29990 52620 30000
rect 52540 29930 52550 29990
rect 52610 29930 52620 29990
rect 52540 29920 52620 29930
rect 52340 29520 52510 29550
rect 52160 29460 52390 29490
rect 51980 29400 52270 29430
rect 51800 29340 52150 29370
rect 49480 29220 49950 29250
rect 49980 29290 50040 29300
rect 49980 29220 50040 29230
rect 49480 27360 49510 29220
rect 49600 27360 49630 29070
rect 51760 27360 51790 29070
rect 51880 27360 51910 29070
rect 52000 27360 52030 29070
rect 52120 27360 52150 29340
rect 52240 27360 52270 29400
rect 52360 27360 52390 29460
rect 52480 27360 52510 29520
rect 52540 29140 52610 29920
rect 53620 29150 53690 30060
rect 53810 29150 53840 30060
rect 54010 29550 54040 32450
rect 54100 29600 54130 32590
rect 57240 32600 57250 32660
rect 57310 32600 57320 32660
rect 62230 32660 62310 32670
rect 57240 32590 57320 32600
rect 59040 32590 59050 32650
rect 59110 32590 59120 32650
rect 57060 32380 57140 32390
rect 54230 32310 54240 32370
rect 54300 32310 54310 32370
rect 54170 32170 54180 32230
rect 54240 32170 54250 32230
rect 53610 29140 53690 29150
rect 52540 29080 52550 29140
rect 52610 29080 52620 29140
rect 52540 29070 52620 29080
rect 53610 29080 53620 29140
rect 53680 29080 53690 29140
rect 53610 29060 53690 29080
rect 53780 29140 53840 29150
rect 53780 29070 53840 29080
rect 53870 29520 54040 29550
rect 54070 29590 54130 29600
rect 54070 29520 54130 29530
rect 53610 29000 53620 29060
rect 53680 29000 53690 29060
rect 53610 28990 53690 29000
rect 52540 28950 52620 28960
rect 52540 28890 52550 28950
rect 52610 28890 52620 28950
rect 52540 28880 52620 28890
rect 53070 28480 53690 28490
rect 53070 28420 53080 28480
rect 53140 28460 53690 28480
rect 53140 28420 53150 28460
rect 52650 28410 52730 28420
rect 53070 28410 53150 28420
rect 53490 28410 53570 28420
rect 52650 28390 52660 28410
rect 52540 28360 52660 28390
rect 52650 28350 52660 28360
rect 52720 28350 52730 28410
rect 52650 28340 52730 28350
rect 53490 28350 53500 28410
rect 53560 28390 53570 28410
rect 53560 28360 53690 28390
rect 53560 28350 53570 28360
rect 53490 28340 53570 28350
rect 53060 28310 53160 28330
rect 53060 28240 53080 28310
rect 53150 28240 53160 28310
rect 53060 28200 53160 28240
rect 53060 28130 53080 28200
rect 53150 28130 53160 28200
rect 53060 28120 53160 28130
rect 52650 28100 52730 28110
rect 52650 28080 52660 28100
rect 52540 28050 52660 28080
rect 52650 28040 52660 28050
rect 52720 28040 52730 28100
rect 53490 28100 53570 28110
rect 53490 28040 53500 28100
rect 53560 28080 53570 28100
rect 53560 28050 53690 28080
rect 53560 28040 53570 28050
rect 52650 28030 52730 28040
rect 53070 28030 53150 28040
rect 53490 28030 53570 28040
rect 53070 27970 53080 28030
rect 53140 27990 53150 28030
rect 53140 27970 53690 27990
rect 53070 27960 53690 27970
rect 53680 27420 53690 27440
rect 53870 27360 53900 29520
rect 54190 29490 54220 32170
rect 54280 29540 54310 32310
rect 57060 32320 57070 32380
rect 57130 32320 57140 32380
rect 57060 32310 57140 32320
rect 56700 32100 56780 32110
rect 54590 32030 54600 32090
rect 54660 32030 54670 32090
rect 54530 31890 54540 31950
rect 54600 31890 54610 31950
rect 54410 31750 54420 31810
rect 54480 31750 54490 31810
rect 54350 31610 54360 31670
rect 54420 31610 54430 31670
rect 53990 29460 54220 29490
rect 54250 29530 54310 29540
rect 54250 29460 54310 29470
rect 53990 27360 54020 29460
rect 54370 29430 54400 31610
rect 54460 29480 54490 31750
rect 54110 29400 54400 29430
rect 54430 29470 54490 29480
rect 54430 29400 54490 29410
rect 54110 27360 54140 29400
rect 54550 29370 54580 31890
rect 54640 29420 54670 32030
rect 54230 29340 54580 29370
rect 54610 29410 54670 29420
rect 54610 29340 54670 29350
rect 56700 32040 56710 32100
rect 56770 32040 56780 32100
rect 56700 32030 56780 32040
rect 56700 29420 56730 32030
rect 56760 31960 56840 31970
rect 56760 31900 56770 31960
rect 56830 31900 56840 31960
rect 56760 31890 56840 31900
rect 56700 29410 56760 29420
rect 56700 29340 56760 29350
rect 56790 29370 56820 31890
rect 56880 31820 56960 31830
rect 56880 31760 56890 31820
rect 56950 31760 56960 31820
rect 56880 31750 56960 31760
rect 56880 29480 56910 31750
rect 56940 31680 57020 31690
rect 56940 31620 56950 31680
rect 57010 31620 57020 31680
rect 56940 31610 57020 31620
rect 56880 29470 56940 29480
rect 56880 29400 56940 29410
rect 56970 29430 57000 31610
rect 57060 29540 57090 32310
rect 57120 32240 57200 32250
rect 57120 32180 57130 32240
rect 57190 32180 57200 32240
rect 57120 32170 57200 32180
rect 57060 29530 57120 29540
rect 57060 29460 57120 29470
rect 57150 29490 57180 32170
rect 57240 29600 57270 32590
rect 57300 32520 57380 32530
rect 57300 32460 57310 32520
rect 57370 32460 57380 32520
rect 57300 32450 57380 32460
rect 58980 32450 58990 32510
rect 59050 32450 59060 32510
rect 57240 29590 57300 29600
rect 57240 29520 57300 29530
rect 57330 29550 57360 32450
rect 58600 30130 58680 30140
rect 58600 30070 58610 30130
rect 58670 30070 58680 30130
rect 58600 30060 58680 30070
rect 58750 30060 58760 30120
rect 58820 30060 58830 30120
rect 57530 29990 57610 30000
rect 57530 29930 57540 29990
rect 57600 29930 57610 29990
rect 57530 29920 57610 29930
rect 57330 29520 57500 29550
rect 57150 29460 57380 29490
rect 56970 29400 57260 29430
rect 56790 29340 57140 29370
rect 54230 27360 54260 29340
rect 54350 27360 54380 29070
rect 54470 27360 54500 29070
rect 54590 27360 54620 29070
rect 56750 27360 56780 29070
rect 56870 27360 56900 29070
rect 56990 27360 57020 29070
rect 57110 27360 57140 29340
rect 57230 27360 57260 29400
rect 57350 27360 57380 29460
rect 57470 27360 57500 29520
rect 57530 29140 57600 29920
rect 58610 29150 58680 30060
rect 58800 29150 58830 30060
rect 59000 29550 59030 32450
rect 59090 29600 59120 32590
rect 62230 32600 62240 32660
rect 62300 32600 62310 32660
rect 67220 32660 67300 32670
rect 62230 32590 62310 32600
rect 64030 32590 64040 32650
rect 64100 32590 64110 32650
rect 62050 32380 62130 32390
rect 59220 32310 59230 32370
rect 59290 32310 59300 32370
rect 59160 32170 59170 32230
rect 59230 32170 59240 32230
rect 58600 29140 58680 29150
rect 57530 29080 57540 29140
rect 57600 29080 57610 29140
rect 57530 29070 57610 29080
rect 58600 29080 58610 29140
rect 58670 29080 58680 29140
rect 58600 29060 58680 29080
rect 58770 29140 58830 29150
rect 58770 29070 58830 29080
rect 58860 29520 59030 29550
rect 59060 29590 59120 29600
rect 59060 29520 59120 29530
rect 58600 29000 58610 29060
rect 58670 29000 58680 29060
rect 58600 28990 58680 29000
rect 57530 28950 57610 28960
rect 57530 28890 57540 28950
rect 57600 28890 57610 28950
rect 57530 28880 57610 28890
rect 58060 28480 58680 28490
rect 58060 28420 58070 28480
rect 58130 28460 58680 28480
rect 58130 28420 58140 28460
rect 57640 28410 57720 28420
rect 58060 28410 58140 28420
rect 58480 28410 58560 28420
rect 57640 28390 57650 28410
rect 57530 28360 57650 28390
rect 57640 28350 57650 28360
rect 57710 28350 57720 28410
rect 57640 28340 57720 28350
rect 58480 28350 58490 28410
rect 58550 28390 58560 28410
rect 58550 28360 58680 28390
rect 58550 28350 58560 28360
rect 58480 28340 58560 28350
rect 58050 28310 58150 28330
rect 58050 28240 58070 28310
rect 58140 28240 58150 28310
rect 58050 28200 58150 28240
rect 58050 28130 58070 28200
rect 58140 28130 58150 28200
rect 58050 28120 58150 28130
rect 57640 28100 57720 28110
rect 57640 28080 57650 28100
rect 57530 28050 57650 28080
rect 57640 28040 57650 28050
rect 57710 28040 57720 28100
rect 58480 28100 58560 28110
rect 58480 28040 58490 28100
rect 58550 28080 58560 28100
rect 58550 28050 58680 28080
rect 58550 28040 58560 28050
rect 57640 28030 57720 28040
rect 58060 28030 58140 28040
rect 58480 28030 58560 28040
rect 58060 27970 58070 28030
rect 58130 27990 58140 28030
rect 58130 27970 58680 27990
rect 58060 27960 58680 27970
rect 58670 27420 58680 27440
rect 58860 27360 58890 29520
rect 59180 29490 59210 32170
rect 59270 29540 59300 32310
rect 62050 32320 62060 32380
rect 62120 32320 62130 32380
rect 62050 32310 62130 32320
rect 59580 32030 59590 32090
rect 59650 32030 59660 32090
rect 59520 31890 59530 31950
rect 59590 31890 59600 31950
rect 59400 31750 59410 31810
rect 59470 31750 59480 31810
rect 59340 31610 59350 31670
rect 59410 31610 59420 31670
rect 58980 29460 59210 29490
rect 59240 29530 59300 29540
rect 59240 29460 59300 29470
rect 58980 27360 59010 29460
rect 59360 29430 59390 31610
rect 59450 29480 59480 31750
rect 59100 29400 59390 29430
rect 59420 29470 59480 29480
rect 59420 29400 59480 29410
rect 59100 27360 59130 29400
rect 59540 29370 59570 31890
rect 59630 29420 59660 32030
rect 62050 29540 62080 32310
rect 62110 32240 62190 32250
rect 62110 32180 62120 32240
rect 62180 32180 62190 32240
rect 62110 32170 62190 32180
rect 62050 29530 62110 29540
rect 62050 29460 62110 29470
rect 62140 29490 62170 32170
rect 62230 29600 62260 32590
rect 62290 32520 62370 32530
rect 62290 32460 62300 32520
rect 62360 32460 62370 32520
rect 62290 32450 62370 32460
rect 63970 32450 63980 32510
rect 64040 32450 64050 32510
rect 62230 29590 62290 29600
rect 62230 29520 62290 29530
rect 62320 29550 62350 32450
rect 63590 30130 63670 30140
rect 63590 30070 63600 30130
rect 63660 30070 63670 30130
rect 63590 30060 63670 30070
rect 63740 30060 63750 30120
rect 63810 30060 63820 30120
rect 62520 29990 62600 30000
rect 62520 29930 62530 29990
rect 62590 29930 62600 29990
rect 62520 29920 62600 29930
rect 62320 29520 62490 29550
rect 62140 29460 62370 29490
rect 59220 29340 59570 29370
rect 59600 29410 59660 29420
rect 59600 29340 59660 29350
rect 59220 27360 59250 29340
rect 59340 27360 59370 29070
rect 59460 27360 59490 29070
rect 59580 27360 59610 29070
rect 61740 27360 61770 29070
rect 61860 27360 61890 29070
rect 61980 27360 62010 29070
rect 62100 27360 62130 29070
rect 62220 27360 62250 29070
rect 62340 27360 62370 29460
rect 62460 27360 62490 29520
rect 62520 29140 62590 29920
rect 63600 29150 63670 30060
rect 63790 29150 63820 30060
rect 63990 29550 64020 32450
rect 64080 29600 64110 32590
rect 67220 32600 67230 32660
rect 67290 32600 67300 32660
rect 72210 32660 72290 32670
rect 67220 32590 67300 32600
rect 69020 32590 69030 32650
rect 69090 32590 69100 32650
rect 67040 32380 67120 32390
rect 64210 32310 64220 32370
rect 64280 32310 64290 32370
rect 64150 32170 64160 32230
rect 64220 32170 64230 32230
rect 63590 29140 63670 29150
rect 62520 29080 62530 29140
rect 62590 29080 62600 29140
rect 62520 29070 62600 29080
rect 63590 29080 63600 29140
rect 63660 29080 63670 29140
rect 63590 29060 63670 29080
rect 63760 29140 63820 29150
rect 63760 29070 63820 29080
rect 63850 29520 64020 29550
rect 64050 29590 64110 29600
rect 64050 29520 64110 29530
rect 63590 29000 63600 29060
rect 63660 29000 63670 29060
rect 63590 28990 63670 29000
rect 62520 28950 62600 28960
rect 62520 28890 62530 28950
rect 62590 28890 62600 28950
rect 62520 28880 62600 28890
rect 63050 28480 63670 28490
rect 63050 28420 63060 28480
rect 63120 28460 63670 28480
rect 63120 28420 63130 28460
rect 62630 28410 62710 28420
rect 63050 28410 63130 28420
rect 63470 28410 63550 28420
rect 62630 28390 62640 28410
rect 62520 28360 62640 28390
rect 62630 28350 62640 28360
rect 62700 28350 62710 28410
rect 62630 28340 62710 28350
rect 63470 28350 63480 28410
rect 63540 28390 63550 28410
rect 63540 28360 63670 28390
rect 63540 28350 63550 28360
rect 63470 28340 63550 28350
rect 63040 28310 63140 28330
rect 63040 28240 63060 28310
rect 63130 28240 63140 28310
rect 63040 28200 63140 28240
rect 63040 28130 63060 28200
rect 63130 28130 63140 28200
rect 63040 28120 63140 28130
rect 62630 28100 62710 28110
rect 62630 28080 62640 28100
rect 62520 28050 62640 28080
rect 62630 28040 62640 28050
rect 62700 28040 62710 28100
rect 63470 28100 63550 28110
rect 63470 28040 63480 28100
rect 63540 28080 63550 28100
rect 63540 28050 63670 28080
rect 63540 28040 63550 28050
rect 62630 28030 62710 28040
rect 63050 28030 63130 28040
rect 63470 28030 63550 28040
rect 63050 27970 63060 28030
rect 63120 27990 63130 28030
rect 63120 27970 63670 27990
rect 63050 27960 63670 27970
rect 63660 27420 63670 27440
rect 63850 27360 63880 29520
rect 64170 29490 64200 32170
rect 64260 29540 64290 32310
rect 63970 29460 64200 29490
rect 64230 29530 64290 29540
rect 64230 29460 64290 29470
rect 67040 32320 67050 32380
rect 67110 32320 67120 32380
rect 67040 32310 67120 32320
rect 67040 29540 67070 32310
rect 67100 32240 67180 32250
rect 67100 32180 67110 32240
rect 67170 32180 67180 32240
rect 67100 32170 67180 32180
rect 67040 29530 67100 29540
rect 67040 29460 67100 29470
rect 67130 29490 67160 32170
rect 67220 29600 67250 32590
rect 67280 32520 67360 32530
rect 67280 32460 67290 32520
rect 67350 32460 67360 32520
rect 67280 32450 67360 32460
rect 68960 32450 68970 32510
rect 69030 32450 69040 32510
rect 67220 29590 67280 29600
rect 67220 29520 67280 29530
rect 67310 29550 67340 32450
rect 68580 30130 68660 30140
rect 68580 30070 68590 30130
rect 68650 30070 68660 30130
rect 68580 30060 68660 30070
rect 68730 30060 68740 30120
rect 68800 30060 68810 30120
rect 67510 29990 67590 30000
rect 67510 29930 67520 29990
rect 67580 29930 67590 29990
rect 67510 29920 67590 29930
rect 67310 29520 67480 29550
rect 67130 29460 67360 29490
rect 63970 27360 64000 29460
rect 64090 27360 64120 29070
rect 64210 27360 64240 29070
rect 64330 27360 64360 29070
rect 64450 27360 64480 29070
rect 64570 27360 64600 29070
rect 66730 27360 66760 29070
rect 66850 27360 66880 29070
rect 66970 27360 67000 29070
rect 67090 27360 67120 29070
rect 67210 27360 67240 29070
rect 67330 27360 67360 29460
rect 67450 27360 67480 29520
rect 67510 29140 67580 29920
rect 68590 29150 68660 30060
rect 68780 29150 68810 30060
rect 68980 29550 69010 32450
rect 69070 29600 69100 32590
rect 72210 32600 72220 32660
rect 72280 32600 72290 32660
rect 77200 32660 77280 32670
rect 72210 32590 72290 32600
rect 74010 32590 74020 32650
rect 74080 32590 74090 32650
rect 69200 32310 69210 32370
rect 69270 32310 69280 32370
rect 69140 32170 69150 32230
rect 69210 32170 69220 32230
rect 68580 29140 68660 29150
rect 67510 29080 67520 29140
rect 67580 29080 67590 29140
rect 67510 29070 67590 29080
rect 68580 29080 68590 29140
rect 68650 29080 68660 29140
rect 68580 29060 68660 29080
rect 68750 29140 68810 29150
rect 68750 29070 68810 29080
rect 68840 29520 69010 29550
rect 69040 29590 69100 29600
rect 69040 29520 69100 29530
rect 68580 29000 68590 29060
rect 68650 29000 68660 29060
rect 68580 28990 68660 29000
rect 67510 28950 67590 28960
rect 67510 28890 67520 28950
rect 67580 28890 67590 28950
rect 67510 28880 67590 28890
rect 68040 28480 68660 28490
rect 68040 28420 68050 28480
rect 68110 28460 68660 28480
rect 68110 28420 68120 28460
rect 67620 28410 67700 28420
rect 68040 28410 68120 28420
rect 68460 28410 68540 28420
rect 67620 28390 67630 28410
rect 67510 28360 67630 28390
rect 67620 28350 67630 28360
rect 67690 28350 67700 28410
rect 67620 28340 67700 28350
rect 68460 28350 68470 28410
rect 68530 28390 68540 28410
rect 68530 28360 68660 28390
rect 68530 28350 68540 28360
rect 68460 28340 68540 28350
rect 68030 28310 68130 28330
rect 68030 28240 68050 28310
rect 68120 28240 68130 28310
rect 68030 28200 68130 28240
rect 68030 28130 68050 28200
rect 68120 28130 68130 28200
rect 68030 28120 68130 28130
rect 67620 28100 67700 28110
rect 67620 28080 67630 28100
rect 67510 28050 67630 28080
rect 67620 28040 67630 28050
rect 67690 28040 67700 28100
rect 68460 28100 68540 28110
rect 68460 28040 68470 28100
rect 68530 28080 68540 28100
rect 68530 28050 68660 28080
rect 68530 28040 68540 28050
rect 67620 28030 67700 28040
rect 68040 28030 68120 28040
rect 68460 28030 68540 28040
rect 68040 27970 68050 28030
rect 68110 27990 68120 28030
rect 68110 27970 68660 27990
rect 68040 27960 68660 27970
rect 68650 27420 68660 27440
rect 68840 27360 68870 29520
rect 69160 29490 69190 32170
rect 69250 29540 69280 32310
rect 68960 29460 69190 29490
rect 69220 29530 69280 29540
rect 72210 29600 72240 32590
rect 72270 32520 72350 32530
rect 72270 32460 72280 32520
rect 72340 32460 72350 32520
rect 72270 32450 72350 32460
rect 73950 32450 73960 32510
rect 74020 32450 74030 32510
rect 72210 29590 72270 29600
rect 72210 29520 72270 29530
rect 72300 29550 72330 32450
rect 73570 30130 73650 30140
rect 73570 30070 73580 30130
rect 73640 30070 73650 30130
rect 73570 30060 73650 30070
rect 73720 30060 73730 30120
rect 73790 30060 73800 30120
rect 72500 29990 72580 30000
rect 72500 29930 72510 29990
rect 72570 29930 72580 29990
rect 72500 29920 72580 29930
rect 72300 29520 72470 29550
rect 69220 29460 69280 29470
rect 68960 27360 68990 29460
rect 69080 27360 69110 29070
rect 69200 27360 69230 29070
rect 69320 27360 69350 29070
rect 69440 27360 69470 29070
rect 69560 27360 69590 29070
rect 71720 27360 71750 29070
rect 71840 27360 71870 29070
rect 71960 27360 71990 29070
rect 72080 27360 72110 29070
rect 72200 27360 72230 29070
rect 72320 27360 72350 29070
rect 72440 27360 72470 29520
rect 72500 29140 72570 29920
rect 73580 29150 73650 30060
rect 73770 29150 73800 30060
rect 73970 29550 74000 32450
rect 74060 29600 74090 32590
rect 73570 29140 73650 29150
rect 72500 29080 72510 29140
rect 72570 29080 72580 29140
rect 72500 29070 72580 29080
rect 73570 29080 73580 29140
rect 73640 29080 73650 29140
rect 73570 29060 73650 29080
rect 73740 29140 73800 29150
rect 73740 29070 73800 29080
rect 73830 29520 74000 29550
rect 74030 29590 74090 29600
rect 74030 29520 74090 29530
rect 77200 32600 77210 32660
rect 77270 32600 77280 32660
rect 77200 32590 77280 32600
rect 79000 32590 79010 32650
rect 79070 32590 79080 32650
rect 77200 29600 77230 32590
rect 77260 32520 77340 32530
rect 77260 32460 77270 32520
rect 77330 32460 77340 32520
rect 77260 32450 77340 32460
rect 78940 32450 78950 32510
rect 79010 32450 79020 32510
rect 77200 29590 77260 29600
rect 77200 29520 77260 29530
rect 77290 29550 77320 32450
rect 78560 30130 78640 30140
rect 78560 30070 78570 30130
rect 78630 30070 78640 30130
rect 78560 30060 78640 30070
rect 78710 30060 78720 30120
rect 78780 30060 78790 30120
rect 77490 29990 77570 30000
rect 77490 29930 77500 29990
rect 77560 29930 77570 29990
rect 77490 29920 77570 29930
rect 77290 29520 77460 29550
rect 73570 29000 73580 29060
rect 73640 29000 73650 29060
rect 73570 28990 73650 29000
rect 72500 28950 72580 28960
rect 72500 28890 72510 28950
rect 72570 28890 72580 28950
rect 72500 28880 72580 28890
rect 73030 28480 73650 28490
rect 73030 28420 73040 28480
rect 73100 28460 73650 28480
rect 73100 28420 73110 28460
rect 72610 28410 72690 28420
rect 73030 28410 73110 28420
rect 73450 28410 73530 28420
rect 72610 28390 72620 28410
rect 72500 28360 72620 28390
rect 72610 28350 72620 28360
rect 72680 28350 72690 28410
rect 72610 28340 72690 28350
rect 73450 28350 73460 28410
rect 73520 28390 73530 28410
rect 73520 28360 73650 28390
rect 73520 28350 73530 28360
rect 73450 28340 73530 28350
rect 73020 28310 73120 28330
rect 73020 28240 73040 28310
rect 73110 28240 73120 28310
rect 73020 28200 73120 28240
rect 73020 28130 73040 28200
rect 73110 28130 73120 28200
rect 73020 28120 73120 28130
rect 72610 28100 72690 28110
rect 72610 28080 72620 28100
rect 72500 28050 72620 28080
rect 72610 28040 72620 28050
rect 72680 28040 72690 28100
rect 73450 28100 73530 28110
rect 73450 28040 73460 28100
rect 73520 28080 73530 28100
rect 73520 28050 73650 28080
rect 73520 28040 73530 28050
rect 72610 28030 72690 28040
rect 73030 28030 73110 28040
rect 73450 28030 73530 28040
rect 73030 27970 73040 28030
rect 73100 27990 73110 28030
rect 73100 27970 73650 27990
rect 73030 27960 73650 27970
rect 73640 27420 73650 27440
rect 73830 27360 73860 29520
rect 73950 27360 73980 29070
rect 74070 27360 74100 29070
rect 74190 27360 74220 29070
rect 74310 27360 74340 29070
rect 74430 27360 74460 29070
rect 74550 27360 74580 29070
rect 76710 27360 76740 29070
rect 76830 27360 76860 29070
rect 76950 27360 76980 29070
rect 77070 27360 77100 29070
rect 77190 27360 77220 29070
rect 77310 27360 77340 29070
rect 77430 27360 77460 29520
rect 77490 29140 77560 29920
rect 78570 29150 78640 30060
rect 78760 29150 78790 30060
rect 78960 29550 78990 32450
rect 79050 29600 79080 32590
rect 78560 29140 78640 29150
rect 77490 29080 77500 29140
rect 77560 29080 77570 29140
rect 77490 29070 77570 29080
rect 78560 29080 78570 29140
rect 78630 29080 78640 29140
rect 78560 29060 78640 29080
rect 78730 29140 78790 29150
rect 78730 29070 78790 29080
rect 78820 29520 78990 29550
rect 79020 29590 79080 29600
rect 79020 29520 79080 29530
rect 82210 29990 82290 30000
rect 82210 29930 82220 29990
rect 82280 29930 82290 29990
rect 82210 29920 82290 29930
rect 78560 29000 78570 29060
rect 78630 29000 78640 29060
rect 78560 28990 78640 29000
rect 77490 28950 77570 28960
rect 77490 28890 77500 28950
rect 77560 28890 77570 28950
rect 77490 28880 77570 28890
rect 78020 28480 78640 28490
rect 78020 28420 78030 28480
rect 78090 28460 78640 28480
rect 78090 28420 78100 28460
rect 77600 28410 77680 28420
rect 78020 28410 78100 28420
rect 78440 28410 78520 28420
rect 77600 28390 77610 28410
rect 77490 28360 77610 28390
rect 77600 28350 77610 28360
rect 77670 28350 77680 28410
rect 77600 28340 77680 28350
rect 78440 28350 78450 28410
rect 78510 28390 78520 28410
rect 78510 28360 78640 28390
rect 78510 28350 78520 28360
rect 78440 28340 78520 28350
rect 78010 28310 78110 28330
rect 78010 28240 78030 28310
rect 78100 28240 78110 28310
rect 78010 28200 78110 28240
rect 78010 28130 78030 28200
rect 78100 28130 78110 28200
rect 78010 28120 78110 28130
rect 77600 28100 77680 28110
rect 77600 28080 77610 28100
rect 77490 28050 77610 28080
rect 77600 28040 77610 28050
rect 77670 28040 77680 28100
rect 78440 28100 78520 28110
rect 78440 28040 78450 28100
rect 78510 28080 78520 28100
rect 78510 28050 78640 28080
rect 78510 28040 78520 28050
rect 77600 28030 77680 28040
rect 78020 28030 78100 28040
rect 78440 28030 78520 28040
rect 78020 27970 78030 28030
rect 78090 27990 78100 28030
rect 78090 27970 78640 27990
rect 78020 27960 78640 27970
rect 78630 27420 78640 27440
rect 78820 27360 78850 29520
rect 82210 29140 82280 29920
rect 82210 29080 82220 29140
rect 82280 29080 82290 29140
rect 82210 29070 82290 29080
rect 78940 27360 78970 29070
rect 79060 27360 79090 29070
rect 79180 27360 79210 29070
rect 79300 27360 79330 29070
rect 79420 27360 79450 29070
rect 79540 27360 79570 29070
rect -2860 -1710 -2830 23940
rect -2740 -1710 -2710 23940
rect -2620 -1710 -2590 23940
rect -2500 -1710 -2470 23940
rect -2380 -1710 -2350 23940
rect -2260 -1710 -2230 23940
rect -2140 -1710 -2110 23940
rect -1010 23930 -930 23940
rect -1010 23870 -1000 23930
rect -940 23870 -930 23930
rect -1010 23860 -930 23870
rect -2080 23820 -2000 23830
rect -2080 23760 -2070 23820
rect -2010 23760 -2000 23820
rect -2080 23750 -2000 23760
rect -1550 23350 -930 23360
rect -1550 23290 -1540 23350
rect -1480 23330 -930 23350
rect -1480 23290 -1470 23330
rect -1970 23280 -1890 23290
rect -1550 23280 -1470 23290
rect -1130 23280 -1050 23290
rect -1970 23260 -1960 23280
rect -2080 23230 -1960 23260
rect -1970 23220 -1960 23230
rect -1900 23220 -1890 23280
rect -1970 23210 -1890 23220
rect -1130 23220 -1120 23280
rect -1060 23260 -1050 23280
rect -1060 23230 -930 23260
rect -1060 23220 -1050 23230
rect -1130 23210 -1050 23220
rect -1560 23180 -1460 23200
rect -1560 23110 -1540 23180
rect -1470 23110 -1460 23180
rect -1560 23070 -1460 23110
rect -1560 23000 -1540 23070
rect -1470 23000 -1460 23070
rect -1560 22990 -1460 23000
rect -1970 22970 -1890 22980
rect -1970 22950 -1960 22970
rect -2080 22920 -1960 22950
rect -1970 22910 -1960 22920
rect -1900 22910 -1890 22970
rect -1130 22970 -1050 22980
rect -1130 22910 -1120 22970
rect -1060 22950 -1050 22970
rect -1060 22920 -930 22950
rect -1060 22910 -1050 22920
rect -1970 22900 -1890 22910
rect -1550 22900 -1470 22910
rect -1130 22900 -1050 22910
rect -1550 22840 -1540 22900
rect -1480 22860 -1470 22900
rect -1480 22840 -930 22860
rect -1550 22830 -930 22840
rect -1020 22360 -930 22370
rect -1020 22300 -1010 22360
rect -940 22300 -930 22360
rect -1020 22290 -930 22300
rect -1010 22220 -930 22230
rect -1010 22160 -1000 22220
rect -940 22160 -930 22220
rect -1010 22150 -930 22160
rect -2080 22110 -2000 22120
rect -2080 22050 -2070 22110
rect -2010 22050 -2000 22110
rect -2080 22040 -2000 22050
rect -1550 21640 -930 21650
rect -1550 21580 -1540 21640
rect -1480 21620 -930 21640
rect -1480 21580 -1470 21620
rect -1970 21570 -1890 21580
rect -1550 21570 -1470 21580
rect -1130 21570 -1050 21580
rect -1970 21550 -1960 21570
rect -2080 21520 -1960 21550
rect -1970 21510 -1960 21520
rect -1900 21510 -1890 21570
rect -1970 21500 -1890 21510
rect -1130 21510 -1120 21570
rect -1060 21550 -1050 21570
rect -1060 21520 -930 21550
rect -1060 21510 -1050 21520
rect -1130 21500 -1050 21510
rect -1560 21470 -1460 21490
rect -1560 21400 -1540 21470
rect -1470 21400 -1460 21470
rect -1560 21360 -1460 21400
rect -1560 21290 -1540 21360
rect -1470 21290 -1460 21360
rect -1560 21280 -1460 21290
rect -1970 21260 -1890 21270
rect -1970 21240 -1960 21260
rect -2080 21210 -1960 21240
rect -1970 21200 -1960 21210
rect -1900 21200 -1890 21260
rect -1130 21260 -1050 21270
rect -1130 21200 -1120 21260
rect -1060 21240 -1050 21260
rect -1060 21210 -930 21240
rect -1060 21200 -1050 21210
rect -1970 21190 -1890 21200
rect -1550 21190 -1470 21200
rect -1130 21190 -1050 21200
rect -1550 21130 -1540 21190
rect -1480 21150 -1470 21190
rect -1480 21130 -930 21150
rect -1550 21120 -930 21130
rect -1020 20650 -930 20660
rect -1020 20590 -1010 20650
rect -940 20590 -930 20650
rect -1020 20580 -930 20590
rect -1010 20510 -930 20520
rect -1010 20450 -1000 20510
rect -940 20450 -930 20510
rect -1010 20440 -930 20450
rect -2080 20400 -2000 20410
rect -2080 20340 -2070 20400
rect -2010 20340 -2000 20400
rect -2080 20330 -2000 20340
rect -1550 19930 -930 19940
rect -1550 19870 -1540 19930
rect -1480 19910 -930 19930
rect -1480 19870 -1470 19910
rect -1970 19860 -1890 19870
rect -1550 19860 -1470 19870
rect -1130 19860 -1050 19870
rect -1970 19840 -1960 19860
rect -2080 19810 -1960 19840
rect -1970 19800 -1960 19810
rect -1900 19800 -1890 19860
rect -1970 19790 -1890 19800
rect -1130 19800 -1120 19860
rect -1060 19840 -1050 19860
rect -1060 19810 -930 19840
rect -1060 19800 -1050 19810
rect -1130 19790 -1050 19800
rect -1560 19760 -1460 19780
rect -1560 19690 -1540 19760
rect -1470 19690 -1460 19760
rect -1560 19650 -1460 19690
rect -1560 19580 -1540 19650
rect -1470 19580 -1460 19650
rect -1560 19570 -1460 19580
rect -1970 19550 -1890 19560
rect -1970 19530 -1960 19550
rect -2080 19500 -1960 19530
rect -1970 19490 -1960 19500
rect -1900 19490 -1890 19550
rect -1130 19550 -1050 19560
rect -1130 19490 -1120 19550
rect -1060 19530 -1050 19550
rect -1060 19500 -930 19530
rect -1060 19490 -1050 19500
rect -1970 19480 -1890 19490
rect -1550 19480 -1470 19490
rect -1130 19480 -1050 19490
rect -1550 19420 -1540 19480
rect -1480 19440 -1470 19480
rect -1480 19420 -930 19440
rect -1550 19410 -930 19420
rect -1020 18940 -930 18950
rect -1020 18880 -1010 18940
rect -940 18880 -930 18940
rect -1020 18870 -930 18880
rect -1010 18800 -930 18810
rect -1010 18740 -1000 18800
rect -940 18740 -930 18800
rect -1010 18730 -930 18740
rect -2080 18690 -2000 18700
rect -2080 18630 -2070 18690
rect -2010 18630 -2000 18690
rect -2080 18620 -2000 18630
rect -1550 18220 -930 18230
rect -1550 18160 -1540 18220
rect -1480 18200 -930 18220
rect -1480 18160 -1470 18200
rect -1970 18150 -1890 18160
rect -1550 18150 -1470 18160
rect -1130 18150 -1050 18160
rect -1970 18130 -1960 18150
rect -2080 18100 -1960 18130
rect -1970 18090 -1960 18100
rect -1900 18090 -1890 18150
rect -1970 18080 -1890 18090
rect -1130 18090 -1120 18150
rect -1060 18130 -1050 18150
rect -1060 18100 -930 18130
rect -1060 18090 -1050 18100
rect -1130 18080 -1050 18090
rect -1560 18050 -1460 18070
rect -1560 17980 -1540 18050
rect -1470 17980 -1460 18050
rect -1560 17940 -1460 17980
rect -1560 17870 -1540 17940
rect -1470 17870 -1460 17940
rect -1560 17860 -1460 17870
rect -1970 17840 -1890 17850
rect -1970 17820 -1960 17840
rect -2080 17790 -1960 17820
rect -1970 17780 -1960 17790
rect -1900 17780 -1890 17840
rect -1130 17840 -1050 17850
rect -1130 17780 -1120 17840
rect -1060 17820 -1050 17840
rect -1060 17790 -930 17820
rect -1060 17780 -1050 17790
rect -1970 17770 -1890 17780
rect -1550 17770 -1470 17780
rect -1130 17770 -1050 17780
rect -1550 17710 -1540 17770
rect -1480 17730 -1470 17770
rect -1480 17710 -930 17730
rect -1550 17700 -930 17710
rect -1020 17230 -930 17240
rect -1020 17170 -1010 17230
rect -940 17170 -930 17230
rect -1020 17160 -930 17170
rect -1010 17090 -930 17100
rect -1010 17030 -1000 17090
rect -940 17030 -930 17090
rect -1010 17020 -930 17030
rect -2080 16980 -2000 16990
rect -2080 16920 -2070 16980
rect -2010 16920 -2000 16980
rect -2080 16910 -2000 16920
rect -1550 16510 -930 16520
rect -1550 16450 -1540 16510
rect -1480 16490 -930 16510
rect -1480 16450 -1470 16490
rect -1970 16440 -1890 16450
rect -1550 16440 -1470 16450
rect -1130 16440 -1050 16450
rect -1970 16420 -1960 16440
rect -2080 16390 -1960 16420
rect -1970 16380 -1960 16390
rect -1900 16380 -1890 16440
rect -1970 16370 -1890 16380
rect -1130 16380 -1120 16440
rect -1060 16420 -1050 16440
rect -1060 16390 -930 16420
rect -1060 16380 -1050 16390
rect -1130 16370 -1050 16380
rect -1560 16340 -1460 16360
rect -1560 16270 -1540 16340
rect -1470 16270 -1460 16340
rect -1560 16230 -1460 16270
rect -1560 16160 -1540 16230
rect -1470 16160 -1460 16230
rect -1560 16150 -1460 16160
rect -1970 16130 -1890 16140
rect -1970 16110 -1960 16130
rect -2080 16080 -1960 16110
rect -1970 16070 -1960 16080
rect -1900 16070 -1890 16130
rect -1130 16130 -1050 16140
rect -1130 16070 -1120 16130
rect -1060 16110 -1050 16130
rect -1060 16080 -930 16110
rect -1060 16070 -1050 16080
rect -1970 16060 -1890 16070
rect -1550 16060 -1470 16070
rect -1130 16060 -1050 16070
rect -1550 16000 -1540 16060
rect -1480 16020 -1470 16060
rect -1480 16000 -930 16020
rect -1550 15990 -930 16000
rect -1020 15520 -930 15530
rect -1020 15460 -1010 15520
rect -940 15460 -930 15520
rect -1020 15450 -930 15460
rect -1010 15380 -930 15390
rect -1010 15320 -1000 15380
rect -940 15320 -930 15380
rect -1010 15310 -930 15320
rect -2080 15270 -2000 15280
rect -2080 15210 -2070 15270
rect -2010 15210 -2000 15270
rect -2080 15200 -2000 15210
rect -1550 14800 -930 14810
rect -1550 14740 -1540 14800
rect -1480 14780 -930 14800
rect -1480 14740 -1470 14780
rect -1970 14730 -1890 14740
rect -1550 14730 -1470 14740
rect -1130 14730 -1050 14740
rect -1970 14710 -1960 14730
rect -2080 14680 -1960 14710
rect -1970 14670 -1960 14680
rect -1900 14670 -1890 14730
rect -1970 14660 -1890 14670
rect -1130 14670 -1120 14730
rect -1060 14710 -1050 14730
rect -1060 14680 -930 14710
rect -1060 14670 -1050 14680
rect -1130 14660 -1050 14670
rect -1560 14630 -1460 14650
rect -1560 14560 -1540 14630
rect -1470 14560 -1460 14630
rect -1560 14520 -1460 14560
rect -1560 14450 -1540 14520
rect -1470 14450 -1460 14520
rect -1560 14440 -1460 14450
rect -1970 14420 -1890 14430
rect -1970 14400 -1960 14420
rect -2080 14370 -1960 14400
rect -1970 14360 -1960 14370
rect -1900 14360 -1890 14420
rect -1130 14420 -1050 14430
rect -1130 14360 -1120 14420
rect -1060 14400 -1050 14420
rect -1060 14370 -930 14400
rect -1060 14360 -1050 14370
rect -1970 14350 -1890 14360
rect -1550 14350 -1470 14360
rect -1130 14350 -1050 14360
rect -1550 14290 -1540 14350
rect -1480 14310 -1470 14350
rect -1480 14290 -930 14310
rect -1550 14280 -930 14290
rect -1020 13810 -930 13820
rect -1020 13750 -1010 13810
rect -940 13750 -930 13810
rect -1020 13740 -930 13750
rect -1010 13670 -930 13680
rect -1010 13610 -1000 13670
rect -940 13610 -930 13670
rect -1010 13600 -930 13610
rect -2080 13560 -2000 13570
rect -2080 13500 -2070 13560
rect -2010 13500 -2000 13560
rect -2080 13490 -2000 13500
rect -1550 13090 -930 13100
rect -1550 13030 -1540 13090
rect -1480 13070 -930 13090
rect -1480 13030 -1470 13070
rect -1970 13020 -1890 13030
rect -1550 13020 -1470 13030
rect -1130 13020 -1050 13030
rect -1970 13000 -1960 13020
rect -2080 12970 -1960 13000
rect -1970 12960 -1960 12970
rect -1900 12960 -1890 13020
rect -1970 12950 -1890 12960
rect -1130 12960 -1120 13020
rect -1060 13000 -1050 13020
rect -1060 12970 -930 13000
rect -1060 12960 -1050 12970
rect -1130 12950 -1050 12960
rect -1560 12920 -1460 12940
rect -1560 12850 -1540 12920
rect -1470 12850 -1460 12920
rect -1560 12810 -1460 12850
rect -1560 12740 -1540 12810
rect -1470 12740 -1460 12810
rect -1560 12730 -1460 12740
rect -1970 12710 -1890 12720
rect -1970 12690 -1960 12710
rect -2080 12660 -1960 12690
rect -1970 12650 -1960 12660
rect -1900 12650 -1890 12710
rect -1130 12710 -1050 12720
rect -1130 12650 -1120 12710
rect -1060 12690 -1050 12710
rect -1060 12660 -930 12690
rect -1060 12650 -1050 12660
rect -1970 12640 -1890 12650
rect -1550 12640 -1470 12650
rect -1130 12640 -1050 12650
rect -1550 12580 -1540 12640
rect -1480 12600 -1470 12640
rect -1480 12580 -930 12600
rect -1550 12570 -930 12580
rect -1020 12100 -930 12110
rect -1020 12040 -1010 12100
rect -940 12040 -930 12100
rect -1020 12030 -930 12040
rect -1010 11960 -930 11970
rect -1010 11900 -1000 11960
rect -940 11900 -930 11960
rect -1010 11890 -930 11900
rect -2080 11850 -2000 11860
rect -2080 11790 -2070 11850
rect -2010 11790 -2000 11850
rect -2080 11780 -2000 11790
rect -1550 11380 -930 11390
rect -1550 11320 -1540 11380
rect -1480 11360 -930 11380
rect -1480 11320 -1470 11360
rect -1970 11310 -1890 11320
rect -1550 11310 -1470 11320
rect -1130 11310 -1050 11320
rect -1970 11290 -1960 11310
rect -2080 11260 -1960 11290
rect -1970 11250 -1960 11260
rect -1900 11250 -1890 11310
rect -1970 11240 -1890 11250
rect -1130 11250 -1120 11310
rect -1060 11290 -1050 11310
rect -1060 11260 -930 11290
rect -1060 11250 -1050 11260
rect -1130 11240 -1050 11250
rect -1560 11210 -1460 11230
rect -1560 11140 -1540 11210
rect -1470 11140 -1460 11210
rect -1560 11100 -1460 11140
rect -1560 11030 -1540 11100
rect -1470 11030 -1460 11100
rect -1560 11020 -1460 11030
rect -1970 11000 -1890 11010
rect -1970 10980 -1960 11000
rect -2080 10950 -1960 10980
rect -1970 10940 -1960 10950
rect -1900 10940 -1890 11000
rect -1130 11000 -1050 11010
rect -1130 10940 -1120 11000
rect -1060 10980 -1050 11000
rect -1060 10950 -930 10980
rect -1060 10940 -1050 10950
rect -1970 10930 -1890 10940
rect -1550 10930 -1470 10940
rect -1130 10930 -1050 10940
rect -1550 10870 -1540 10930
rect -1480 10890 -1470 10930
rect -1480 10870 -930 10890
rect -1550 10860 -930 10870
rect -1020 10390 -930 10400
rect -1020 10330 -1010 10390
rect -940 10330 -930 10390
rect -1020 10320 -930 10330
rect -1010 10250 -930 10260
rect -1010 10190 -1000 10250
rect -940 10190 -930 10250
rect -1010 10180 -930 10190
rect -2080 10140 -2000 10150
rect -2080 10080 -2070 10140
rect -2010 10080 -2000 10140
rect -2080 10070 -2000 10080
rect -1550 9670 -930 9680
rect -1550 9610 -1540 9670
rect -1480 9650 -930 9670
rect -1480 9610 -1470 9650
rect -1970 9600 -1890 9610
rect -1550 9600 -1470 9610
rect -1130 9600 -1050 9610
rect -1970 9580 -1960 9600
rect -2080 9550 -1960 9580
rect -1970 9540 -1960 9550
rect -1900 9540 -1890 9600
rect -1970 9530 -1890 9540
rect -1130 9540 -1120 9600
rect -1060 9580 -1050 9600
rect -1060 9550 -930 9580
rect -1060 9540 -1050 9550
rect -1130 9530 -1050 9540
rect -1560 9500 -1460 9520
rect -1560 9430 -1540 9500
rect -1470 9430 -1460 9500
rect -1560 9390 -1460 9430
rect -1560 9320 -1540 9390
rect -1470 9320 -1460 9390
rect -1560 9310 -1460 9320
rect -1970 9290 -1890 9300
rect -1970 9270 -1960 9290
rect -2080 9240 -1960 9270
rect -1970 9230 -1960 9240
rect -1900 9230 -1890 9290
rect -1130 9290 -1050 9300
rect -1130 9230 -1120 9290
rect -1060 9270 -1050 9290
rect -1060 9240 -930 9270
rect -1060 9230 -1050 9240
rect -1970 9220 -1890 9230
rect -1550 9220 -1470 9230
rect -1130 9220 -1050 9230
rect -1550 9160 -1540 9220
rect -1480 9180 -1470 9220
rect -1480 9160 -930 9180
rect -1550 9150 -930 9160
rect -1020 8680 -930 8690
rect -1020 8620 -1010 8680
rect -940 8620 -930 8680
rect -1020 8610 -930 8620
rect -1010 8540 -930 8550
rect -1010 8480 -1000 8540
rect -940 8480 -930 8540
rect -1010 8470 -930 8480
rect -2080 8430 -2000 8440
rect -2080 8370 -2070 8430
rect -2010 8370 -2000 8430
rect -2080 8360 -2000 8370
rect -1550 7960 -930 7970
rect -1550 7900 -1540 7960
rect -1480 7940 -930 7960
rect -1480 7900 -1470 7940
rect -1970 7890 -1890 7900
rect -1550 7890 -1470 7900
rect -1130 7890 -1050 7900
rect -1970 7870 -1960 7890
rect -2080 7840 -1960 7870
rect -1970 7830 -1960 7840
rect -1900 7830 -1890 7890
rect -1970 7820 -1890 7830
rect -1130 7830 -1120 7890
rect -1060 7870 -1050 7890
rect -1060 7840 -930 7870
rect -1060 7830 -1050 7840
rect -1130 7820 -1050 7830
rect -1560 7790 -1460 7810
rect -1560 7720 -1540 7790
rect -1470 7720 -1460 7790
rect -1560 7680 -1460 7720
rect -1560 7610 -1540 7680
rect -1470 7610 -1460 7680
rect -1560 7600 -1460 7610
rect -1970 7580 -1890 7590
rect -1970 7560 -1960 7580
rect -2080 7530 -1960 7560
rect -1970 7520 -1960 7530
rect -1900 7520 -1890 7580
rect -1130 7580 -1050 7590
rect -1130 7520 -1120 7580
rect -1060 7560 -1050 7580
rect -1060 7530 -930 7560
rect -1060 7520 -1050 7530
rect -1970 7510 -1890 7520
rect -1550 7510 -1470 7520
rect -1130 7510 -1050 7520
rect -1550 7450 -1540 7510
rect -1480 7470 -1470 7510
rect -1480 7450 -930 7470
rect -1550 7440 -930 7450
rect -1020 6970 -930 6980
rect -1020 6910 -1010 6970
rect -940 6910 -930 6970
rect -1020 6900 -930 6910
rect -1010 6830 -930 6840
rect -1010 6770 -1000 6830
rect -940 6770 -930 6830
rect -1010 6760 -930 6770
rect -2080 6720 -2000 6730
rect -2080 6660 -2070 6720
rect -2010 6660 -2000 6720
rect -2080 6650 -2000 6660
rect -1550 6250 -930 6260
rect -1550 6190 -1540 6250
rect -1480 6230 -930 6250
rect -1480 6190 -1470 6230
rect -1970 6180 -1890 6190
rect -1550 6180 -1470 6190
rect -1130 6180 -1050 6190
rect -1970 6160 -1960 6180
rect -2080 6130 -1960 6160
rect -1970 6120 -1960 6130
rect -1900 6120 -1890 6180
rect -1970 6110 -1890 6120
rect -1130 6120 -1120 6180
rect -1060 6160 -1050 6180
rect -1060 6130 -930 6160
rect -1060 6120 -1050 6130
rect -1130 6110 -1050 6120
rect -1560 6080 -1460 6100
rect -1560 6010 -1540 6080
rect -1470 6010 -1460 6080
rect -1560 5970 -1460 6010
rect -1560 5900 -1540 5970
rect -1470 5900 -1460 5970
rect -1560 5890 -1460 5900
rect -1970 5870 -1890 5880
rect -1970 5850 -1960 5870
rect -2080 5820 -1960 5850
rect -1970 5810 -1960 5820
rect -1900 5810 -1890 5870
rect -1130 5870 -1050 5880
rect -1130 5810 -1120 5870
rect -1060 5850 -1050 5870
rect -1060 5820 -930 5850
rect -1060 5810 -1050 5820
rect -1970 5800 -1890 5810
rect -1550 5800 -1470 5810
rect -1130 5800 -1050 5810
rect -1550 5740 -1540 5800
rect -1480 5760 -1470 5800
rect -1480 5740 -930 5760
rect -1550 5730 -930 5740
rect -1020 5260 -930 5270
rect -1020 5200 -1010 5260
rect -940 5200 -930 5260
rect -1020 5190 -930 5200
rect -1010 5120 -930 5130
rect -1010 5060 -1000 5120
rect -940 5060 -930 5120
rect -1010 5050 -930 5060
rect -2080 5010 -2000 5020
rect -2080 4950 -2070 5010
rect -2010 4950 -2000 5010
rect -2080 4940 -2000 4950
rect -1550 4540 -930 4550
rect -1550 4480 -1540 4540
rect -1480 4520 -930 4540
rect -1480 4480 -1470 4520
rect -1970 4470 -1890 4480
rect -1550 4470 -1470 4480
rect -1130 4470 -1050 4480
rect -1970 4450 -1960 4470
rect -2080 4420 -1960 4450
rect -1970 4410 -1960 4420
rect -1900 4410 -1890 4470
rect -1970 4400 -1890 4410
rect -1130 4410 -1120 4470
rect -1060 4450 -1050 4470
rect -1060 4420 -930 4450
rect -1060 4410 -1050 4420
rect -1130 4400 -1050 4410
rect -1560 4370 -1460 4390
rect -1560 4300 -1540 4370
rect -1470 4300 -1460 4370
rect -1560 4260 -1460 4300
rect -1560 4190 -1540 4260
rect -1470 4190 -1460 4260
rect -1560 4180 -1460 4190
rect -1970 4160 -1890 4170
rect -1970 4140 -1960 4160
rect -2080 4110 -1960 4140
rect -1970 4100 -1960 4110
rect -1900 4100 -1890 4160
rect -1130 4160 -1050 4170
rect -1130 4100 -1120 4160
rect -1060 4140 -1050 4160
rect -1060 4110 -930 4140
rect -1060 4100 -1050 4110
rect -1970 4090 -1890 4100
rect -1550 4090 -1470 4100
rect -1130 4090 -1050 4100
rect -1550 4030 -1540 4090
rect -1480 4050 -1470 4090
rect -1480 4030 -930 4050
rect -1550 4020 -930 4030
rect -1020 3550 -930 3560
rect -1020 3490 -1010 3550
rect -940 3490 -930 3550
rect -1020 3480 -930 3490
rect -1010 3410 -930 3420
rect -1010 3350 -1000 3410
rect -940 3350 -930 3410
rect -1010 3340 -930 3350
rect -2080 3300 -2000 3310
rect -2080 3240 -2070 3300
rect -2010 3240 -2000 3300
rect -2080 3230 -2000 3240
rect -1550 2830 -930 2840
rect -1550 2770 -1540 2830
rect -1480 2810 -930 2830
rect -1480 2770 -1470 2810
rect -1970 2760 -1890 2770
rect -1550 2760 -1470 2770
rect -1130 2760 -1050 2770
rect -1970 2740 -1960 2760
rect -2080 2710 -1960 2740
rect -1970 2700 -1960 2710
rect -1900 2700 -1890 2760
rect -1970 2690 -1890 2700
rect -1130 2700 -1120 2760
rect -1060 2740 -1050 2760
rect -1060 2710 -930 2740
rect -1060 2700 -1050 2710
rect -1130 2690 -1050 2700
rect -1560 2660 -1460 2680
rect -1560 2590 -1540 2660
rect -1470 2590 -1460 2660
rect -1560 2550 -1460 2590
rect -1560 2480 -1540 2550
rect -1470 2480 -1460 2550
rect -1560 2470 -1460 2480
rect -1970 2450 -1890 2460
rect -1970 2430 -1960 2450
rect -2080 2400 -1960 2430
rect -1970 2390 -1960 2400
rect -1900 2390 -1890 2450
rect -1130 2450 -1050 2460
rect -1130 2390 -1120 2450
rect -1060 2430 -1050 2450
rect -1060 2400 -930 2430
rect -1060 2390 -1050 2400
rect -1970 2380 -1890 2390
rect -1550 2380 -1470 2390
rect -1130 2380 -1050 2390
rect -1550 2320 -1540 2380
rect -1480 2340 -1470 2380
rect -1480 2320 -930 2340
rect -1550 2310 -930 2320
rect -1020 1840 -930 1850
rect -1020 1780 -1010 1840
rect -940 1780 -930 1840
rect -1020 1770 -930 1780
rect -1010 1700 -930 1710
rect -1010 1640 -1000 1700
rect -940 1640 -930 1700
rect -1010 1630 -930 1640
rect -2080 1590 -2000 1600
rect -2080 1530 -2070 1590
rect -2010 1530 -2000 1590
rect -2080 1520 -2000 1530
rect -1550 1120 -930 1130
rect -1550 1060 -1540 1120
rect -1480 1100 -930 1120
rect -1480 1060 -1470 1100
rect -1970 1050 -1890 1060
rect -1550 1050 -1470 1060
rect -1130 1050 -1050 1060
rect -1970 1030 -1960 1050
rect -2080 1000 -1960 1030
rect -1970 990 -1960 1000
rect -1900 990 -1890 1050
rect -1970 980 -1890 990
rect -1130 990 -1120 1050
rect -1060 1030 -1050 1050
rect -1060 1000 -930 1030
rect -1060 990 -1050 1000
rect -1130 980 -1050 990
rect -1560 950 -1460 970
rect -1560 880 -1540 950
rect -1470 880 -1460 950
rect -1560 840 -1460 880
rect -1560 770 -1540 840
rect -1470 770 -1460 840
rect -1560 760 -1460 770
rect -1970 740 -1890 750
rect -1970 720 -1960 740
rect -2080 690 -1960 720
rect -1970 680 -1960 690
rect -1900 680 -1890 740
rect -1130 740 -1050 750
rect -1130 680 -1120 740
rect -1060 720 -1050 740
rect -1060 690 -930 720
rect -1060 680 -1050 690
rect -1970 670 -1890 680
rect -1550 670 -1470 680
rect -1130 670 -1050 680
rect -1550 610 -1540 670
rect -1480 630 -1470 670
rect -1480 610 -930 630
rect -1550 600 -930 610
rect -2080 140 -2000 150
rect -750 140 -720 23940
rect -630 140 -600 23940
rect -510 140 -480 23940
rect -390 140 -360 23940
rect -270 140 -240 23940
rect -150 140 -120 23940
rect -30 140 0 23940
rect -2080 80 -2070 140
rect -2010 80 -2000 140
rect -2080 70 -2000 80
rect -1020 130 -930 140
rect -1020 70 -1010 130
rect -940 70 -930 130
rect -1020 60 -930 70
rect -1010 -10 -930 0
rect -1010 -70 -1000 -10
rect -940 -70 -930 -10
rect -1010 -80 -930 -70
rect -2080 -120 -2000 -110
rect -2080 -180 -2070 -120
rect -2010 -180 -2000 -120
rect -2080 -190 -2000 -180
rect -1550 -590 -930 -580
rect -1550 -650 -1540 -590
rect -1480 -610 -930 -590
rect -1480 -650 -1470 -610
rect -1970 -660 -1890 -650
rect -1550 -660 -1470 -650
rect -1130 -660 -1050 -650
rect -1970 -680 -1960 -660
rect -2080 -710 -1960 -680
rect -1970 -720 -1960 -710
rect -1900 -720 -1890 -660
rect -1970 -730 -1890 -720
rect -1130 -720 -1120 -660
rect -1060 -680 -1050 -660
rect -1060 -710 -930 -680
rect -1060 -720 -1050 -710
rect -1130 -730 -1050 -720
rect -1560 -760 -1460 -740
rect -1560 -830 -1540 -760
rect -1470 -830 -1460 -760
rect -1560 -870 -1460 -830
rect -1560 -940 -1540 -870
rect -1470 -940 -1460 -870
rect -1560 -950 -1460 -940
rect -1970 -970 -1890 -960
rect -1970 -990 -1960 -970
rect -2080 -1020 -1960 -990
rect -1970 -1030 -1960 -1020
rect -1900 -1030 -1890 -970
rect -1130 -970 -1050 -960
rect -1130 -1030 -1120 -970
rect -1060 -990 -1050 -970
rect -1060 -1020 -930 -990
rect -1060 -1030 -1050 -1020
rect -1970 -1040 -1890 -1030
rect -1550 -1040 -1470 -1030
rect -1130 -1040 -1050 -1030
rect -1550 -1100 -1540 -1040
rect -1480 -1080 -1470 -1040
rect -1480 -1100 -930 -1080
rect -1550 -1110 -930 -1100
rect -1020 -1580 -930 -1570
rect -1020 -1640 -1010 -1580
rect -940 -1640 -930 -1580
rect -1020 -1650 -930 -1640
rect -750 -1710 -720 -110
rect -630 -1710 -600 -110
rect -510 -1710 -480 -110
rect -390 -1710 -360 -110
rect -270 -1710 -240 -110
rect -150 -1710 -120 -110
rect -30 -1710 0 -110
rect 1860 -1710 1890 150
rect 1980 -1710 2010 150
rect 2100 -1710 2130 150
rect 2220 -1710 2250 150
rect 2340 -1710 2370 150
rect 2460 -1710 2490 150
rect 2580 -1710 2610 150
rect 2640 140 2720 150
rect 2640 80 2650 140
rect 2710 80 2720 140
rect 2640 70 2720 80
rect 3820 40 3940 70
rect 3710 -10 3790 0
rect 3710 -70 3720 -10
rect 3780 -70 3790 -10
rect 3820 -20 3860 40
rect 3920 -20 3940 40
rect 3820 -50 3940 -20
rect 3710 -80 3790 -70
rect 2640 -120 2720 -110
rect 2640 -180 2650 -120
rect 2710 -180 2720 -120
rect 2640 -190 2720 -180
rect 3170 -590 3790 -580
rect 3170 -650 3180 -590
rect 3240 -610 3790 -590
rect 3240 -650 3250 -610
rect 2750 -660 2830 -650
rect 3170 -660 3250 -650
rect 3590 -660 3670 -650
rect 2750 -680 2760 -660
rect 2640 -710 2760 -680
rect 2750 -720 2760 -710
rect 2820 -720 2830 -660
rect 2750 -730 2830 -720
rect 3590 -720 3600 -660
rect 3660 -680 3670 -660
rect 3660 -710 3790 -680
rect 3660 -720 3670 -710
rect 3590 -730 3670 -720
rect 3160 -760 3260 -740
rect 3160 -830 3180 -760
rect 3250 -830 3260 -760
rect 3160 -870 3260 -830
rect 3160 -940 3180 -870
rect 3250 -940 3260 -870
rect 3160 -950 3260 -940
rect 2750 -970 2830 -960
rect 2750 -990 2760 -970
rect 2640 -1020 2760 -990
rect 2750 -1030 2760 -1020
rect 2820 -1030 2830 -970
rect 3590 -970 3670 -960
rect 3590 -1030 3600 -970
rect 3660 -990 3670 -970
rect 3660 -1020 3790 -990
rect 3660 -1030 3670 -1020
rect 2750 -1040 2830 -1030
rect 3170 -1040 3250 -1030
rect 3590 -1040 3670 -1030
rect 3170 -1100 3180 -1040
rect 3240 -1080 3250 -1040
rect 3240 -1100 3790 -1080
rect 3170 -1110 3790 -1100
rect 3710 -1640 3790 -1630
rect 3710 -1700 3720 -1640
rect 3780 -1700 3790 -1640
rect 3710 -1710 3790 -1700
rect 3970 -1710 4000 0
rect 4090 -1710 4120 0
rect 4210 -1710 4240 0
rect 4330 -1710 4360 0
rect 4450 -1710 4480 0
rect 4570 -1710 4600 0
rect 4690 -1710 4720 0
rect 6850 -1710 6880 150
rect 6970 -1710 7000 150
rect 7090 -1710 7120 150
rect 7210 -1710 7240 150
rect 7330 -1710 7360 150
rect 7450 -1710 7480 150
rect 7570 -1710 7600 150
rect 7630 140 7710 150
rect 7630 80 7640 140
rect 7700 80 7710 140
rect 7630 70 7710 80
rect 8810 40 8930 70
rect 8700 -10 8780 0
rect 8700 -70 8710 -10
rect 8770 -70 8780 -10
rect 8810 -20 8850 40
rect 8910 -20 8930 40
rect 8810 -50 8930 -20
rect 8700 -80 8780 -70
rect 7630 -120 7710 -110
rect 7630 -180 7640 -120
rect 7700 -180 7710 -120
rect 7630 -190 7710 -180
rect 8160 -590 8780 -580
rect 8160 -650 8170 -590
rect 8230 -610 8780 -590
rect 8230 -650 8240 -610
rect 7740 -660 7820 -650
rect 8160 -660 8240 -650
rect 8580 -660 8660 -650
rect 7740 -680 7750 -660
rect 7630 -710 7750 -680
rect 7740 -720 7750 -710
rect 7810 -720 7820 -660
rect 7740 -730 7820 -720
rect 8580 -720 8590 -660
rect 8650 -680 8660 -660
rect 8650 -710 8780 -680
rect 8650 -720 8660 -710
rect 8580 -730 8660 -720
rect 8150 -760 8250 -740
rect 8150 -830 8170 -760
rect 8240 -830 8250 -760
rect 8150 -870 8250 -830
rect 8150 -940 8170 -870
rect 8240 -940 8250 -870
rect 8150 -950 8250 -940
rect 7740 -970 7820 -960
rect 7740 -990 7750 -970
rect 7630 -1020 7750 -990
rect 7740 -1030 7750 -1020
rect 7810 -1030 7820 -970
rect 8580 -970 8660 -960
rect 8580 -1030 8590 -970
rect 8650 -990 8660 -970
rect 8650 -1020 8780 -990
rect 8650 -1030 8660 -1020
rect 7740 -1040 7820 -1030
rect 8160 -1040 8240 -1030
rect 8580 -1040 8660 -1030
rect 8160 -1100 8170 -1040
rect 8230 -1080 8240 -1040
rect 8230 -1100 8780 -1080
rect 8160 -1110 8780 -1100
rect 8700 -1640 8780 -1630
rect 8700 -1700 8710 -1640
rect 8770 -1700 8780 -1640
rect 8700 -1710 8780 -1700
rect 8960 -1710 8990 130
rect 9080 -1710 9110 0
rect 9200 -1710 9230 0
rect 9320 -1710 9350 0
rect 9440 -1710 9470 0
rect 9560 -1710 9590 0
rect 9680 -1710 9710 0
rect 11840 -1710 11870 150
rect 11960 -1710 11990 150
rect 12080 -1710 12110 150
rect 12200 -1710 12230 150
rect 12320 -1710 12350 150
rect 12440 -1710 12470 150
rect 12560 -1710 12590 150
rect 12620 140 12700 150
rect 12620 80 12630 140
rect 12690 80 12700 140
rect 12620 70 12700 80
rect 13800 40 13920 70
rect 13690 -10 13770 0
rect 13690 -70 13700 -10
rect 13760 -70 13770 -10
rect 13800 -20 13840 40
rect 13900 -20 13920 40
rect 13800 -50 13920 -20
rect 13690 -80 13770 -70
rect 12620 -120 12700 -110
rect 12620 -180 12630 -120
rect 12690 -180 12700 -120
rect 12620 -190 12700 -180
rect 13150 -590 13770 -580
rect 13150 -650 13160 -590
rect 13220 -610 13770 -590
rect 13220 -650 13230 -610
rect 12730 -660 12810 -650
rect 13150 -660 13230 -650
rect 13570 -660 13650 -650
rect 12730 -680 12740 -660
rect 12620 -710 12740 -680
rect 12730 -720 12740 -710
rect 12800 -720 12810 -660
rect 12730 -730 12810 -720
rect 13570 -720 13580 -660
rect 13640 -680 13650 -660
rect 13640 -710 13770 -680
rect 13640 -720 13650 -710
rect 13570 -730 13650 -720
rect 13140 -760 13240 -740
rect 13140 -830 13160 -760
rect 13230 -830 13240 -760
rect 13140 -870 13240 -830
rect 13140 -940 13160 -870
rect 13230 -940 13240 -870
rect 13140 -950 13240 -940
rect 12730 -970 12810 -960
rect 12730 -990 12740 -970
rect 12620 -1020 12740 -990
rect 12730 -1030 12740 -1020
rect 12800 -1030 12810 -970
rect 13570 -970 13650 -960
rect 13570 -1030 13580 -970
rect 13640 -990 13650 -970
rect 13640 -1020 13770 -990
rect 13640 -1030 13650 -1020
rect 12730 -1040 12810 -1030
rect 13150 -1040 13230 -1030
rect 13570 -1040 13650 -1030
rect 13150 -1100 13160 -1040
rect 13220 -1080 13230 -1040
rect 13220 -1100 13770 -1080
rect 13150 -1110 13770 -1100
rect 13690 -1640 13770 -1630
rect 13690 -1700 13700 -1640
rect 13760 -1700 13770 -1640
rect 13690 -1710 13770 -1700
rect 13950 -1710 13980 130
rect 14070 -1710 14100 0
rect 14190 -1710 14220 0
rect 14310 -1710 14340 0
rect 14430 -1710 14460 0
rect 14550 -1710 14580 0
rect 14670 -1710 14700 0
rect 16830 -1710 16860 150
rect 16950 -1710 16980 150
rect 17070 -1710 17100 150
rect 17190 -1710 17220 150
rect 17310 -1710 17340 150
rect 17430 -1710 17460 150
rect 17550 -1710 17580 150
rect 17610 140 17690 150
rect 17610 80 17620 140
rect 17680 80 17690 140
rect 17610 70 17690 80
rect 18790 40 18910 70
rect 18680 -10 18760 0
rect 18680 -70 18690 -10
rect 18750 -70 18760 -10
rect 18790 -20 18830 40
rect 18890 -20 18910 40
rect 18790 -50 18910 -20
rect 18680 -80 18760 -70
rect 17610 -120 17690 -110
rect 17610 -180 17620 -120
rect 17680 -180 17690 -120
rect 17610 -190 17690 -180
rect 18140 -590 18760 -580
rect 18140 -650 18150 -590
rect 18210 -610 18760 -590
rect 18210 -650 18220 -610
rect 17720 -660 17800 -650
rect 18140 -660 18220 -650
rect 18560 -660 18640 -650
rect 17720 -680 17730 -660
rect 17610 -710 17730 -680
rect 17720 -720 17730 -710
rect 17790 -720 17800 -660
rect 17720 -730 17800 -720
rect 18560 -720 18570 -660
rect 18630 -680 18640 -660
rect 18630 -710 18760 -680
rect 18630 -720 18640 -710
rect 18560 -730 18640 -720
rect 18130 -760 18230 -740
rect 18130 -830 18150 -760
rect 18220 -830 18230 -760
rect 18130 -870 18230 -830
rect 18130 -940 18150 -870
rect 18220 -940 18230 -870
rect 18130 -950 18230 -940
rect 17720 -970 17800 -960
rect 17720 -990 17730 -970
rect 17610 -1020 17730 -990
rect 17720 -1030 17730 -1020
rect 17790 -1030 17800 -970
rect 18560 -970 18640 -960
rect 18560 -1030 18570 -970
rect 18630 -990 18640 -970
rect 18630 -1020 18760 -990
rect 18630 -1030 18640 -1020
rect 17720 -1040 17800 -1030
rect 18140 -1040 18220 -1030
rect 18560 -1040 18640 -1030
rect 18140 -1100 18150 -1040
rect 18210 -1080 18220 -1040
rect 18210 -1100 18760 -1080
rect 18140 -1110 18760 -1100
rect 18680 -1640 18760 -1630
rect 18680 -1700 18690 -1640
rect 18750 -1700 18760 -1640
rect 18680 -1710 18760 -1700
rect 18940 -1710 18970 130
rect 19060 -1710 19090 0
rect 19180 -1710 19210 0
rect 19300 -1710 19330 0
rect 19420 -1710 19450 0
rect 19540 -1710 19570 0
rect 19660 -1710 19690 0
rect 21820 -1710 21850 150
rect 21940 -1710 21970 150
rect 22060 -1710 22090 150
rect 22180 -1710 22210 150
rect 22300 -1710 22330 150
rect 22420 -1710 22450 150
rect 22540 -1710 22570 150
rect 22600 140 22680 150
rect 22600 80 22610 140
rect 22670 80 22680 140
rect 22600 70 22680 80
rect 23780 40 23900 70
rect 23670 -10 23750 0
rect 23670 -70 23680 -10
rect 23740 -70 23750 -10
rect 23780 -20 23820 40
rect 23880 -20 23900 40
rect 23780 -50 23900 -20
rect 23670 -80 23750 -70
rect 22600 -120 22680 -110
rect 22600 -180 22610 -120
rect 22670 -180 22680 -120
rect 22600 -190 22680 -180
rect 23130 -590 23750 -580
rect 23130 -650 23140 -590
rect 23200 -610 23750 -590
rect 23200 -650 23210 -610
rect 22710 -660 22790 -650
rect 23130 -660 23210 -650
rect 23550 -660 23630 -650
rect 22710 -680 22720 -660
rect 22600 -710 22720 -680
rect 22710 -720 22720 -710
rect 22780 -720 22790 -660
rect 22710 -730 22790 -720
rect 23550 -720 23560 -660
rect 23620 -680 23630 -660
rect 23620 -710 23750 -680
rect 23620 -720 23630 -710
rect 23550 -730 23630 -720
rect 23120 -760 23220 -740
rect 23120 -830 23140 -760
rect 23210 -830 23220 -760
rect 23120 -870 23220 -830
rect 23120 -940 23140 -870
rect 23210 -940 23220 -870
rect 23120 -950 23220 -940
rect 22710 -970 22790 -960
rect 22710 -990 22720 -970
rect 22600 -1020 22720 -990
rect 22710 -1030 22720 -1020
rect 22780 -1030 22790 -970
rect 23550 -970 23630 -960
rect 23550 -1030 23560 -970
rect 23620 -990 23630 -970
rect 23620 -1020 23750 -990
rect 23620 -1030 23630 -1020
rect 22710 -1040 22790 -1030
rect 23130 -1040 23210 -1030
rect 23550 -1040 23630 -1030
rect 23130 -1100 23140 -1040
rect 23200 -1080 23210 -1040
rect 23200 -1100 23750 -1080
rect 23130 -1110 23750 -1100
rect 23670 -1640 23750 -1630
rect 23670 -1700 23680 -1640
rect 23740 -1700 23750 -1640
rect 23670 -1710 23750 -1700
rect 23930 -1710 23960 130
rect 24050 -1710 24080 0
rect 24170 -1710 24200 0
rect 24290 -1710 24320 0
rect 24410 -1710 24440 0
rect 24530 -1710 24560 0
rect 24650 -1710 24680 0
rect 26810 -1710 26840 150
rect 26930 -1710 26960 150
rect 27050 -1710 27080 150
rect 27170 -1710 27200 150
rect 27290 -1710 27320 150
rect 27410 -1710 27440 150
rect 27530 -1710 27560 150
rect 27590 140 27670 150
rect 27590 80 27600 140
rect 27660 80 27670 140
rect 27590 70 27670 80
rect 28770 40 28890 70
rect 28660 -10 28740 0
rect 28660 -70 28670 -10
rect 28730 -70 28740 -10
rect 28770 -20 28810 40
rect 28870 -20 28890 40
rect 28770 -50 28890 -20
rect 28660 -80 28740 -70
rect 27590 -120 27670 -110
rect 27590 -180 27600 -120
rect 27660 -180 27670 -120
rect 27590 -190 27670 -180
rect 28120 -590 28740 -580
rect 28120 -650 28130 -590
rect 28190 -610 28740 -590
rect 28190 -650 28200 -610
rect 27700 -660 27780 -650
rect 28120 -660 28200 -650
rect 28540 -660 28620 -650
rect 27700 -680 27710 -660
rect 27590 -710 27710 -680
rect 27700 -720 27710 -710
rect 27770 -720 27780 -660
rect 27700 -730 27780 -720
rect 28540 -720 28550 -660
rect 28610 -680 28620 -660
rect 28610 -710 28740 -680
rect 28610 -720 28620 -710
rect 28540 -730 28620 -720
rect 28110 -760 28210 -740
rect 28110 -830 28130 -760
rect 28200 -830 28210 -760
rect 28110 -870 28210 -830
rect 28110 -940 28130 -870
rect 28200 -940 28210 -870
rect 28110 -950 28210 -940
rect 27700 -970 27780 -960
rect 27700 -990 27710 -970
rect 27590 -1020 27710 -990
rect 27700 -1030 27710 -1020
rect 27770 -1030 27780 -970
rect 28540 -970 28620 -960
rect 28540 -1030 28550 -970
rect 28610 -990 28620 -970
rect 28610 -1020 28740 -990
rect 28610 -1030 28620 -1020
rect 27700 -1040 27780 -1030
rect 28120 -1040 28200 -1030
rect 28540 -1040 28620 -1030
rect 28120 -1100 28130 -1040
rect 28190 -1080 28200 -1040
rect 28190 -1100 28740 -1080
rect 28120 -1110 28740 -1100
rect 28660 -1640 28740 -1630
rect 28660 -1700 28670 -1640
rect 28730 -1700 28740 -1640
rect 28660 -1710 28740 -1700
rect 28920 -1710 28950 130
rect 29040 -1710 29070 0
rect 29160 -1710 29190 0
rect 29280 -1710 29310 0
rect 29400 -1710 29430 0
rect 29520 -1710 29550 0
rect 29640 -1710 29670 0
rect 31800 -1710 31830 150
rect 31920 -1710 31950 150
rect 32040 -1710 32070 150
rect 32160 -1710 32190 150
rect 32280 -1710 32310 150
rect 32400 -1710 32430 150
rect 32520 -1710 32550 150
rect 32580 140 32660 150
rect 32580 80 32590 140
rect 32650 80 32660 140
rect 32580 70 32660 80
rect 33760 40 33880 70
rect 33650 -10 33730 0
rect 33650 -70 33660 -10
rect 33720 -70 33730 -10
rect 33760 -20 33800 40
rect 33860 -20 33880 40
rect 33760 -50 33880 -20
rect 33650 -80 33730 -70
rect 32580 -120 32660 -110
rect 32580 -180 32590 -120
rect 32650 -180 32660 -120
rect 32580 -190 32660 -180
rect 33110 -590 33730 -580
rect 33110 -650 33120 -590
rect 33180 -610 33730 -590
rect 33180 -650 33190 -610
rect 32690 -660 32770 -650
rect 33110 -660 33190 -650
rect 33530 -660 33610 -650
rect 32690 -680 32700 -660
rect 32580 -710 32700 -680
rect 32690 -720 32700 -710
rect 32760 -720 32770 -660
rect 32690 -730 32770 -720
rect 33530 -720 33540 -660
rect 33600 -680 33610 -660
rect 33600 -710 33730 -680
rect 33600 -720 33610 -710
rect 33530 -730 33610 -720
rect 33100 -760 33200 -740
rect 33100 -830 33120 -760
rect 33190 -830 33200 -760
rect 33100 -870 33200 -830
rect 33100 -940 33120 -870
rect 33190 -940 33200 -870
rect 33100 -950 33200 -940
rect 32690 -970 32770 -960
rect 32690 -990 32700 -970
rect 32580 -1020 32700 -990
rect 32690 -1030 32700 -1020
rect 32760 -1030 32770 -970
rect 33530 -970 33610 -960
rect 33530 -1030 33540 -970
rect 33600 -990 33610 -970
rect 33600 -1020 33730 -990
rect 33600 -1030 33610 -1020
rect 32690 -1040 32770 -1030
rect 33110 -1040 33190 -1030
rect 33530 -1040 33610 -1030
rect 33110 -1100 33120 -1040
rect 33180 -1080 33190 -1040
rect 33180 -1100 33730 -1080
rect 33110 -1110 33730 -1100
rect 33650 -1640 33730 -1630
rect 33650 -1700 33660 -1640
rect 33720 -1700 33730 -1640
rect 33650 -1710 33730 -1700
rect 33910 -1710 33940 130
rect 34030 -1710 34060 0
rect 34150 -1710 34180 0
rect 34270 -1710 34300 0
rect 34390 -1710 34420 0
rect 34510 -1710 34540 0
rect 34630 -1710 34660 0
rect 36790 -1710 36820 150
rect 36910 -1710 36940 150
rect 37030 -1710 37060 150
rect 37150 -1710 37180 150
rect 37270 -1710 37300 150
rect 37390 -1710 37420 150
rect 37510 -1710 37540 150
rect 37570 140 37650 150
rect 37570 80 37580 140
rect 37640 80 37650 140
rect 37570 70 37650 80
rect 38750 40 38870 70
rect 38640 -10 38720 0
rect 38640 -70 38650 -10
rect 38710 -70 38720 -10
rect 38750 -20 38790 40
rect 38850 -20 38870 40
rect 38750 -50 38870 -20
rect 38640 -80 38720 -70
rect 37570 -120 37650 -110
rect 37570 -180 37580 -120
rect 37640 -180 37650 -120
rect 37570 -190 37650 -180
rect 38100 -590 38720 -580
rect 38100 -650 38110 -590
rect 38170 -610 38720 -590
rect 38170 -650 38180 -610
rect 37680 -660 37760 -650
rect 38100 -660 38180 -650
rect 38520 -660 38600 -650
rect 37680 -680 37690 -660
rect 37570 -710 37690 -680
rect 37680 -720 37690 -710
rect 37750 -720 37760 -660
rect 37680 -730 37760 -720
rect 38520 -720 38530 -660
rect 38590 -680 38600 -660
rect 38590 -710 38720 -680
rect 38590 -720 38600 -710
rect 38520 -730 38600 -720
rect 38090 -760 38190 -740
rect 38090 -830 38110 -760
rect 38180 -830 38190 -760
rect 38090 -870 38190 -830
rect 38090 -940 38110 -870
rect 38180 -940 38190 -870
rect 38090 -950 38190 -940
rect 37680 -970 37760 -960
rect 37680 -990 37690 -970
rect 37570 -1020 37690 -990
rect 37680 -1030 37690 -1020
rect 37750 -1030 37760 -970
rect 38520 -970 38600 -960
rect 38520 -1030 38530 -970
rect 38590 -990 38600 -970
rect 38590 -1020 38720 -990
rect 38590 -1030 38600 -1020
rect 37680 -1040 37760 -1030
rect 38100 -1040 38180 -1030
rect 38520 -1040 38600 -1030
rect 38100 -1100 38110 -1040
rect 38170 -1080 38180 -1040
rect 38170 -1100 38720 -1080
rect 38100 -1110 38720 -1100
rect 38640 -1640 38720 -1630
rect 38640 -1700 38650 -1640
rect 38710 -1700 38720 -1640
rect 38640 -1710 38720 -1700
rect 38900 -1710 38930 130
rect 39020 -1710 39050 0
rect 39140 -1710 39170 0
rect 39260 -1710 39290 0
rect 39380 -1710 39410 0
rect 39500 -1710 39530 0
rect 39620 -1710 39650 0
rect 41780 -1710 41810 150
rect 41900 -1710 41930 150
rect 42020 -1710 42050 150
rect 42140 -1710 42170 150
rect 42260 -1710 42290 150
rect 42380 -1710 42410 150
rect 42500 -1710 42530 150
rect 42560 140 42640 150
rect 42560 80 42570 140
rect 42630 80 42640 140
rect 42560 70 42640 80
rect 43740 40 43860 70
rect 43630 -10 43710 0
rect 43630 -70 43640 -10
rect 43700 -70 43710 -10
rect 43740 -20 43780 40
rect 43840 -20 43860 40
rect 43740 -50 43860 -20
rect 43630 -80 43710 -70
rect 42560 -120 42640 -110
rect 42560 -180 42570 -120
rect 42630 -180 42640 -120
rect 42560 -190 42640 -180
rect 43090 -590 43710 -580
rect 43090 -650 43100 -590
rect 43160 -610 43710 -590
rect 43160 -650 43170 -610
rect 42670 -660 42750 -650
rect 43090 -660 43170 -650
rect 43510 -660 43590 -650
rect 42670 -680 42680 -660
rect 42560 -710 42680 -680
rect 42670 -720 42680 -710
rect 42740 -720 42750 -660
rect 42670 -730 42750 -720
rect 43510 -720 43520 -660
rect 43580 -680 43590 -660
rect 43580 -710 43710 -680
rect 43580 -720 43590 -710
rect 43510 -730 43590 -720
rect 43080 -760 43180 -740
rect 43080 -830 43100 -760
rect 43170 -830 43180 -760
rect 43080 -870 43180 -830
rect 43080 -940 43100 -870
rect 43170 -940 43180 -870
rect 43080 -950 43180 -940
rect 42670 -970 42750 -960
rect 42670 -990 42680 -970
rect 42560 -1020 42680 -990
rect 42670 -1030 42680 -1020
rect 42740 -1030 42750 -970
rect 43510 -970 43590 -960
rect 43510 -1030 43520 -970
rect 43580 -990 43590 -970
rect 43580 -1020 43710 -990
rect 43580 -1030 43590 -1020
rect 42670 -1040 42750 -1030
rect 43090 -1040 43170 -1030
rect 43510 -1040 43590 -1030
rect 43090 -1100 43100 -1040
rect 43160 -1080 43170 -1040
rect 43160 -1100 43710 -1080
rect 43090 -1110 43710 -1100
rect 43630 -1640 43710 -1630
rect 43630 -1700 43640 -1640
rect 43700 -1700 43710 -1640
rect 43630 -1710 43710 -1700
rect 43890 -1710 43920 130
rect 44010 -1710 44040 0
rect 44130 -1710 44160 0
rect 44250 -1710 44280 0
rect 44370 -1710 44400 0
rect 44490 -1710 44520 0
rect 44610 -1710 44640 0
rect 46770 -1710 46800 150
rect 46890 -1710 46920 150
rect 47010 -1710 47040 150
rect 47130 -1710 47160 150
rect 47250 -1710 47280 150
rect 47370 -1710 47400 150
rect 47490 -1710 47520 150
rect 47550 140 47630 150
rect 47550 80 47560 140
rect 47620 80 47630 140
rect 47550 70 47630 80
rect 48730 40 48850 70
rect 48620 -10 48700 0
rect 48620 -70 48630 -10
rect 48690 -70 48700 -10
rect 48730 -20 48770 40
rect 48830 -20 48850 40
rect 48730 -50 48850 -20
rect 48620 -80 48700 -70
rect 47550 -120 47630 -110
rect 47550 -180 47560 -120
rect 47620 -180 47630 -120
rect 47550 -190 47630 -180
rect 48080 -590 48700 -580
rect 48080 -650 48090 -590
rect 48150 -610 48700 -590
rect 48150 -650 48160 -610
rect 47660 -660 47740 -650
rect 48080 -660 48160 -650
rect 48500 -660 48580 -650
rect 47660 -680 47670 -660
rect 47550 -710 47670 -680
rect 47660 -720 47670 -710
rect 47730 -720 47740 -660
rect 47660 -730 47740 -720
rect 48500 -720 48510 -660
rect 48570 -680 48580 -660
rect 48570 -710 48700 -680
rect 48570 -720 48580 -710
rect 48500 -730 48580 -720
rect 48070 -760 48170 -740
rect 48070 -830 48090 -760
rect 48160 -830 48170 -760
rect 48070 -870 48170 -830
rect 48070 -940 48090 -870
rect 48160 -940 48170 -870
rect 48070 -950 48170 -940
rect 47660 -970 47740 -960
rect 47660 -990 47670 -970
rect 47550 -1020 47670 -990
rect 47660 -1030 47670 -1020
rect 47730 -1030 47740 -970
rect 48500 -970 48580 -960
rect 48500 -1030 48510 -970
rect 48570 -990 48580 -970
rect 48570 -1020 48700 -990
rect 48570 -1030 48580 -1020
rect 47660 -1040 47740 -1030
rect 48080 -1040 48160 -1030
rect 48500 -1040 48580 -1030
rect 48080 -1100 48090 -1040
rect 48150 -1080 48160 -1040
rect 48150 -1100 48700 -1080
rect 48080 -1110 48700 -1100
rect 48620 -1640 48700 -1630
rect 48620 -1700 48630 -1640
rect 48690 -1700 48700 -1640
rect 48620 -1710 48700 -1700
rect 48880 -1710 48910 130
rect 49000 -1710 49030 0
rect 49120 -1710 49150 0
rect 49240 -1710 49270 0
rect 49360 -1710 49390 0
rect 49480 -1710 49510 0
rect 49600 -1710 49630 0
rect 51760 -1710 51790 150
rect 51880 -1710 51910 150
rect 52000 -1710 52030 150
rect 52120 -1710 52150 150
rect 52240 -1710 52270 150
rect 52360 -1710 52390 150
rect 52480 -1710 52510 150
rect 52540 140 52620 150
rect 52540 80 52550 140
rect 52610 80 52620 140
rect 52540 70 52620 80
rect 53720 40 53840 70
rect 53610 -10 53690 0
rect 53610 -70 53620 -10
rect 53680 -70 53690 -10
rect 53720 -20 53760 40
rect 53820 -20 53840 40
rect 53720 -50 53840 -20
rect 53610 -80 53690 -70
rect 52540 -120 52620 -110
rect 52540 -180 52550 -120
rect 52610 -180 52620 -120
rect 52540 -190 52620 -180
rect 53070 -590 53690 -580
rect 53070 -650 53080 -590
rect 53140 -610 53690 -590
rect 53140 -650 53150 -610
rect 52650 -660 52730 -650
rect 53070 -660 53150 -650
rect 53490 -660 53570 -650
rect 52650 -680 52660 -660
rect 52540 -710 52660 -680
rect 52650 -720 52660 -710
rect 52720 -720 52730 -660
rect 52650 -730 52730 -720
rect 53490 -720 53500 -660
rect 53560 -680 53570 -660
rect 53560 -710 53690 -680
rect 53560 -720 53570 -710
rect 53490 -730 53570 -720
rect 53060 -760 53160 -740
rect 53060 -830 53080 -760
rect 53150 -830 53160 -760
rect 53060 -870 53160 -830
rect 53060 -940 53080 -870
rect 53150 -940 53160 -870
rect 53060 -950 53160 -940
rect 52650 -970 52730 -960
rect 52650 -990 52660 -970
rect 52540 -1020 52660 -990
rect 52650 -1030 52660 -1020
rect 52720 -1030 52730 -970
rect 53490 -970 53570 -960
rect 53490 -1030 53500 -970
rect 53560 -990 53570 -970
rect 53560 -1020 53690 -990
rect 53560 -1030 53570 -1020
rect 52650 -1040 52730 -1030
rect 53070 -1040 53150 -1030
rect 53490 -1040 53570 -1030
rect 53070 -1100 53080 -1040
rect 53140 -1080 53150 -1040
rect 53140 -1100 53690 -1080
rect 53070 -1110 53690 -1100
rect 53610 -1640 53690 -1630
rect 53610 -1700 53620 -1640
rect 53680 -1700 53690 -1640
rect 53610 -1710 53690 -1700
rect 53870 -1710 53900 130
rect 53990 -1710 54020 0
rect 54110 -1710 54140 0
rect 54230 -1710 54260 0
rect 54350 -1710 54380 0
rect 54470 -1710 54500 0
rect 54590 -1710 54620 0
rect 56750 -1710 56780 150
rect 56870 -1710 56900 150
rect 56990 -1710 57020 150
rect 57110 -1710 57140 150
rect 57230 -1710 57260 150
rect 57350 -1710 57380 150
rect 57470 -1710 57500 150
rect 57530 140 57610 150
rect 57530 80 57540 140
rect 57600 80 57610 140
rect 57530 70 57610 80
rect 58710 40 58830 70
rect 58600 -10 58680 0
rect 58600 -70 58610 -10
rect 58670 -70 58680 -10
rect 58710 -20 58750 40
rect 58810 -20 58830 40
rect 58710 -50 58830 -20
rect 58600 -80 58680 -70
rect 57530 -120 57610 -110
rect 57530 -180 57540 -120
rect 57600 -180 57610 -120
rect 57530 -190 57610 -180
rect 58060 -590 58680 -580
rect 58060 -650 58070 -590
rect 58130 -610 58680 -590
rect 58130 -650 58140 -610
rect 57640 -660 57720 -650
rect 58060 -660 58140 -650
rect 58480 -660 58560 -650
rect 57640 -680 57650 -660
rect 57530 -710 57650 -680
rect 57640 -720 57650 -710
rect 57710 -720 57720 -660
rect 57640 -730 57720 -720
rect 58480 -720 58490 -660
rect 58550 -680 58560 -660
rect 58550 -710 58680 -680
rect 58550 -720 58560 -710
rect 58480 -730 58560 -720
rect 58050 -760 58150 -740
rect 58050 -830 58070 -760
rect 58140 -830 58150 -760
rect 58050 -870 58150 -830
rect 58050 -940 58070 -870
rect 58140 -940 58150 -870
rect 58050 -950 58150 -940
rect 57640 -970 57720 -960
rect 57640 -990 57650 -970
rect 57530 -1020 57650 -990
rect 57640 -1030 57650 -1020
rect 57710 -1030 57720 -970
rect 58480 -970 58560 -960
rect 58480 -1030 58490 -970
rect 58550 -990 58560 -970
rect 58550 -1020 58680 -990
rect 58550 -1030 58560 -1020
rect 57640 -1040 57720 -1030
rect 58060 -1040 58140 -1030
rect 58480 -1040 58560 -1030
rect 58060 -1100 58070 -1040
rect 58130 -1080 58140 -1040
rect 58130 -1100 58680 -1080
rect 58060 -1110 58680 -1100
rect 58600 -1640 58680 -1630
rect 58600 -1700 58610 -1640
rect 58670 -1700 58680 -1640
rect 58600 -1710 58680 -1700
rect 58860 -1710 58890 130
rect 58980 -1710 59010 0
rect 59100 -1710 59130 0
rect 59220 -1710 59250 0
rect 59340 -1710 59370 0
rect 59460 -1710 59490 0
rect 59580 -1710 59610 0
rect 61740 -1710 61770 150
rect 61860 -1710 61890 150
rect 61980 -1710 62010 150
rect 62100 -1710 62130 150
rect 62220 -1710 62250 150
rect 62340 -1710 62370 150
rect 62460 -1710 62490 150
rect 62520 140 62600 150
rect 62520 80 62530 140
rect 62590 80 62600 140
rect 62520 70 62600 80
rect 63700 40 63820 70
rect 63590 -10 63670 0
rect 63590 -70 63600 -10
rect 63660 -70 63670 -10
rect 63700 -20 63740 40
rect 63800 -20 63820 40
rect 63700 -50 63820 -20
rect 63590 -80 63670 -70
rect 62520 -120 62600 -110
rect 62520 -180 62530 -120
rect 62590 -180 62600 -120
rect 62520 -190 62600 -180
rect 63050 -590 63670 -580
rect 63050 -650 63060 -590
rect 63120 -610 63670 -590
rect 63120 -650 63130 -610
rect 62630 -660 62710 -650
rect 63050 -660 63130 -650
rect 63470 -660 63550 -650
rect 62630 -680 62640 -660
rect 62520 -710 62640 -680
rect 62630 -720 62640 -710
rect 62700 -720 62710 -660
rect 62630 -730 62710 -720
rect 63470 -720 63480 -660
rect 63540 -680 63550 -660
rect 63540 -710 63670 -680
rect 63540 -720 63550 -710
rect 63470 -730 63550 -720
rect 63040 -760 63140 -740
rect 63040 -830 63060 -760
rect 63130 -830 63140 -760
rect 63040 -870 63140 -830
rect 63040 -940 63060 -870
rect 63130 -940 63140 -870
rect 63040 -950 63140 -940
rect 62630 -970 62710 -960
rect 62630 -990 62640 -970
rect 62520 -1020 62640 -990
rect 62630 -1030 62640 -1020
rect 62700 -1030 62710 -970
rect 63470 -970 63550 -960
rect 63470 -1030 63480 -970
rect 63540 -990 63550 -970
rect 63540 -1020 63670 -990
rect 63540 -1030 63550 -1020
rect 62630 -1040 62710 -1030
rect 63050 -1040 63130 -1030
rect 63470 -1040 63550 -1030
rect 63050 -1100 63060 -1040
rect 63120 -1080 63130 -1040
rect 63120 -1100 63670 -1080
rect 63050 -1110 63670 -1100
rect 63590 -1640 63670 -1630
rect 63590 -1700 63600 -1640
rect 63660 -1700 63670 -1640
rect 63590 -1710 63670 -1700
rect 63850 -1710 63880 130
rect 63970 -1710 64000 0
rect 64090 -1710 64120 0
rect 64210 -1710 64240 0
rect 64330 -1710 64360 0
rect 64450 -1710 64480 0
rect 64570 -1710 64600 0
rect 66730 -1710 66760 150
rect 66850 -1710 66880 150
rect 66970 -1710 67000 150
rect 67090 -1710 67120 150
rect 67210 -1710 67240 150
rect 67330 -1710 67360 150
rect 67450 -1710 67480 150
rect 67510 140 67590 150
rect 67510 80 67520 140
rect 67580 80 67590 140
rect 67510 70 67590 80
rect 68690 40 68810 70
rect 68580 -10 68660 0
rect 68580 -70 68590 -10
rect 68650 -70 68660 -10
rect 68690 -20 68730 40
rect 68790 -20 68810 40
rect 68690 -50 68810 -20
rect 68580 -80 68660 -70
rect 67510 -120 67590 -110
rect 67510 -180 67520 -120
rect 67580 -180 67590 -120
rect 67510 -190 67590 -180
rect 68040 -590 68660 -580
rect 68040 -650 68050 -590
rect 68110 -610 68660 -590
rect 68110 -650 68120 -610
rect 67620 -660 67700 -650
rect 68040 -660 68120 -650
rect 68460 -660 68540 -650
rect 67620 -680 67630 -660
rect 67510 -710 67630 -680
rect 67620 -720 67630 -710
rect 67690 -720 67700 -660
rect 67620 -730 67700 -720
rect 68460 -720 68470 -660
rect 68530 -680 68540 -660
rect 68530 -710 68660 -680
rect 68530 -720 68540 -710
rect 68460 -730 68540 -720
rect 68030 -760 68130 -740
rect 68030 -830 68050 -760
rect 68120 -830 68130 -760
rect 68030 -870 68130 -830
rect 68030 -940 68050 -870
rect 68120 -940 68130 -870
rect 68030 -950 68130 -940
rect 67620 -970 67700 -960
rect 67620 -990 67630 -970
rect 67510 -1020 67630 -990
rect 67620 -1030 67630 -1020
rect 67690 -1030 67700 -970
rect 68460 -970 68540 -960
rect 68460 -1030 68470 -970
rect 68530 -990 68540 -970
rect 68530 -1020 68660 -990
rect 68530 -1030 68540 -1020
rect 67620 -1040 67700 -1030
rect 68040 -1040 68120 -1030
rect 68460 -1040 68540 -1030
rect 68040 -1100 68050 -1040
rect 68110 -1080 68120 -1040
rect 68110 -1100 68660 -1080
rect 68040 -1110 68660 -1100
rect 68580 -1640 68660 -1630
rect 68580 -1700 68590 -1640
rect 68650 -1700 68660 -1640
rect 68580 -1710 68660 -1700
rect 68840 -1710 68870 130
rect 68960 -1710 68990 0
rect 69080 -1710 69110 0
rect 69200 -1710 69230 0
rect 69320 -1710 69350 0
rect 69440 -1710 69470 0
rect 69560 -1710 69590 0
rect 71720 -1710 71750 150
rect 71840 -1710 71870 150
rect 71960 -1710 71990 150
rect 72080 -1710 72110 150
rect 72200 -1710 72230 150
rect 72320 -1710 72350 150
rect 72440 -1710 72470 150
rect 72500 140 72580 150
rect 72500 80 72510 140
rect 72570 80 72580 140
rect 72500 70 72580 80
rect 73680 40 73800 70
rect 73570 -10 73650 0
rect 73570 -70 73580 -10
rect 73640 -70 73650 -10
rect 73680 -20 73720 40
rect 73780 -20 73800 40
rect 73680 -50 73800 -20
rect 73570 -80 73650 -70
rect 72500 -120 72580 -110
rect 72500 -180 72510 -120
rect 72570 -180 72580 -120
rect 72500 -190 72580 -180
rect 73030 -590 73650 -580
rect 73030 -650 73040 -590
rect 73100 -610 73650 -590
rect 73100 -650 73110 -610
rect 72610 -660 72690 -650
rect 73030 -660 73110 -650
rect 73450 -660 73530 -650
rect 72610 -680 72620 -660
rect 72500 -710 72620 -680
rect 72610 -720 72620 -710
rect 72680 -720 72690 -660
rect 72610 -730 72690 -720
rect 73450 -720 73460 -660
rect 73520 -680 73530 -660
rect 73520 -710 73650 -680
rect 73520 -720 73530 -710
rect 73450 -730 73530 -720
rect 73020 -760 73120 -740
rect 73020 -830 73040 -760
rect 73110 -830 73120 -760
rect 73020 -870 73120 -830
rect 73020 -940 73040 -870
rect 73110 -940 73120 -870
rect 73020 -950 73120 -940
rect 72610 -970 72690 -960
rect 72610 -990 72620 -970
rect 72500 -1020 72620 -990
rect 72610 -1030 72620 -1020
rect 72680 -1030 72690 -970
rect 73450 -970 73530 -960
rect 73450 -1030 73460 -970
rect 73520 -990 73530 -970
rect 73520 -1020 73650 -990
rect 73520 -1030 73530 -1020
rect 72610 -1040 72690 -1030
rect 73030 -1040 73110 -1030
rect 73450 -1040 73530 -1030
rect 73030 -1100 73040 -1040
rect 73100 -1080 73110 -1040
rect 73100 -1100 73650 -1080
rect 73030 -1110 73650 -1100
rect 73570 -1640 73650 -1630
rect 73570 -1700 73580 -1640
rect 73640 -1700 73650 -1640
rect 73570 -1710 73650 -1700
rect 73830 -1710 73860 130
rect 73950 -1710 73980 0
rect 74070 -1710 74100 0
rect 74190 -1710 74220 0
rect 74310 -1710 74340 0
rect 74430 -1710 74460 0
rect 74550 -1710 74580 0
rect 76710 -1710 76740 150
rect 76830 -1710 76860 150
rect 76950 -1710 76980 150
rect 77070 -1710 77100 150
rect 77190 -1710 77220 150
rect 77310 -1710 77340 150
rect 77430 -1710 77460 150
rect 77490 140 77570 150
rect 77490 80 77500 140
rect 77560 80 77570 140
rect 77490 70 77570 80
rect 78560 -10 78640 0
rect 78560 -70 78570 -10
rect 78630 -70 78640 -10
rect 78560 -80 78640 -70
rect 77490 -120 77570 -110
rect 77490 -180 77500 -120
rect 77560 -180 77570 -120
rect 77490 -190 77570 -180
rect 78020 -590 78640 -580
rect 78020 -650 78030 -590
rect 78090 -610 78640 -590
rect 78090 -650 78100 -610
rect 77600 -660 77680 -650
rect 78020 -660 78100 -650
rect 78440 -660 78520 -650
rect 77600 -680 77610 -660
rect 77490 -710 77610 -680
rect 77600 -720 77610 -710
rect 77670 -720 77680 -660
rect 77600 -730 77680 -720
rect 78440 -720 78450 -660
rect 78510 -680 78520 -660
rect 78510 -710 78640 -680
rect 78510 -720 78520 -710
rect 78440 -730 78520 -720
rect 78010 -760 78110 -740
rect 78010 -830 78030 -760
rect 78100 -830 78110 -760
rect 78010 -870 78110 -830
rect 78010 -940 78030 -870
rect 78100 -940 78110 -870
rect 78010 -950 78110 -940
rect 77600 -970 77680 -960
rect 77600 -990 77610 -970
rect 77490 -1020 77610 -990
rect 77600 -1030 77610 -1020
rect 77670 -1030 77680 -970
rect 78440 -970 78520 -960
rect 78440 -1030 78450 -970
rect 78510 -990 78520 -970
rect 78510 -1020 78640 -990
rect 78510 -1030 78520 -1020
rect 77600 -1040 77680 -1030
rect 78020 -1040 78100 -1030
rect 78440 -1040 78520 -1030
rect 78020 -1100 78030 -1040
rect 78090 -1080 78100 -1040
rect 78090 -1100 78640 -1080
rect 78020 -1110 78640 -1100
rect 78560 -1640 78640 -1630
rect 78560 -1700 78570 -1640
rect 78630 -1700 78640 -1640
rect 78560 -1710 78640 -1700
rect 78820 -1710 78850 -260
rect 78940 -1710 78970 -260
rect 79060 -1710 79090 -260
rect 79180 -1710 79210 -260
rect 79300 -1710 79330 -260
rect 79420 -1710 79450 -260
rect 79540 -1710 79570 -260
rect 81430 -1710 81460 29070
rect 81550 -1710 81580 29070
rect 81670 -1710 81700 29070
rect 81790 -1710 81820 29070
rect 81910 -1710 81940 29070
rect 82030 -1710 82060 29070
rect 82150 -1710 82180 29070
rect 83280 29060 83360 29070
rect 83280 29000 83290 29060
rect 83350 29000 83360 29060
rect 83280 28990 83360 29000
rect 82210 28950 82290 28960
rect 82210 28890 82220 28950
rect 82280 28890 82290 28950
rect 82210 28880 82290 28890
rect 82740 28480 83360 28490
rect 82740 28420 82750 28480
rect 82810 28460 83360 28480
rect 82810 28420 82820 28460
rect 82320 28410 82400 28420
rect 82740 28410 82820 28420
rect 83160 28410 83240 28420
rect 82320 28390 82330 28410
rect 82210 28360 82330 28390
rect 82320 28350 82330 28360
rect 82390 28350 82400 28410
rect 82320 28340 82400 28350
rect 83160 28350 83170 28410
rect 83230 28390 83240 28410
rect 83230 28360 83360 28390
rect 83230 28350 83240 28360
rect 83160 28340 83240 28350
rect 82730 28310 82830 28330
rect 82730 28240 82750 28310
rect 82820 28240 82830 28310
rect 82730 28200 82830 28240
rect 82730 28130 82750 28200
rect 82820 28130 82830 28200
rect 82730 28120 82830 28130
rect 82320 28100 82400 28110
rect 82320 28080 82330 28100
rect 82210 28050 82330 28080
rect 82320 28040 82330 28050
rect 82390 28040 82400 28100
rect 83160 28100 83240 28110
rect 83160 28040 83170 28100
rect 83230 28080 83240 28100
rect 83230 28050 83360 28080
rect 83230 28040 83240 28050
rect 82320 28030 82400 28040
rect 82740 28030 82820 28040
rect 83160 28030 83240 28040
rect 82740 27970 82750 28030
rect 82810 27990 82820 28030
rect 82810 27970 83360 27990
rect 82740 27960 83360 27970
rect 83270 27490 83360 27500
rect 83270 27430 83280 27490
rect 83350 27430 83360 27490
rect 83270 27420 83360 27430
rect 83280 27350 83360 27360
rect 83280 27290 83290 27350
rect 83350 27290 83360 27350
rect 83280 27280 83360 27290
rect 82210 27240 82290 27250
rect 82210 27180 82220 27240
rect 82280 27180 82290 27240
rect 82210 27170 82290 27180
rect 82740 26770 83360 26780
rect 82740 26710 82750 26770
rect 82810 26750 83360 26770
rect 82810 26710 82820 26750
rect 82320 26700 82400 26710
rect 82740 26700 82820 26710
rect 83160 26700 83240 26710
rect 82320 26680 82330 26700
rect 82210 26650 82330 26680
rect 82320 26640 82330 26650
rect 82390 26640 82400 26700
rect 82320 26630 82400 26640
rect 83160 26640 83170 26700
rect 83230 26680 83240 26700
rect 83230 26650 83360 26680
rect 83230 26640 83240 26650
rect 83160 26630 83240 26640
rect 82730 26600 82830 26620
rect 82730 26530 82750 26600
rect 82820 26530 82830 26600
rect 82730 26490 82830 26530
rect 82730 26420 82750 26490
rect 82820 26420 82830 26490
rect 82730 26410 82830 26420
rect 82320 26390 82400 26400
rect 82320 26370 82330 26390
rect 82210 26340 82330 26370
rect 82320 26330 82330 26340
rect 82390 26330 82400 26390
rect 83160 26390 83240 26400
rect 83160 26330 83170 26390
rect 83230 26370 83240 26390
rect 83230 26340 83360 26370
rect 83230 26330 83240 26340
rect 82320 26320 82400 26330
rect 82740 26320 82820 26330
rect 83160 26320 83240 26330
rect 82740 26260 82750 26320
rect 82810 26280 82820 26320
rect 82810 26260 83360 26280
rect 82740 26250 83360 26260
rect 83270 25780 83360 25790
rect 83270 25720 83280 25780
rect 83350 25720 83360 25780
rect 83270 25710 83360 25720
rect 83280 25640 83360 25650
rect 83280 25580 83290 25640
rect 83350 25580 83360 25640
rect 83280 25570 83360 25580
rect 82210 25530 82290 25540
rect 82210 25470 82220 25530
rect 82280 25470 82290 25530
rect 82210 25460 82290 25470
rect 82740 25060 83360 25070
rect 82740 25000 82750 25060
rect 82810 25040 83360 25060
rect 82810 25000 82820 25040
rect 82320 24990 82400 25000
rect 82740 24990 82820 25000
rect 83160 24990 83240 25000
rect 82320 24970 82330 24990
rect 82210 24940 82330 24970
rect 82320 24930 82330 24940
rect 82390 24930 82400 24990
rect 82320 24920 82400 24930
rect 83160 24930 83170 24990
rect 83230 24970 83240 24990
rect 83230 24940 83360 24970
rect 83230 24930 83240 24940
rect 83160 24920 83240 24930
rect 82730 24890 82830 24910
rect 82730 24820 82750 24890
rect 82820 24820 82830 24890
rect 82730 24780 82830 24820
rect 82730 24710 82750 24780
rect 82820 24710 82830 24780
rect 82730 24700 82830 24710
rect 82320 24680 82400 24690
rect 82320 24660 82330 24680
rect 82210 24630 82330 24660
rect 82320 24620 82330 24630
rect 82390 24620 82400 24680
rect 83160 24680 83240 24690
rect 83160 24620 83170 24680
rect 83230 24660 83240 24680
rect 83230 24630 83360 24660
rect 83230 24620 83240 24630
rect 82320 24610 82400 24620
rect 82740 24610 82820 24620
rect 83160 24610 83240 24620
rect 82740 24550 82750 24610
rect 82810 24570 82820 24610
rect 82810 24550 83360 24570
rect 82740 24540 83360 24550
rect 83270 24070 83360 24080
rect 83270 24010 83280 24070
rect 83350 24010 83360 24070
rect 83270 24000 83360 24010
rect 83280 23930 83360 23940
rect 83280 23870 83290 23930
rect 83350 23870 83360 23930
rect 83280 23860 83360 23870
rect 82210 23820 82290 23830
rect 82210 23760 82220 23820
rect 82280 23760 82290 23820
rect 82210 23750 82290 23760
rect 82740 23350 83360 23360
rect 82740 23290 82750 23350
rect 82810 23330 83360 23350
rect 82810 23290 82820 23330
rect 82320 23280 82400 23290
rect 82740 23280 82820 23290
rect 83160 23280 83240 23290
rect 82320 23260 82330 23280
rect 82210 23230 82330 23260
rect 82320 23220 82330 23230
rect 82390 23220 82400 23280
rect 82320 23210 82400 23220
rect 83160 23220 83170 23280
rect 83230 23260 83240 23280
rect 83230 23230 83360 23260
rect 83230 23220 83240 23230
rect 83160 23210 83240 23220
rect 82730 23180 82830 23200
rect 82730 23110 82750 23180
rect 82820 23110 82830 23180
rect 82730 23070 82830 23110
rect 82730 23000 82750 23070
rect 82820 23000 82830 23070
rect 82730 22990 82830 23000
rect 82320 22970 82400 22980
rect 82320 22950 82330 22970
rect 82210 22920 82330 22950
rect 82320 22910 82330 22920
rect 82390 22910 82400 22970
rect 83160 22970 83240 22980
rect 83160 22910 83170 22970
rect 83230 22950 83240 22970
rect 83230 22920 83360 22950
rect 83230 22910 83240 22920
rect 82320 22900 82400 22910
rect 82740 22900 82820 22910
rect 83160 22900 83240 22910
rect 82740 22840 82750 22900
rect 82810 22860 82820 22900
rect 82810 22840 83360 22860
rect 82740 22830 83360 22840
rect 83270 22360 83360 22370
rect 83270 22300 83280 22360
rect 83350 22300 83360 22360
rect 83270 22290 83360 22300
rect 83280 22220 83360 22230
rect 83280 22160 83290 22220
rect 83350 22160 83360 22220
rect 83280 22150 83360 22160
rect 82210 22110 82290 22120
rect 82210 22050 82220 22110
rect 82280 22050 82290 22110
rect 82210 22040 82290 22050
rect 82740 21640 83360 21650
rect 82740 21580 82750 21640
rect 82810 21620 83360 21640
rect 82810 21580 82820 21620
rect 82320 21570 82400 21580
rect 82740 21570 82820 21580
rect 83160 21570 83240 21580
rect 82320 21550 82330 21570
rect 82210 21520 82330 21550
rect 82320 21510 82330 21520
rect 82390 21510 82400 21570
rect 82320 21500 82400 21510
rect 83160 21510 83170 21570
rect 83230 21550 83240 21570
rect 83230 21520 83360 21550
rect 83230 21510 83240 21520
rect 83160 21500 83240 21510
rect 82730 21470 82830 21490
rect 82730 21400 82750 21470
rect 82820 21400 82830 21470
rect 82730 21360 82830 21400
rect 82730 21290 82750 21360
rect 82820 21290 82830 21360
rect 82730 21280 82830 21290
rect 82320 21260 82400 21270
rect 82320 21240 82330 21260
rect 82210 21210 82330 21240
rect 82320 21200 82330 21210
rect 82390 21200 82400 21260
rect 83160 21260 83240 21270
rect 83160 21200 83170 21260
rect 83230 21240 83240 21260
rect 83230 21210 83360 21240
rect 83230 21200 83240 21210
rect 82320 21190 82400 21200
rect 82740 21190 82820 21200
rect 83160 21190 83240 21200
rect 82740 21130 82750 21190
rect 82810 21150 82820 21190
rect 82810 21130 83360 21150
rect 82740 21120 83360 21130
rect 83270 20650 83360 20660
rect 83270 20590 83280 20650
rect 83350 20590 83360 20650
rect 83270 20580 83360 20590
rect 83280 20510 83360 20520
rect 83280 20450 83290 20510
rect 83350 20450 83360 20510
rect 83280 20440 83360 20450
rect 82210 20400 82290 20410
rect 82210 20340 82220 20400
rect 82280 20340 82290 20400
rect 82210 20330 82290 20340
rect 82740 19930 83360 19940
rect 82740 19870 82750 19930
rect 82810 19910 83360 19930
rect 82810 19870 82820 19910
rect 82320 19860 82400 19870
rect 82740 19860 82820 19870
rect 83160 19860 83240 19870
rect 82320 19840 82330 19860
rect 82210 19810 82330 19840
rect 82320 19800 82330 19810
rect 82390 19800 82400 19860
rect 82320 19790 82400 19800
rect 83160 19800 83170 19860
rect 83230 19840 83240 19860
rect 83230 19810 83360 19840
rect 83230 19800 83240 19810
rect 83160 19790 83240 19800
rect 82730 19760 82830 19780
rect 82730 19690 82750 19760
rect 82820 19690 82830 19760
rect 82730 19650 82830 19690
rect 82730 19580 82750 19650
rect 82820 19580 82830 19650
rect 82730 19570 82830 19580
rect 82320 19550 82400 19560
rect 82320 19530 82330 19550
rect 82210 19500 82330 19530
rect 82320 19490 82330 19500
rect 82390 19490 82400 19550
rect 83160 19550 83240 19560
rect 83160 19490 83170 19550
rect 83230 19530 83240 19550
rect 83230 19500 83360 19530
rect 83230 19490 83240 19500
rect 82320 19480 82400 19490
rect 82740 19480 82820 19490
rect 83160 19480 83240 19490
rect 82740 19420 82750 19480
rect 82810 19440 82820 19480
rect 82810 19420 83360 19440
rect 82740 19410 83360 19420
rect 83270 18940 83360 18950
rect 83270 18880 83280 18940
rect 83350 18880 83360 18940
rect 83270 18870 83360 18880
rect 83280 18800 83360 18810
rect 83280 18740 83290 18800
rect 83350 18740 83360 18800
rect 83280 18730 83360 18740
rect 82210 18690 82290 18700
rect 82210 18630 82220 18690
rect 82280 18630 82290 18690
rect 82210 18620 82290 18630
rect 82740 18220 83360 18230
rect 82740 18160 82750 18220
rect 82810 18200 83360 18220
rect 82810 18160 82820 18200
rect 82320 18150 82400 18160
rect 82740 18150 82820 18160
rect 83160 18150 83240 18160
rect 82320 18130 82330 18150
rect 82210 18100 82330 18130
rect 82320 18090 82330 18100
rect 82390 18090 82400 18150
rect 82320 18080 82400 18090
rect 83160 18090 83170 18150
rect 83230 18130 83240 18150
rect 83230 18100 83360 18130
rect 83230 18090 83240 18100
rect 83160 18080 83240 18090
rect 82730 18050 82830 18070
rect 82730 17980 82750 18050
rect 82820 17980 82830 18050
rect 82730 17940 82830 17980
rect 82730 17870 82750 17940
rect 82820 17870 82830 17940
rect 82730 17860 82830 17870
rect 82320 17840 82400 17850
rect 82320 17820 82330 17840
rect 82210 17790 82330 17820
rect 82320 17780 82330 17790
rect 82390 17780 82400 17840
rect 83160 17840 83240 17850
rect 83160 17780 83170 17840
rect 83230 17820 83240 17840
rect 83230 17790 83360 17820
rect 83230 17780 83240 17790
rect 82320 17770 82400 17780
rect 82740 17770 82820 17780
rect 83160 17770 83240 17780
rect 82740 17710 82750 17770
rect 82810 17730 82820 17770
rect 82810 17710 83360 17730
rect 82740 17700 83360 17710
rect 83270 17230 83360 17240
rect 83270 17170 83280 17230
rect 83350 17170 83360 17230
rect 83270 17160 83360 17170
rect 83280 17090 83360 17100
rect 83280 17030 83290 17090
rect 83350 17030 83360 17090
rect 83280 17020 83360 17030
rect 82210 16980 82290 16990
rect 82210 16920 82220 16980
rect 82280 16920 82290 16980
rect 82210 16910 82290 16920
rect 82740 16510 83360 16520
rect 82740 16450 82750 16510
rect 82810 16490 83360 16510
rect 82810 16450 82820 16490
rect 82320 16440 82400 16450
rect 82740 16440 82820 16450
rect 83160 16440 83240 16450
rect 82320 16420 82330 16440
rect 82210 16390 82330 16420
rect 82320 16380 82330 16390
rect 82390 16380 82400 16440
rect 82320 16370 82400 16380
rect 83160 16380 83170 16440
rect 83230 16420 83240 16440
rect 83230 16390 83360 16420
rect 83230 16380 83240 16390
rect 83160 16370 83240 16380
rect 82730 16340 82830 16360
rect 82730 16270 82750 16340
rect 82820 16270 82830 16340
rect 82730 16230 82830 16270
rect 82730 16160 82750 16230
rect 82820 16160 82830 16230
rect 82730 16150 82830 16160
rect 82320 16130 82400 16140
rect 82320 16110 82330 16130
rect 82210 16080 82330 16110
rect 82320 16070 82330 16080
rect 82390 16070 82400 16130
rect 83160 16130 83240 16140
rect 83160 16070 83170 16130
rect 83230 16110 83240 16130
rect 83230 16080 83360 16110
rect 83230 16070 83240 16080
rect 82320 16060 82400 16070
rect 82740 16060 82820 16070
rect 83160 16060 83240 16070
rect 82740 16000 82750 16060
rect 82810 16020 82820 16060
rect 82810 16000 83360 16020
rect 82740 15990 83360 16000
rect 83270 15520 83360 15530
rect 83270 15460 83280 15520
rect 83350 15460 83360 15520
rect 83270 15450 83360 15460
rect 83280 15380 83360 15390
rect 83280 15320 83290 15380
rect 83350 15320 83360 15380
rect 83280 15310 83360 15320
rect 82210 15270 82290 15280
rect 82210 15210 82220 15270
rect 82280 15210 82290 15270
rect 82210 15200 82290 15210
rect 82740 14800 83360 14810
rect 82740 14740 82750 14800
rect 82810 14780 83360 14800
rect 82810 14740 82820 14780
rect 82320 14730 82400 14740
rect 82740 14730 82820 14740
rect 83160 14730 83240 14740
rect 82320 14710 82330 14730
rect 82210 14680 82330 14710
rect 82320 14670 82330 14680
rect 82390 14670 82400 14730
rect 82320 14660 82400 14670
rect 83160 14670 83170 14730
rect 83230 14710 83240 14730
rect 83230 14680 83360 14710
rect 83230 14670 83240 14680
rect 83160 14660 83240 14670
rect 82730 14630 82830 14650
rect 82730 14560 82750 14630
rect 82820 14560 82830 14630
rect 82730 14520 82830 14560
rect 82730 14450 82750 14520
rect 82820 14450 82830 14520
rect 82730 14440 82830 14450
rect 82320 14420 82400 14430
rect 82320 14400 82330 14420
rect 82210 14370 82330 14400
rect 82320 14360 82330 14370
rect 82390 14360 82400 14420
rect 83160 14420 83240 14430
rect 83160 14360 83170 14420
rect 83230 14400 83240 14420
rect 83230 14370 83360 14400
rect 83230 14360 83240 14370
rect 82320 14350 82400 14360
rect 82740 14350 82820 14360
rect 83160 14350 83240 14360
rect 82740 14290 82750 14350
rect 82810 14310 82820 14350
rect 82810 14290 83360 14310
rect 82740 14280 83360 14290
rect 83270 13810 83360 13820
rect 83270 13750 83280 13810
rect 83350 13750 83360 13810
rect 83270 13740 83360 13750
rect 83280 13670 83360 13680
rect 83280 13610 83290 13670
rect 83350 13610 83360 13670
rect 83280 13600 83360 13610
rect 82210 13560 82290 13570
rect 82210 13500 82220 13560
rect 82280 13500 82290 13560
rect 82210 13490 82290 13500
rect 82740 13090 83360 13100
rect 82740 13030 82750 13090
rect 82810 13070 83360 13090
rect 82810 13030 82820 13070
rect 82320 13020 82400 13030
rect 82740 13020 82820 13030
rect 83160 13020 83240 13030
rect 82320 13000 82330 13020
rect 82210 12970 82330 13000
rect 82320 12960 82330 12970
rect 82390 12960 82400 13020
rect 82320 12950 82400 12960
rect 83160 12960 83170 13020
rect 83230 13000 83240 13020
rect 83230 12970 83360 13000
rect 83230 12960 83240 12970
rect 83160 12950 83240 12960
rect 82730 12920 82830 12940
rect 82730 12850 82750 12920
rect 82820 12850 82830 12920
rect 82730 12810 82830 12850
rect 82730 12740 82750 12810
rect 82820 12740 82830 12810
rect 82730 12730 82830 12740
rect 82320 12710 82400 12720
rect 82320 12690 82330 12710
rect 82210 12660 82330 12690
rect 82320 12650 82330 12660
rect 82390 12650 82400 12710
rect 83160 12710 83240 12720
rect 83160 12650 83170 12710
rect 83230 12690 83240 12710
rect 83230 12660 83360 12690
rect 83230 12650 83240 12660
rect 82320 12640 82400 12650
rect 82740 12640 82820 12650
rect 83160 12640 83240 12650
rect 82740 12580 82750 12640
rect 82810 12600 82820 12640
rect 82810 12580 83360 12600
rect 82740 12570 83360 12580
rect 83270 12100 83360 12110
rect 83270 12040 83280 12100
rect 83350 12040 83360 12100
rect 83270 12030 83360 12040
rect 83280 11960 83360 11970
rect 83280 11900 83290 11960
rect 83350 11900 83360 11960
rect 83280 11890 83360 11900
rect 82210 11850 82290 11860
rect 82210 11790 82220 11850
rect 82280 11790 82290 11850
rect 82210 11780 82290 11790
rect 82740 11380 83360 11390
rect 82740 11320 82750 11380
rect 82810 11360 83360 11380
rect 82810 11320 82820 11360
rect 82320 11310 82400 11320
rect 82740 11310 82820 11320
rect 83160 11310 83240 11320
rect 82320 11290 82330 11310
rect 82210 11260 82330 11290
rect 82320 11250 82330 11260
rect 82390 11250 82400 11310
rect 82320 11240 82400 11250
rect 83160 11250 83170 11310
rect 83230 11290 83240 11310
rect 83230 11260 83360 11290
rect 83230 11250 83240 11260
rect 83160 11240 83240 11250
rect 82730 11210 82830 11230
rect 82730 11140 82750 11210
rect 82820 11140 82830 11210
rect 82730 11100 82830 11140
rect 82730 11030 82750 11100
rect 82820 11030 82830 11100
rect 82730 11020 82830 11030
rect 82320 11000 82400 11010
rect 82320 10980 82330 11000
rect 82210 10950 82330 10980
rect 82320 10940 82330 10950
rect 82390 10940 82400 11000
rect 83160 11000 83240 11010
rect 83160 10940 83170 11000
rect 83230 10980 83240 11000
rect 83230 10950 83360 10980
rect 83230 10940 83240 10950
rect 82320 10930 82400 10940
rect 82740 10930 82820 10940
rect 83160 10930 83240 10940
rect 82740 10870 82750 10930
rect 82810 10890 82820 10930
rect 82810 10870 83360 10890
rect 82740 10860 83360 10870
rect 83270 10390 83360 10400
rect 83270 10330 83280 10390
rect 83350 10330 83360 10390
rect 83270 10320 83360 10330
rect 83280 10250 83360 10260
rect 83280 10190 83290 10250
rect 83350 10190 83360 10250
rect 83280 10180 83360 10190
rect 82210 10140 82290 10150
rect 82210 10080 82220 10140
rect 82280 10080 82290 10140
rect 82210 10070 82290 10080
rect 82740 9670 83360 9680
rect 82740 9610 82750 9670
rect 82810 9650 83360 9670
rect 82810 9610 82820 9650
rect 82320 9600 82400 9610
rect 82740 9600 82820 9610
rect 83160 9600 83240 9610
rect 82320 9580 82330 9600
rect 82210 9550 82330 9580
rect 82320 9540 82330 9550
rect 82390 9540 82400 9600
rect 82320 9530 82400 9540
rect 83160 9540 83170 9600
rect 83230 9580 83240 9600
rect 83230 9550 83360 9580
rect 83230 9540 83240 9550
rect 83160 9530 83240 9540
rect 82730 9500 82830 9520
rect 82730 9430 82750 9500
rect 82820 9430 82830 9500
rect 82730 9390 82830 9430
rect 82730 9320 82750 9390
rect 82820 9320 82830 9390
rect 82730 9310 82830 9320
rect 82320 9290 82400 9300
rect 82320 9270 82330 9290
rect 82210 9240 82330 9270
rect 82320 9230 82330 9240
rect 82390 9230 82400 9290
rect 83160 9290 83240 9300
rect 83160 9230 83170 9290
rect 83230 9270 83240 9290
rect 83230 9240 83360 9270
rect 83230 9230 83240 9240
rect 82320 9220 82400 9230
rect 82740 9220 82820 9230
rect 83160 9220 83240 9230
rect 82740 9160 82750 9220
rect 82810 9180 82820 9220
rect 82810 9160 83360 9180
rect 82740 9150 83360 9160
rect 83270 8680 83360 8690
rect 83270 8620 83280 8680
rect 83350 8620 83360 8680
rect 83270 8610 83360 8620
rect 83280 8540 83360 8550
rect 83280 8480 83290 8540
rect 83350 8480 83360 8540
rect 83280 8470 83360 8480
rect 82210 8430 82290 8440
rect 82210 8370 82220 8430
rect 82280 8370 82290 8430
rect 82210 8360 82290 8370
rect 82740 7960 83360 7970
rect 82740 7900 82750 7960
rect 82810 7940 83360 7960
rect 82810 7900 82820 7940
rect 82320 7890 82400 7900
rect 82740 7890 82820 7900
rect 83160 7890 83240 7900
rect 82320 7870 82330 7890
rect 82210 7840 82330 7870
rect 82320 7830 82330 7840
rect 82390 7830 82400 7890
rect 82320 7820 82400 7830
rect 83160 7830 83170 7890
rect 83230 7870 83240 7890
rect 83230 7840 83360 7870
rect 83230 7830 83240 7840
rect 83160 7820 83240 7830
rect 82730 7790 82830 7810
rect 82730 7720 82750 7790
rect 82820 7720 82830 7790
rect 82730 7680 82830 7720
rect 82730 7610 82750 7680
rect 82820 7610 82830 7680
rect 82730 7600 82830 7610
rect 82320 7580 82400 7590
rect 82320 7560 82330 7580
rect 82210 7530 82330 7560
rect 82320 7520 82330 7530
rect 82390 7520 82400 7580
rect 83160 7580 83240 7590
rect 83160 7520 83170 7580
rect 83230 7560 83240 7580
rect 83230 7530 83360 7560
rect 83230 7520 83240 7530
rect 82320 7510 82400 7520
rect 82740 7510 82820 7520
rect 83160 7510 83240 7520
rect 82740 7450 82750 7510
rect 82810 7470 82820 7510
rect 82810 7450 83360 7470
rect 82740 7440 83360 7450
rect 83270 6970 83360 6980
rect 83270 6910 83280 6970
rect 83350 6910 83360 6970
rect 83270 6900 83360 6910
rect 83280 6830 83360 6840
rect 83280 6770 83290 6830
rect 83350 6770 83360 6830
rect 83280 6760 83360 6770
rect 82210 6720 82290 6730
rect 82210 6660 82220 6720
rect 82280 6660 82290 6720
rect 82210 6650 82290 6660
rect 82740 6250 83360 6260
rect 82740 6190 82750 6250
rect 82810 6230 83360 6250
rect 82810 6190 82820 6230
rect 82320 6180 82400 6190
rect 82740 6180 82820 6190
rect 83160 6180 83240 6190
rect 82320 6160 82330 6180
rect 82210 6130 82330 6160
rect 82320 6120 82330 6130
rect 82390 6120 82400 6180
rect 82320 6110 82400 6120
rect 83160 6120 83170 6180
rect 83230 6160 83240 6180
rect 83230 6130 83360 6160
rect 83230 6120 83240 6130
rect 83160 6110 83240 6120
rect 82730 6080 82830 6100
rect 82730 6010 82750 6080
rect 82820 6010 82830 6080
rect 82730 5970 82830 6010
rect 82730 5900 82750 5970
rect 82820 5900 82830 5970
rect 82730 5890 82830 5900
rect 82320 5870 82400 5880
rect 82320 5850 82330 5870
rect 82210 5820 82330 5850
rect 82320 5810 82330 5820
rect 82390 5810 82400 5870
rect 83160 5870 83240 5880
rect 83160 5810 83170 5870
rect 83230 5850 83240 5870
rect 83230 5820 83360 5850
rect 83230 5810 83240 5820
rect 82320 5800 82400 5810
rect 82740 5800 82820 5810
rect 83160 5800 83240 5810
rect 82740 5740 82750 5800
rect 82810 5760 82820 5800
rect 82810 5740 83360 5760
rect 82740 5730 83360 5740
rect 83270 5260 83360 5270
rect 83270 5200 83280 5260
rect 83350 5200 83360 5260
rect 83270 5190 83360 5200
rect 83280 5120 83360 5130
rect 83280 5060 83290 5120
rect 83350 5060 83360 5120
rect 83280 5050 83360 5060
rect 82210 5010 82290 5020
rect 82210 4950 82220 5010
rect 82280 4950 82290 5010
rect 82210 4940 82290 4950
rect 82740 4540 83360 4550
rect 82740 4480 82750 4540
rect 82810 4520 83360 4540
rect 82810 4480 82820 4520
rect 82320 4470 82400 4480
rect 82740 4470 82820 4480
rect 83160 4470 83240 4480
rect 82320 4450 82330 4470
rect 82210 4420 82330 4450
rect 82320 4410 82330 4420
rect 82390 4410 82400 4470
rect 82320 4400 82400 4410
rect 83160 4410 83170 4470
rect 83230 4450 83240 4470
rect 83230 4420 83360 4450
rect 83230 4410 83240 4420
rect 83160 4400 83240 4410
rect 82730 4370 82830 4390
rect 82730 4300 82750 4370
rect 82820 4300 82830 4370
rect 82730 4260 82830 4300
rect 82730 4190 82750 4260
rect 82820 4190 82830 4260
rect 82730 4180 82830 4190
rect 82320 4160 82400 4170
rect 82320 4140 82330 4160
rect 82210 4110 82330 4140
rect 82320 4100 82330 4110
rect 82390 4100 82400 4160
rect 83160 4160 83240 4170
rect 83160 4100 83170 4160
rect 83230 4140 83240 4160
rect 83230 4110 83360 4140
rect 83230 4100 83240 4110
rect 82320 4090 82400 4100
rect 82740 4090 82820 4100
rect 83160 4090 83240 4100
rect 82740 4030 82750 4090
rect 82810 4050 82820 4090
rect 82810 4030 83360 4050
rect 82740 4020 83360 4030
rect 83270 3550 83360 3560
rect 83270 3490 83280 3550
rect 83350 3490 83360 3550
rect 83270 3480 83360 3490
rect 83280 3410 83360 3420
rect 83280 3350 83290 3410
rect 83350 3350 83360 3410
rect 83280 3340 83360 3350
rect 82210 3300 82290 3310
rect 82210 3240 82220 3300
rect 82280 3240 82290 3300
rect 82210 3230 82290 3240
rect 82740 2830 83360 2840
rect 82740 2770 82750 2830
rect 82810 2810 83360 2830
rect 82810 2770 82820 2810
rect 82320 2760 82400 2770
rect 82740 2760 82820 2770
rect 83160 2760 83240 2770
rect 82320 2740 82330 2760
rect 82210 2710 82330 2740
rect 82320 2700 82330 2710
rect 82390 2700 82400 2760
rect 82320 2690 82400 2700
rect 83160 2700 83170 2760
rect 83230 2740 83240 2760
rect 83230 2710 83360 2740
rect 83230 2700 83240 2710
rect 83160 2690 83240 2700
rect 82730 2660 82830 2680
rect 82730 2590 82750 2660
rect 82820 2590 82830 2660
rect 82730 2550 82830 2590
rect 82730 2480 82750 2550
rect 82820 2480 82830 2550
rect 82730 2470 82830 2480
rect 82320 2450 82400 2460
rect 82320 2430 82330 2450
rect 82210 2400 82330 2430
rect 82320 2390 82330 2400
rect 82390 2390 82400 2450
rect 83160 2450 83240 2460
rect 83160 2390 83170 2450
rect 83230 2430 83240 2450
rect 83230 2400 83360 2430
rect 83230 2390 83240 2400
rect 82320 2380 82400 2390
rect 82740 2380 82820 2390
rect 83160 2380 83240 2390
rect 82740 2320 82750 2380
rect 82810 2340 82820 2380
rect 82810 2320 83360 2340
rect 82740 2310 83360 2320
rect 83270 1840 83360 1850
rect 83270 1780 83280 1840
rect 83350 1780 83360 1840
rect 83270 1770 83360 1780
rect 83280 1700 83360 1710
rect 83280 1640 83290 1700
rect 83350 1640 83360 1700
rect 83280 1630 83360 1640
rect 82210 1590 82290 1600
rect 82210 1530 82220 1590
rect 82280 1530 82290 1590
rect 82210 1520 82290 1530
rect 82740 1120 83360 1130
rect 82740 1060 82750 1120
rect 82810 1100 83360 1120
rect 82810 1060 82820 1100
rect 82320 1050 82400 1060
rect 82740 1050 82820 1060
rect 83160 1050 83240 1060
rect 82320 1030 82330 1050
rect 82210 1000 82330 1030
rect 82320 990 82330 1000
rect 82390 990 82400 1050
rect 82320 980 82400 990
rect 83160 990 83170 1050
rect 83230 1030 83240 1050
rect 83230 1000 83360 1030
rect 83230 990 83240 1000
rect 83160 980 83240 990
rect 82730 950 82830 970
rect 82730 880 82750 950
rect 82820 880 82830 950
rect 82730 840 82830 880
rect 82730 770 82750 840
rect 82820 770 82830 840
rect 82730 760 82830 770
rect 82320 740 82400 750
rect 82320 720 82330 740
rect 82210 690 82330 720
rect 82320 680 82330 690
rect 82390 680 82400 740
rect 83160 740 83240 750
rect 83160 680 83170 740
rect 83230 720 83240 740
rect 83230 690 83360 720
rect 83230 680 83240 690
rect 82320 670 82400 680
rect 82740 670 82820 680
rect 83160 670 83240 680
rect 82740 610 82750 670
rect 82810 630 82820 670
rect 82810 610 83360 630
rect 82740 600 83360 610
rect 82210 140 82290 150
rect 83540 140 83570 29070
rect 83660 140 83690 29070
rect 83780 140 83810 29070
rect 83900 140 83930 29070
rect 84020 140 84050 29070
rect 84140 140 84170 29070
rect 84260 140 84290 29070
rect 82210 80 82220 140
rect 82280 80 82290 140
rect 82210 70 82290 80
rect 83270 130 83360 140
rect 83270 70 83280 130
rect 83350 70 83360 130
rect 83270 60 83360 70
rect 83280 -10 83360 0
rect 83280 -70 83290 -10
rect 83350 -70 83360 -10
rect 83280 -80 83360 -70
rect 82210 -120 82290 -110
rect 82210 -180 82220 -120
rect 82280 -180 82290 -120
rect 82210 -190 82290 -180
rect 82740 -590 83360 -580
rect 82740 -650 82750 -590
rect 82810 -610 83360 -590
rect 82810 -650 82820 -610
rect 82320 -660 82400 -650
rect 82740 -660 82820 -650
rect 83160 -660 83240 -650
rect 82320 -680 82330 -660
rect 82210 -710 82330 -680
rect 82320 -720 82330 -710
rect 82390 -720 82400 -660
rect 82320 -730 82400 -720
rect 83160 -720 83170 -660
rect 83230 -680 83240 -660
rect 83230 -710 83360 -680
rect 83230 -720 83240 -710
rect 83160 -730 83240 -720
rect 82730 -760 82830 -740
rect 82730 -830 82750 -760
rect 82820 -830 82830 -760
rect 82730 -870 82830 -830
rect 82730 -940 82750 -870
rect 82820 -940 82830 -870
rect 82730 -950 82830 -940
rect 82320 -970 82400 -960
rect 82320 -990 82330 -970
rect 82210 -1020 82330 -990
rect 82320 -1030 82330 -1020
rect 82390 -1030 82400 -970
rect 83160 -970 83240 -960
rect 83160 -1030 83170 -970
rect 83230 -990 83240 -970
rect 83230 -1020 83360 -990
rect 83230 -1030 83240 -1020
rect 82320 -1040 82400 -1030
rect 82740 -1040 82820 -1030
rect 83160 -1040 83240 -1030
rect 82740 -1100 82750 -1040
rect 82810 -1080 82820 -1040
rect 82810 -1100 83360 -1080
rect 82740 -1110 83360 -1100
rect 83270 -1580 83360 -1570
rect 83270 -1640 83280 -1580
rect 83350 -1640 83360 -1580
rect 83270 -1650 83360 -1640
rect 83540 -1710 83570 -110
rect 83660 -1710 83690 -110
rect 83780 -1710 83810 -110
rect 83900 -1710 83930 -110
rect 84020 -1710 84050 -110
rect 84140 -1710 84170 -110
rect 84260 -1710 84290 -110
<< via2 >>
rect 2360 32600 2420 32660
rect -5510 30060 -5450 30120
rect -5240 29930 -5180 29990
rect -5100 29930 -5040 29990
rect -2070 29930 -2010 29990
rect -5360 29790 -5300 29850
rect 2420 32460 2480 32520
rect 3720 30070 3780 30130
rect 2650 29930 2710 29990
rect 7350 32600 7410 32660
rect 7410 32460 7470 32520
rect 8710 30070 8770 30130
rect 7640 29930 7700 29990
rect 3720 29000 3780 29060
rect 2650 28890 2710 28950
rect 3180 28250 3240 28310
rect 3240 28250 3250 28310
rect 3180 28240 3250 28250
rect 3180 28140 3240 28200
rect 3240 28140 3250 28200
rect 3180 28130 3250 28140
rect 12340 32600 12400 32660
rect 12160 32320 12220 32380
rect 12220 32180 12280 32240
rect 8710 29000 8770 29060
rect 7640 28890 7700 28950
rect 8170 28250 8230 28310
rect 8230 28250 8240 28310
rect 8170 28240 8240 28250
rect 8170 28140 8230 28200
rect 8230 28140 8240 28200
rect 8170 28130 8240 28140
rect 12400 32460 12460 32520
rect 13700 30070 13760 30130
rect 12630 29930 12690 29990
rect 17330 32600 17390 32660
rect 13700 29000 13760 29060
rect 12630 28890 12690 28950
rect 13160 28250 13220 28310
rect 13220 28250 13230 28310
rect 13160 28240 13230 28250
rect 13160 28140 13220 28200
rect 13220 28140 13230 28200
rect 13160 28130 13230 28140
rect 17150 32320 17210 32380
rect 17210 32180 17270 32240
rect 17390 32460 17450 32520
rect 18690 30070 18750 30130
rect 17620 29930 17680 29990
rect 22320 32600 22380 32660
rect 18690 29000 18750 29060
rect 17620 28890 17680 28950
rect 18150 28250 18210 28310
rect 18210 28250 18220 28310
rect 18150 28240 18220 28250
rect 18150 28140 18210 28200
rect 18210 28140 18220 28200
rect 18150 28130 18220 28140
rect 22140 32320 22200 32380
rect 21780 32040 21840 32100
rect 21840 31900 21900 31960
rect 21960 31760 22020 31820
rect 22020 31620 22080 31680
rect 22200 32180 22260 32240
rect 22380 32460 22440 32520
rect 23680 30070 23740 30130
rect 22610 29930 22670 29990
rect 27310 32600 27370 32660
rect 23680 29000 23740 29060
rect 22610 28890 22670 28950
rect 23140 28250 23200 28310
rect 23200 28250 23210 28310
rect 23140 28240 23210 28250
rect 23140 28140 23200 28200
rect 23200 28140 23210 28200
rect 23140 28130 23210 28140
rect 27130 32320 27190 32380
rect 26770 32040 26830 32100
rect 26830 31900 26890 31960
rect 26950 31760 27010 31820
rect 27010 31620 27070 31680
rect 27190 32180 27250 32240
rect 27370 32460 27430 32520
rect 28670 30070 28730 30130
rect 27600 29930 27660 29990
rect 32300 32600 32360 32660
rect 28670 29000 28730 29060
rect 27600 28890 27660 28950
rect 28130 28250 28190 28310
rect 28190 28250 28200 28310
rect 28130 28240 28200 28250
rect 28130 28140 28190 28200
rect 28190 28140 28200 28200
rect 28130 28130 28200 28140
rect 32120 32320 32180 32380
rect 31940 32040 32000 32100
rect 31760 31760 31820 31820
rect 31400 31480 31460 31540
rect 31460 31340 31520 31400
rect 31580 31200 31640 31260
rect 31640 31060 31700 31120
rect 31820 31620 31880 31680
rect 32000 31900 32060 31960
rect 32180 32180 32240 32240
rect 32360 32460 32420 32520
rect 33660 30070 33720 30130
rect 32590 29930 32650 29990
rect 37290 32600 37350 32660
rect 33660 29000 33720 29060
rect 32590 28890 32650 28950
rect 33120 28250 33180 28310
rect 33180 28250 33190 28310
rect 33120 28240 33190 28250
rect 33120 28140 33180 28200
rect 33180 28140 33190 28200
rect 33120 28130 33190 28140
rect 37110 32320 37170 32380
rect 36930 32040 36990 32100
rect 36750 31760 36810 31820
rect 36570 31480 36630 31540
rect 36390 30920 36450 30980
rect 36210 30360 36270 30420
rect 36270 30220 36330 30280
rect 36450 30780 36510 30840
rect 36630 31340 36690 31400
rect 36810 31620 36870 31680
rect 36990 31900 37050 31960
rect 37170 32180 37230 32240
rect 37350 32460 37410 32520
rect 38650 30070 38710 30130
rect 37580 29930 37640 29990
rect 42280 32600 42340 32660
rect 38650 29000 38710 29060
rect 37580 28890 37640 28950
rect 38110 28250 38170 28310
rect 38170 28250 38180 28310
rect 38110 28240 38180 28250
rect 38110 28140 38170 28200
rect 38170 28140 38180 28200
rect 38110 28130 38180 28140
rect 42100 32320 42160 32380
rect 41920 32040 41980 32100
rect 41740 31760 41800 31820
rect 41560 31480 41620 31540
rect 41200 30920 41260 30980
rect 41260 30780 41320 30840
rect 41350 30640 41410 30700
rect 41440 30500 41500 30560
rect 41620 31340 41680 31400
rect 41800 31620 41860 31680
rect 41980 31900 42040 31960
rect 42160 32180 42220 32240
rect 42340 32460 42400 32520
rect 43640 30070 43700 30130
rect 42570 29930 42630 29990
rect 47270 32600 47330 32660
rect 43640 29000 43700 29060
rect 42570 28890 42630 28950
rect 43100 28250 43160 28310
rect 43160 28250 43170 28310
rect 43100 28240 43170 28250
rect 43100 28140 43160 28200
rect 43160 28140 43170 28200
rect 43100 28130 43170 28140
rect 47090 32320 47150 32380
rect 46910 32040 46970 32100
rect 46730 31760 46790 31820
rect 46370 31480 46430 31540
rect 46430 31340 46490 31400
rect 46550 31200 46610 31260
rect 46610 31060 46670 31120
rect 46790 31620 46850 31680
rect 46970 31900 47030 31960
rect 47150 32180 47210 32240
rect 47330 32460 47390 32520
rect 48630 30070 48690 30130
rect 47560 29930 47620 29990
rect 52260 32600 52320 32660
rect 48630 29000 48690 29060
rect 47560 28890 47620 28950
rect 48090 28250 48150 28310
rect 48150 28250 48160 28310
rect 48090 28240 48160 28250
rect 48090 28140 48150 28200
rect 48150 28140 48160 28200
rect 48090 28130 48160 28140
rect 52080 32320 52140 32380
rect 51720 32040 51780 32100
rect 51780 31900 51840 31960
rect 51900 31760 51960 31820
rect 51960 31620 52020 31680
rect 52140 32180 52200 32240
rect 52320 32460 52380 32520
rect 53620 30070 53680 30130
rect 52550 29930 52610 29990
rect 57250 32600 57310 32660
rect 53620 29000 53680 29060
rect 52550 28890 52610 28950
rect 53080 28250 53140 28310
rect 53140 28250 53150 28310
rect 53080 28240 53150 28250
rect 53080 28140 53140 28200
rect 53140 28140 53150 28200
rect 53080 28130 53150 28140
rect 57070 32320 57130 32380
rect 56710 32040 56770 32100
rect 56770 31900 56830 31960
rect 56890 31760 56950 31820
rect 56950 31620 57010 31680
rect 57130 32180 57190 32240
rect 57310 32460 57370 32520
rect 58610 30070 58670 30130
rect 57540 29930 57600 29990
rect 62240 32600 62300 32660
rect 58610 29000 58670 29060
rect 57540 28890 57600 28950
rect 58070 28250 58130 28310
rect 58130 28250 58140 28310
rect 58070 28240 58140 28250
rect 58070 28140 58130 28200
rect 58130 28140 58140 28200
rect 58070 28130 58140 28140
rect 62060 32320 62120 32380
rect 62120 32180 62180 32240
rect 62300 32460 62360 32520
rect 63600 30070 63660 30130
rect 62530 29930 62590 29990
rect 67230 32600 67290 32660
rect 63600 29000 63660 29060
rect 62530 28890 62590 28950
rect 63060 28250 63120 28310
rect 63120 28250 63130 28310
rect 63060 28240 63130 28250
rect 63060 28140 63120 28200
rect 63120 28140 63130 28200
rect 63060 28130 63130 28140
rect 67050 32320 67110 32380
rect 67110 32180 67170 32240
rect 67290 32460 67350 32520
rect 68590 30070 68650 30130
rect 67520 29930 67580 29990
rect 72220 32600 72280 32660
rect 68590 29000 68650 29060
rect 67520 28890 67580 28950
rect 68050 28250 68110 28310
rect 68110 28250 68120 28310
rect 68050 28240 68120 28250
rect 68050 28140 68110 28200
rect 68110 28140 68120 28200
rect 68050 28130 68120 28140
rect 72280 32460 72340 32520
rect 73580 30070 73640 30130
rect 72510 29930 72570 29990
rect 77210 32600 77270 32660
rect 77270 32460 77330 32520
rect 78570 30070 78630 30130
rect 77500 29930 77560 29990
rect 73580 29000 73640 29060
rect 72510 28890 72570 28950
rect 73040 28250 73100 28310
rect 73100 28250 73110 28310
rect 73040 28240 73110 28250
rect 73040 28140 73100 28200
rect 73100 28140 73110 28200
rect 73040 28130 73110 28140
rect 82220 29930 82280 29990
rect 78570 29000 78630 29060
rect 77500 28890 77560 28950
rect 78030 28250 78090 28310
rect 78090 28250 78100 28310
rect 78030 28240 78100 28250
rect 78030 28140 78090 28200
rect 78090 28140 78100 28200
rect 78030 28130 78100 28140
rect -1000 23870 -940 23930
rect -2070 23760 -2010 23820
rect -1540 23120 -1480 23180
rect -1480 23120 -1470 23180
rect -1540 23110 -1470 23120
rect -1540 23010 -1480 23070
rect -1480 23010 -1470 23070
rect -1540 23000 -1470 23010
rect -1010 22300 -940 22360
rect -1000 22160 -940 22220
rect -2070 22050 -2010 22110
rect -1540 21410 -1480 21470
rect -1480 21410 -1470 21470
rect -1540 21400 -1470 21410
rect -1540 21300 -1480 21360
rect -1480 21300 -1470 21360
rect -1540 21290 -1470 21300
rect -1010 20590 -940 20650
rect -1000 20450 -940 20510
rect -2070 20340 -2010 20400
rect -1540 19700 -1480 19760
rect -1480 19700 -1470 19760
rect -1540 19690 -1470 19700
rect -1540 19590 -1480 19650
rect -1480 19590 -1470 19650
rect -1540 19580 -1470 19590
rect -1010 18880 -940 18940
rect -1000 18740 -940 18800
rect -2070 18630 -2010 18690
rect -1540 17990 -1480 18050
rect -1480 17990 -1470 18050
rect -1540 17980 -1470 17990
rect -1540 17880 -1480 17940
rect -1480 17880 -1470 17940
rect -1540 17870 -1470 17880
rect -1010 17170 -940 17230
rect -1000 17030 -940 17090
rect -2070 16920 -2010 16980
rect -1540 16280 -1480 16340
rect -1480 16280 -1470 16340
rect -1540 16270 -1470 16280
rect -1540 16170 -1480 16230
rect -1480 16170 -1470 16230
rect -1540 16160 -1470 16170
rect -1010 15460 -940 15520
rect -1000 15320 -940 15380
rect -2070 15210 -2010 15270
rect -1540 14570 -1480 14630
rect -1480 14570 -1470 14630
rect -1540 14560 -1470 14570
rect -1540 14460 -1480 14520
rect -1480 14460 -1470 14520
rect -1540 14450 -1470 14460
rect -1010 13750 -940 13810
rect -1000 13610 -940 13670
rect -2070 13500 -2010 13560
rect -1540 12860 -1480 12920
rect -1480 12860 -1470 12920
rect -1540 12850 -1470 12860
rect -1540 12750 -1480 12810
rect -1480 12750 -1470 12810
rect -1540 12740 -1470 12750
rect -1010 12040 -940 12100
rect -1000 11900 -940 11960
rect -2070 11790 -2010 11850
rect -1540 11150 -1480 11210
rect -1480 11150 -1470 11210
rect -1540 11140 -1470 11150
rect -1540 11040 -1480 11100
rect -1480 11040 -1470 11100
rect -1540 11030 -1470 11040
rect -1010 10330 -940 10390
rect -1000 10190 -940 10250
rect -2070 10080 -2010 10140
rect -1540 9440 -1480 9500
rect -1480 9440 -1470 9500
rect -1540 9430 -1470 9440
rect -1540 9330 -1480 9390
rect -1480 9330 -1470 9390
rect -1540 9320 -1470 9330
rect -1010 8620 -940 8680
rect -1000 8480 -940 8540
rect -2070 8370 -2010 8430
rect -1540 7730 -1480 7790
rect -1480 7730 -1470 7790
rect -1540 7720 -1470 7730
rect -1540 7620 -1480 7680
rect -1480 7620 -1470 7680
rect -1540 7610 -1470 7620
rect -1010 6910 -940 6970
rect -1000 6770 -940 6830
rect -2070 6660 -2010 6720
rect -1540 6020 -1480 6080
rect -1480 6020 -1470 6080
rect -1540 6010 -1470 6020
rect -1540 5910 -1480 5970
rect -1480 5910 -1470 5970
rect -1540 5900 -1470 5910
rect -1010 5200 -940 5260
rect -1000 5060 -940 5120
rect -2070 4950 -2010 5010
rect -1540 4310 -1480 4370
rect -1480 4310 -1470 4370
rect -1540 4300 -1470 4310
rect -1540 4200 -1480 4260
rect -1480 4200 -1470 4260
rect -1540 4190 -1470 4200
rect -1010 3490 -940 3550
rect -1000 3350 -940 3410
rect -2070 3240 -2010 3300
rect -1540 2600 -1480 2660
rect -1480 2600 -1470 2660
rect -1540 2590 -1470 2600
rect -1540 2490 -1480 2550
rect -1480 2490 -1470 2550
rect -1540 2480 -1470 2490
rect -1010 1780 -940 1840
rect -1000 1640 -940 1700
rect -2070 1530 -2010 1590
rect -1540 890 -1480 950
rect -1480 890 -1470 950
rect -1540 880 -1470 890
rect -1540 780 -1480 840
rect -1480 780 -1470 840
rect -1540 770 -1470 780
rect -2070 80 -2010 140
rect -1010 70 -940 130
rect -1000 -70 -940 -10
rect -2070 -180 -2010 -120
rect -1540 -820 -1480 -760
rect -1480 -820 -1470 -760
rect -1540 -830 -1470 -820
rect -1540 -930 -1480 -870
rect -1480 -930 -1470 -870
rect -1540 -940 -1470 -930
rect -1010 -1640 -940 -1580
rect 2650 80 2710 140
rect 3720 -70 3780 -10
rect 3860 -20 3920 40
rect 2650 -180 2710 -120
rect 3180 -820 3240 -760
rect 3240 -820 3250 -760
rect 3180 -830 3250 -820
rect 3180 -930 3240 -870
rect 3240 -930 3250 -870
rect 3180 -940 3250 -930
rect 3720 -1700 3780 -1640
rect 7640 80 7700 140
rect 8710 -70 8770 -10
rect 8850 -20 8910 40
rect 7640 -180 7700 -120
rect 8170 -820 8230 -760
rect 8230 -820 8240 -760
rect 8170 -830 8240 -820
rect 8170 -930 8230 -870
rect 8230 -930 8240 -870
rect 8170 -940 8240 -930
rect 8710 -1700 8770 -1640
rect 12630 80 12690 140
rect 13700 -70 13760 -10
rect 13840 -20 13900 40
rect 12630 -180 12690 -120
rect 13160 -820 13220 -760
rect 13220 -820 13230 -760
rect 13160 -830 13230 -820
rect 13160 -930 13220 -870
rect 13220 -930 13230 -870
rect 13160 -940 13230 -930
rect 13700 -1700 13760 -1640
rect 17620 80 17680 140
rect 18690 -70 18750 -10
rect 18830 -20 18890 40
rect 17620 -180 17680 -120
rect 18150 -820 18210 -760
rect 18210 -820 18220 -760
rect 18150 -830 18220 -820
rect 18150 -930 18210 -870
rect 18210 -930 18220 -870
rect 18150 -940 18220 -930
rect 18690 -1700 18750 -1640
rect 22610 80 22670 140
rect 23680 -70 23740 -10
rect 23820 -20 23880 40
rect 22610 -180 22670 -120
rect 23140 -820 23200 -760
rect 23200 -820 23210 -760
rect 23140 -830 23210 -820
rect 23140 -930 23200 -870
rect 23200 -930 23210 -870
rect 23140 -940 23210 -930
rect 23680 -1700 23740 -1640
rect 27600 80 27660 140
rect 28670 -70 28730 -10
rect 28810 -20 28870 40
rect 27600 -180 27660 -120
rect 28130 -820 28190 -760
rect 28190 -820 28200 -760
rect 28130 -830 28200 -820
rect 28130 -930 28190 -870
rect 28190 -930 28200 -870
rect 28130 -940 28200 -930
rect 28670 -1700 28730 -1640
rect 32590 80 32650 140
rect 33660 -70 33720 -10
rect 33800 -20 33860 40
rect 32590 -180 32650 -120
rect 33120 -820 33180 -760
rect 33180 -820 33190 -760
rect 33120 -830 33190 -820
rect 33120 -930 33180 -870
rect 33180 -930 33190 -870
rect 33120 -940 33190 -930
rect 33660 -1700 33720 -1640
rect 37580 80 37640 140
rect 38650 -70 38710 -10
rect 38790 -20 38850 40
rect 37580 -180 37640 -120
rect 38110 -820 38170 -760
rect 38170 -820 38180 -760
rect 38110 -830 38180 -820
rect 38110 -930 38170 -870
rect 38170 -930 38180 -870
rect 38110 -940 38180 -930
rect 38650 -1700 38710 -1640
rect 42570 80 42630 140
rect 43640 -70 43700 -10
rect 43780 -20 43840 40
rect 42570 -180 42630 -120
rect 43100 -820 43160 -760
rect 43160 -820 43170 -760
rect 43100 -830 43170 -820
rect 43100 -930 43160 -870
rect 43160 -930 43170 -870
rect 43100 -940 43170 -930
rect 43640 -1700 43700 -1640
rect 47560 80 47620 140
rect 48630 -70 48690 -10
rect 48770 -20 48830 40
rect 47560 -180 47620 -120
rect 48090 -820 48150 -760
rect 48150 -820 48160 -760
rect 48090 -830 48160 -820
rect 48090 -930 48150 -870
rect 48150 -930 48160 -870
rect 48090 -940 48160 -930
rect 48630 -1700 48690 -1640
rect 52550 80 52610 140
rect 53620 -70 53680 -10
rect 53760 -20 53820 40
rect 52550 -180 52610 -120
rect 53080 -820 53140 -760
rect 53140 -820 53150 -760
rect 53080 -830 53150 -820
rect 53080 -930 53140 -870
rect 53140 -930 53150 -870
rect 53080 -940 53150 -930
rect 53620 -1700 53680 -1640
rect 57540 80 57600 140
rect 58610 -70 58670 -10
rect 58750 -20 58810 40
rect 57540 -180 57600 -120
rect 58070 -820 58130 -760
rect 58130 -820 58140 -760
rect 58070 -830 58140 -820
rect 58070 -930 58130 -870
rect 58130 -930 58140 -870
rect 58070 -940 58140 -930
rect 58610 -1700 58670 -1640
rect 62530 80 62590 140
rect 63600 -70 63660 -10
rect 63740 -20 63800 40
rect 62530 -180 62590 -120
rect 63060 -820 63120 -760
rect 63120 -820 63130 -760
rect 63060 -830 63130 -820
rect 63060 -930 63120 -870
rect 63120 -930 63130 -870
rect 63060 -940 63130 -930
rect 63600 -1700 63660 -1640
rect 67520 80 67580 140
rect 68590 -70 68650 -10
rect 68730 -20 68790 40
rect 67520 -180 67580 -120
rect 68050 -820 68110 -760
rect 68110 -820 68120 -760
rect 68050 -830 68120 -820
rect 68050 -930 68110 -870
rect 68110 -930 68120 -870
rect 68050 -940 68120 -930
rect 68590 -1700 68650 -1640
rect 72510 80 72570 140
rect 73580 -70 73640 -10
rect 73720 -20 73780 40
rect 72510 -180 72570 -120
rect 73040 -820 73100 -760
rect 73100 -820 73110 -760
rect 73040 -830 73110 -820
rect 73040 -930 73100 -870
rect 73100 -930 73110 -870
rect 73040 -940 73110 -930
rect 73580 -1700 73640 -1640
rect 77500 80 77560 140
rect 78570 -70 78630 -10
rect 77500 -180 77560 -120
rect 78030 -820 78090 -760
rect 78090 -820 78100 -760
rect 78030 -830 78100 -820
rect 78030 -930 78090 -870
rect 78090 -930 78100 -870
rect 78030 -940 78100 -930
rect 78570 -1700 78630 -1640
rect 83290 29000 83350 29060
rect 82220 28890 82280 28950
rect 82750 28250 82810 28310
rect 82810 28250 82820 28310
rect 82750 28240 82820 28250
rect 82750 28140 82810 28200
rect 82810 28140 82820 28200
rect 82750 28130 82820 28140
rect 83280 27430 83350 27490
rect 83290 27290 83350 27350
rect 82220 27180 82280 27240
rect 82750 26540 82810 26600
rect 82810 26540 82820 26600
rect 82750 26530 82820 26540
rect 82750 26430 82810 26490
rect 82810 26430 82820 26490
rect 82750 26420 82820 26430
rect 83280 25720 83350 25780
rect 83290 25580 83350 25640
rect 82220 25470 82280 25530
rect 82750 24830 82810 24890
rect 82810 24830 82820 24890
rect 82750 24820 82820 24830
rect 82750 24720 82810 24780
rect 82810 24720 82820 24780
rect 82750 24710 82820 24720
rect 83280 24010 83350 24070
rect 83290 23870 83350 23930
rect 82220 23760 82280 23820
rect 82750 23120 82810 23180
rect 82810 23120 82820 23180
rect 82750 23110 82820 23120
rect 82750 23010 82810 23070
rect 82810 23010 82820 23070
rect 82750 23000 82820 23010
rect 83280 22300 83350 22360
rect 83290 22160 83350 22220
rect 82220 22050 82280 22110
rect 82750 21410 82810 21470
rect 82810 21410 82820 21470
rect 82750 21400 82820 21410
rect 82750 21300 82810 21360
rect 82810 21300 82820 21360
rect 82750 21290 82820 21300
rect 83280 20590 83350 20650
rect 83290 20450 83350 20510
rect 82220 20340 82280 20400
rect 82750 19700 82810 19760
rect 82810 19700 82820 19760
rect 82750 19690 82820 19700
rect 82750 19590 82810 19650
rect 82810 19590 82820 19650
rect 82750 19580 82820 19590
rect 83280 18880 83350 18940
rect 83290 18740 83350 18800
rect 82220 18630 82280 18690
rect 82750 17990 82810 18050
rect 82810 17990 82820 18050
rect 82750 17980 82820 17990
rect 82750 17880 82810 17940
rect 82810 17880 82820 17940
rect 82750 17870 82820 17880
rect 83280 17170 83350 17230
rect 83290 17030 83350 17090
rect 82220 16920 82280 16980
rect 82750 16280 82810 16340
rect 82810 16280 82820 16340
rect 82750 16270 82820 16280
rect 82750 16170 82810 16230
rect 82810 16170 82820 16230
rect 82750 16160 82820 16170
rect 83280 15460 83350 15520
rect 83290 15320 83350 15380
rect 82220 15210 82280 15270
rect 82750 14570 82810 14630
rect 82810 14570 82820 14630
rect 82750 14560 82820 14570
rect 82750 14460 82810 14520
rect 82810 14460 82820 14520
rect 82750 14450 82820 14460
rect 83280 13750 83350 13810
rect 83290 13610 83350 13670
rect 82220 13500 82280 13560
rect 82750 12860 82810 12920
rect 82810 12860 82820 12920
rect 82750 12850 82820 12860
rect 82750 12750 82810 12810
rect 82810 12750 82820 12810
rect 82750 12740 82820 12750
rect 83280 12040 83350 12100
rect 83290 11900 83350 11960
rect 82220 11790 82280 11850
rect 82750 11150 82810 11210
rect 82810 11150 82820 11210
rect 82750 11140 82820 11150
rect 82750 11040 82810 11100
rect 82810 11040 82820 11100
rect 82750 11030 82820 11040
rect 83280 10330 83350 10390
rect 83290 10190 83350 10250
rect 82220 10080 82280 10140
rect 82750 9440 82810 9500
rect 82810 9440 82820 9500
rect 82750 9430 82820 9440
rect 82750 9330 82810 9390
rect 82810 9330 82820 9390
rect 82750 9320 82820 9330
rect 83280 8620 83350 8680
rect 83290 8480 83350 8540
rect 82220 8370 82280 8430
rect 82750 7730 82810 7790
rect 82810 7730 82820 7790
rect 82750 7720 82820 7730
rect 82750 7620 82810 7680
rect 82810 7620 82820 7680
rect 82750 7610 82820 7620
rect 83280 6910 83350 6970
rect 83290 6770 83350 6830
rect 82220 6660 82280 6720
rect 82750 6020 82810 6080
rect 82810 6020 82820 6080
rect 82750 6010 82820 6020
rect 82750 5910 82810 5970
rect 82810 5910 82820 5970
rect 82750 5900 82820 5910
rect 83280 5200 83350 5260
rect 83290 5060 83350 5120
rect 82220 4950 82280 5010
rect 82750 4310 82810 4370
rect 82810 4310 82820 4370
rect 82750 4300 82820 4310
rect 82750 4200 82810 4260
rect 82810 4200 82820 4260
rect 82750 4190 82820 4200
rect 83280 3490 83350 3550
rect 83290 3350 83350 3410
rect 82220 3240 82280 3300
rect 82750 2600 82810 2660
rect 82810 2600 82820 2660
rect 82750 2590 82820 2600
rect 82750 2490 82810 2550
rect 82810 2490 82820 2550
rect 82750 2480 82820 2490
rect 83280 1780 83350 1840
rect 83290 1640 83350 1700
rect 82220 1530 82280 1590
rect 82750 890 82810 950
rect 82810 890 82820 950
rect 82750 880 82820 890
rect 82750 780 82810 840
rect 82810 780 82820 840
rect 82750 770 82820 780
rect 82220 80 82280 140
rect 83280 70 83350 130
rect 83290 -70 83350 -10
rect 82220 -180 82280 -120
rect 82750 -820 82810 -760
rect 82810 -820 82820 -760
rect 82750 -830 82820 -820
rect 82750 -930 82810 -870
rect 82810 -930 82820 -870
rect 82750 -940 82820 -930
rect 83280 -1640 83350 -1580
<< metal3 >>
rect 2350 32660 2430 32670
rect 2350 32650 2360 32660
rect -5140 32600 2360 32650
rect 2420 32650 2430 32660
rect 7340 32660 7420 32670
rect 7340 32650 7350 32660
rect 2420 32600 7350 32650
rect 7410 32650 7420 32660
rect 12330 32660 12410 32670
rect 12330 32650 12340 32660
rect 7410 32600 12340 32650
rect 12400 32650 12410 32660
rect 17320 32660 17400 32670
rect 17320 32650 17330 32660
rect 12400 32600 17330 32650
rect 17390 32650 17400 32660
rect 22310 32660 22390 32670
rect 22310 32650 22320 32660
rect 17390 32600 22320 32650
rect 22380 32650 22390 32660
rect 27300 32660 27380 32670
rect 27300 32650 27310 32660
rect 22380 32600 27310 32650
rect 27370 32650 27380 32660
rect 32290 32660 32370 32670
rect 32290 32650 32300 32660
rect 27370 32600 32300 32650
rect 32360 32650 32370 32660
rect 37280 32660 37360 32670
rect 37280 32650 37290 32660
rect 32360 32600 37290 32650
rect 37350 32650 37360 32660
rect 42270 32660 42350 32670
rect 42270 32650 42280 32660
rect 37350 32600 42280 32650
rect 42340 32650 42350 32660
rect 47260 32660 47340 32670
rect 47260 32650 47270 32660
rect 42340 32600 47270 32650
rect 47330 32650 47340 32660
rect 52250 32660 52330 32670
rect 52250 32650 52260 32660
rect 47330 32600 52260 32650
rect 52320 32650 52330 32660
rect 57240 32660 57320 32670
rect 57240 32650 57250 32660
rect 52320 32600 57250 32650
rect 57310 32650 57320 32660
rect 62230 32660 62310 32670
rect 62230 32650 62240 32660
rect 57310 32600 62240 32650
rect 62300 32650 62310 32660
rect 67220 32660 67300 32670
rect 67220 32650 67230 32660
rect 62300 32600 67230 32650
rect 67290 32650 67300 32660
rect 72210 32660 72290 32670
rect 72210 32650 72220 32660
rect 67290 32600 72220 32650
rect 72280 32650 72290 32660
rect 77200 32660 77280 32670
rect 77200 32650 77210 32660
rect 72280 32600 77210 32650
rect 77270 32650 77280 32660
rect 77270 32600 84650 32650
rect -5140 32590 84650 32600
rect 2410 32520 2490 32530
rect 2410 32510 2420 32520
rect -5140 32460 2420 32510
rect 2480 32510 2490 32520
rect 7400 32520 7480 32530
rect 7400 32510 7410 32520
rect 2480 32460 7410 32510
rect 7470 32510 7480 32520
rect 12390 32520 12470 32530
rect 12390 32510 12400 32520
rect 7470 32460 12400 32510
rect 12460 32510 12470 32520
rect 17380 32520 17460 32530
rect 17380 32510 17390 32520
rect 12460 32460 17390 32510
rect 17450 32510 17460 32520
rect 22370 32520 22450 32530
rect 22370 32510 22380 32520
rect 17450 32460 22380 32510
rect 22440 32510 22450 32520
rect 27360 32520 27440 32530
rect 27360 32510 27370 32520
rect 22440 32460 27370 32510
rect 27430 32510 27440 32520
rect 32350 32520 32430 32530
rect 32350 32510 32360 32520
rect 27430 32460 32360 32510
rect 32420 32510 32430 32520
rect 37340 32520 37420 32530
rect 37340 32510 37350 32520
rect 32420 32460 37350 32510
rect 37410 32510 37420 32520
rect 42330 32520 42410 32530
rect 42330 32510 42340 32520
rect 37410 32460 42340 32510
rect 42400 32510 42410 32520
rect 47320 32520 47400 32530
rect 47320 32510 47330 32520
rect 42400 32460 47330 32510
rect 47390 32510 47400 32520
rect 52310 32520 52390 32530
rect 52310 32510 52320 32520
rect 47390 32460 52320 32510
rect 52380 32510 52390 32520
rect 57300 32520 57380 32530
rect 57300 32510 57310 32520
rect 52380 32460 57310 32510
rect 57370 32510 57380 32520
rect 62290 32520 62370 32530
rect 62290 32510 62300 32520
rect 57370 32460 62300 32510
rect 62360 32510 62370 32520
rect 67280 32520 67360 32530
rect 67280 32510 67290 32520
rect 62360 32460 67290 32510
rect 67350 32510 67360 32520
rect 72270 32520 72350 32530
rect 72270 32510 72280 32520
rect 67350 32460 72280 32510
rect 72340 32510 72350 32520
rect 77260 32520 77340 32530
rect 77260 32510 77270 32520
rect 72340 32460 77270 32510
rect 77330 32510 77340 32520
rect 77330 32460 84650 32510
rect -5140 32450 84650 32460
rect 12150 32380 12230 32390
rect 12150 32370 12160 32380
rect -5140 32320 12160 32370
rect 12220 32370 12230 32380
rect 17140 32380 17220 32390
rect 17140 32370 17150 32380
rect 12220 32320 17150 32370
rect 17210 32370 17220 32380
rect 22130 32380 22210 32390
rect 22130 32370 22140 32380
rect 17210 32320 22140 32370
rect 22200 32370 22210 32380
rect 27120 32380 27200 32390
rect 27120 32370 27130 32380
rect 22200 32320 27130 32370
rect 27190 32370 27200 32380
rect 32110 32380 32190 32390
rect 32110 32370 32120 32380
rect 27190 32320 32120 32370
rect 32180 32370 32190 32380
rect 37100 32380 37180 32390
rect 37100 32370 37110 32380
rect 32180 32320 37110 32370
rect 37170 32370 37180 32380
rect 42090 32380 42170 32390
rect 42090 32370 42100 32380
rect 37170 32320 42100 32370
rect 42160 32370 42170 32380
rect 47080 32380 47160 32390
rect 47080 32370 47090 32380
rect 42160 32320 47090 32370
rect 47150 32370 47160 32380
rect 52070 32380 52150 32390
rect 52070 32370 52080 32380
rect 47150 32320 52080 32370
rect 52140 32370 52150 32380
rect 57060 32380 57140 32390
rect 57060 32370 57070 32380
rect 52140 32320 57070 32370
rect 57130 32370 57140 32380
rect 62050 32380 62130 32390
rect 62050 32370 62060 32380
rect 57130 32320 62060 32370
rect 62120 32370 62130 32380
rect 67040 32380 67120 32390
rect 67040 32370 67050 32380
rect 62120 32320 67050 32370
rect 67110 32370 67120 32380
rect 67110 32320 84650 32370
rect -5140 32310 84650 32320
rect 12210 32240 12290 32250
rect 12210 32230 12220 32240
rect -5140 32180 12220 32230
rect 12280 32230 12290 32240
rect 17200 32240 17280 32250
rect 17200 32230 17210 32240
rect 12280 32180 17210 32230
rect 17270 32230 17280 32240
rect 22190 32240 22270 32250
rect 22190 32230 22200 32240
rect 17270 32180 22200 32230
rect 22260 32230 22270 32240
rect 27180 32240 27260 32250
rect 27180 32230 27190 32240
rect 22260 32180 27190 32230
rect 27250 32230 27260 32240
rect 32170 32240 32250 32250
rect 32170 32230 32180 32240
rect 27250 32180 32180 32230
rect 32240 32230 32250 32240
rect 37160 32240 37240 32250
rect 37160 32230 37170 32240
rect 32240 32180 37170 32230
rect 37230 32230 37240 32240
rect 42150 32240 42230 32250
rect 42150 32230 42160 32240
rect 37230 32180 42160 32230
rect 42220 32230 42230 32240
rect 47140 32240 47220 32250
rect 47140 32230 47150 32240
rect 42220 32180 47150 32230
rect 47210 32230 47220 32240
rect 52130 32240 52210 32250
rect 52130 32230 52140 32240
rect 47210 32180 52140 32230
rect 52200 32230 52210 32240
rect 57120 32240 57200 32250
rect 57120 32230 57130 32240
rect 52200 32180 57130 32230
rect 57190 32230 57200 32240
rect 62110 32240 62190 32250
rect 62110 32230 62120 32240
rect 57190 32180 62120 32230
rect 62180 32230 62190 32240
rect 67100 32240 67180 32250
rect 67100 32230 67110 32240
rect 62180 32180 67110 32230
rect 67170 32230 67180 32240
rect 67170 32180 84650 32230
rect -5140 32170 84650 32180
rect 21770 32100 21850 32110
rect 21770 32090 21780 32100
rect -5140 32040 21780 32090
rect 21840 32090 21850 32100
rect 26760 32100 26840 32110
rect 26760 32090 26770 32100
rect 21840 32040 26770 32090
rect 26830 32090 26840 32100
rect 31930 32100 32010 32110
rect 31930 32090 31940 32100
rect 26830 32040 31940 32090
rect 32000 32090 32010 32100
rect 36920 32100 37000 32110
rect 36920 32090 36930 32100
rect 32000 32040 36930 32090
rect 36990 32090 37000 32100
rect 41910 32100 41990 32110
rect 41910 32090 41920 32100
rect 36990 32040 41920 32090
rect 41980 32090 41990 32100
rect 46900 32100 46980 32110
rect 46900 32090 46910 32100
rect 41980 32040 46910 32090
rect 46970 32090 46980 32100
rect 51710 32100 51790 32110
rect 51710 32090 51720 32100
rect 46970 32040 51720 32090
rect 51780 32090 51790 32100
rect 56700 32100 56780 32110
rect 56700 32090 56710 32100
rect 51780 32040 56710 32090
rect 56770 32090 56780 32100
rect 56770 32040 84650 32090
rect -5140 32030 84650 32040
rect 21830 31960 21910 31970
rect 21830 31950 21840 31960
rect -5140 31900 21840 31950
rect 21900 31950 21910 31960
rect 26820 31960 26900 31970
rect 26820 31950 26830 31960
rect 21900 31900 26830 31950
rect 26890 31950 26900 31960
rect 31990 31960 32070 31970
rect 31990 31950 32000 31960
rect 26890 31900 32000 31950
rect 32060 31950 32070 31960
rect 36980 31960 37060 31970
rect 36980 31950 36990 31960
rect 32060 31900 36990 31950
rect 37050 31950 37060 31960
rect 41970 31960 42050 31970
rect 41970 31950 41980 31960
rect 37050 31900 41980 31950
rect 42040 31950 42050 31960
rect 46960 31960 47040 31970
rect 46960 31950 46970 31960
rect 42040 31900 46970 31950
rect 47030 31950 47040 31960
rect 51770 31960 51850 31970
rect 51770 31950 51780 31960
rect 47030 31900 51780 31950
rect 51840 31950 51850 31960
rect 56760 31960 56840 31970
rect 56760 31950 56770 31960
rect 51840 31900 56770 31950
rect 56830 31950 56840 31960
rect 56830 31900 84650 31950
rect -5140 31890 84650 31900
rect 21950 31820 22030 31830
rect 21950 31810 21960 31820
rect -5140 31760 21960 31810
rect 22020 31810 22030 31820
rect 26940 31820 27020 31830
rect 26940 31810 26950 31820
rect 22020 31760 26950 31810
rect 27010 31810 27020 31820
rect 31750 31820 31830 31830
rect 31750 31810 31760 31820
rect 27010 31760 31760 31810
rect 31820 31810 31830 31820
rect 36740 31820 36820 31830
rect 36740 31810 36750 31820
rect 31820 31760 36750 31810
rect 36810 31810 36820 31820
rect 41730 31820 41810 31830
rect 41730 31810 41740 31820
rect 36810 31760 41740 31810
rect 41800 31810 41810 31820
rect 46720 31820 46800 31830
rect 46720 31810 46730 31820
rect 41800 31760 46730 31810
rect 46790 31810 46800 31820
rect 51890 31820 51970 31830
rect 51890 31810 51900 31820
rect 46790 31760 51900 31810
rect 51960 31810 51970 31820
rect 56880 31820 56960 31830
rect 56880 31810 56890 31820
rect 51960 31760 56890 31810
rect 56950 31810 56960 31820
rect 56950 31760 84650 31810
rect -5140 31750 84650 31760
rect 22010 31680 22090 31690
rect 22010 31670 22020 31680
rect -5140 31620 22020 31670
rect 22080 31670 22090 31680
rect 27000 31680 27080 31690
rect 27000 31670 27010 31680
rect 22080 31620 27010 31670
rect 27070 31670 27080 31680
rect 31810 31680 31890 31690
rect 31810 31670 31820 31680
rect 27070 31620 31820 31670
rect 31880 31670 31890 31680
rect 36800 31680 36880 31690
rect 36800 31670 36810 31680
rect 31880 31620 36810 31670
rect 36870 31670 36880 31680
rect 41790 31680 41870 31690
rect 41790 31670 41800 31680
rect 36870 31620 41800 31670
rect 41860 31670 41870 31680
rect 46780 31680 46860 31690
rect 46780 31670 46790 31680
rect 41860 31620 46790 31670
rect 46850 31670 46860 31680
rect 51950 31680 52030 31690
rect 51950 31670 51960 31680
rect 46850 31620 51960 31670
rect 52020 31670 52030 31680
rect 56940 31680 57020 31690
rect 56940 31670 56950 31680
rect 52020 31620 56950 31670
rect 57010 31670 57020 31680
rect 57010 31620 84650 31670
rect -5140 31610 84650 31620
rect 31390 31540 31470 31550
rect 31390 31530 31400 31540
rect -5140 31480 31400 31530
rect 31460 31530 31470 31540
rect 36560 31540 36640 31550
rect 36560 31530 36570 31540
rect 31460 31480 36570 31530
rect 36630 31530 36640 31540
rect 41550 31540 41630 31550
rect 41550 31530 41560 31540
rect 36630 31480 41560 31530
rect 41620 31530 41630 31540
rect 46360 31540 46440 31550
rect 46360 31530 46370 31540
rect 41620 31480 46370 31530
rect 46430 31530 46440 31540
rect 46430 31480 84650 31530
rect -5140 31470 84650 31480
rect 31450 31400 31530 31410
rect 31450 31390 31460 31400
rect -5140 31340 31460 31390
rect 31520 31390 31530 31400
rect 36620 31400 36700 31410
rect 36620 31390 36630 31400
rect 31520 31340 36630 31390
rect 36690 31390 36700 31400
rect 41610 31400 41690 31410
rect 41610 31390 41620 31400
rect 36690 31340 41620 31390
rect 41680 31390 41690 31400
rect 46420 31400 46500 31410
rect 46420 31390 46430 31400
rect 41680 31340 46430 31390
rect 46490 31390 46500 31400
rect 46490 31340 84650 31390
rect -5140 31330 84650 31340
rect 31570 31260 31650 31270
rect 31570 31250 31580 31260
rect -5140 31200 31580 31250
rect 31640 31250 31650 31260
rect 46540 31260 46620 31270
rect 46540 31250 46550 31260
rect 31640 31200 46550 31250
rect 46610 31250 46620 31260
rect 46610 31200 84650 31250
rect -5140 31190 84650 31200
rect 31630 31120 31710 31130
rect 31630 31110 31640 31120
rect -5140 31060 31640 31110
rect 31700 31110 31710 31120
rect 46600 31120 46680 31130
rect 46600 31110 46610 31120
rect 31700 31060 46610 31110
rect 46670 31110 46680 31120
rect 46670 31060 84650 31110
rect -5140 31050 84650 31060
rect 36380 30980 36460 30990
rect 36380 30970 36390 30980
rect -5140 30920 36390 30970
rect 36450 30970 36460 30980
rect 41190 30980 41270 30990
rect 41190 30970 41200 30980
rect 36450 30920 41200 30970
rect 41260 30970 41270 30980
rect 41260 30920 84650 30970
rect -5140 30910 84650 30920
rect 36440 30840 36520 30850
rect 36440 30830 36450 30840
rect -5140 30780 36450 30830
rect 36510 30830 36520 30840
rect 41250 30840 41330 30850
rect 41250 30830 41260 30840
rect 36510 30780 41260 30830
rect 41320 30830 41330 30840
rect 41320 30780 84650 30830
rect -5140 30770 84650 30780
rect 41340 30700 41420 30710
rect 41340 30690 41350 30700
rect -5140 30640 41350 30690
rect 41410 30690 41420 30700
rect 41410 30640 84650 30690
rect -5140 30630 84650 30640
rect 41430 30560 41510 30570
rect 41430 30550 41440 30560
rect -5140 30500 41440 30550
rect 41500 30550 41510 30560
rect 41500 30500 84650 30550
rect -5140 30490 84650 30500
rect 36200 30420 36280 30430
rect 36200 30410 36210 30420
rect -5180 30400 36210 30410
rect -5580 30360 36210 30400
rect 36270 30410 36280 30420
rect 36270 30360 84650 30410
rect -5580 30350 84650 30360
rect -5580 30340 -5140 30350
rect 36260 30280 36340 30290
rect 36260 30270 36270 30280
rect -5180 30260 36270 30270
rect -5580 30220 36270 30260
rect 36330 30270 36340 30280
rect 36330 30220 84650 30270
rect -5580 30210 84650 30220
rect -5580 30200 -5140 30210
rect -5530 30130 -5430 30140
rect -5530 30050 -5520 30130
rect -5440 30050 -5430 30130
rect 3710 30130 3790 30140
rect 3710 30120 3720 30130
rect -5530 30040 -5430 30050
rect -5370 30070 3720 30120
rect 3780 30120 3790 30130
rect 8700 30130 8780 30140
rect 8700 30120 8710 30130
rect 3780 30070 8710 30120
rect 8770 30120 8780 30130
rect 13690 30130 13770 30140
rect 13690 30120 13700 30130
rect 8770 30070 13700 30120
rect 13760 30120 13770 30130
rect 18680 30130 18760 30140
rect 18680 30120 18690 30130
rect 13760 30070 18690 30120
rect 18750 30120 18760 30130
rect 23670 30130 23750 30140
rect 23670 30120 23680 30130
rect 18750 30070 23680 30120
rect 23740 30120 23750 30130
rect 28660 30130 28740 30140
rect 28660 30120 28670 30130
rect 23740 30070 28670 30120
rect 28730 30120 28740 30130
rect 33650 30130 33730 30140
rect 33650 30120 33660 30130
rect 28730 30070 33660 30120
rect 33720 30120 33730 30130
rect 38640 30130 38720 30140
rect 38640 30120 38650 30130
rect 33720 30070 38650 30120
rect 38710 30120 38720 30130
rect 43630 30130 43710 30140
rect 43630 30120 43640 30130
rect 38710 30070 43640 30120
rect 43700 30120 43710 30130
rect 48620 30130 48700 30140
rect 48620 30120 48630 30130
rect 43700 30070 48630 30120
rect 48690 30120 48700 30130
rect 53610 30130 53690 30140
rect 53610 30120 53620 30130
rect 48690 30070 53620 30120
rect 53680 30120 53690 30130
rect 58600 30130 58680 30140
rect 58600 30120 58610 30130
rect 53680 30070 58610 30120
rect 58670 30120 58680 30130
rect 63590 30130 63670 30140
rect 63590 30120 63600 30130
rect 58670 30070 63600 30120
rect 63660 30120 63670 30130
rect 68580 30130 68660 30140
rect 68580 30120 68590 30130
rect 63660 30070 68590 30120
rect 68650 30120 68660 30130
rect 73570 30130 73650 30140
rect 73570 30120 73580 30130
rect 68650 30070 73580 30120
rect 73640 30120 73650 30130
rect 78560 30130 78640 30140
rect 78560 30120 78570 30130
rect 73640 30070 78570 30120
rect 78630 30120 78640 30130
rect 78630 30070 84650 30120
rect -5370 30060 84650 30070
rect -6370 29900 -6300 29990
rect -5370 29860 -5310 30060
rect -5250 29990 -5170 30000
rect -5250 29930 -5240 29990
rect -5180 29980 -5170 29990
rect -5110 29990 -5030 30000
rect -5110 29980 -5100 29990
rect -5180 29930 -5100 29980
rect -5040 29980 -5030 29990
rect -2080 29990 -2000 30000
rect -2080 29980 -2070 29990
rect -5040 29930 -2070 29980
rect -2010 29980 -2000 29990
rect 2640 29990 2720 30000
rect 2640 29980 2650 29990
rect -2010 29930 2650 29980
rect 2710 29980 2720 29990
rect 7630 29990 7710 30000
rect 7630 29980 7640 29990
rect 2710 29930 7640 29980
rect 7700 29980 7710 29990
rect 12620 29990 12700 30000
rect 12620 29980 12630 29990
rect 7700 29930 12630 29980
rect 12690 29980 12700 29990
rect 17610 29990 17690 30000
rect 17610 29980 17620 29990
rect 12690 29930 17620 29980
rect 17680 29980 17690 29990
rect 22600 29990 22680 30000
rect 22600 29980 22610 29990
rect 17680 29930 22610 29980
rect 22670 29980 22680 29990
rect 27590 29990 27670 30000
rect 27590 29980 27600 29990
rect 22670 29930 27600 29980
rect 27660 29980 27670 29990
rect 32580 29990 32660 30000
rect 32580 29980 32590 29990
rect 27660 29930 32590 29980
rect 32650 29980 32660 29990
rect 37570 29990 37650 30000
rect 37570 29980 37580 29990
rect 32650 29930 37580 29980
rect 37640 29980 37650 29990
rect 42560 29990 42640 30000
rect 42560 29980 42570 29990
rect 37640 29930 42570 29980
rect 42630 29980 42640 29990
rect 47550 29990 47630 30000
rect 47550 29980 47560 29990
rect 42630 29930 47560 29980
rect 47620 29980 47630 29990
rect 52540 29990 52620 30000
rect 52540 29980 52550 29990
rect 47620 29930 52550 29980
rect 52610 29980 52620 29990
rect 57530 29990 57610 30000
rect 57530 29980 57540 29990
rect 52610 29930 57540 29980
rect 57600 29980 57610 29990
rect 62520 29990 62600 30000
rect 62520 29980 62530 29990
rect 57600 29930 62530 29980
rect 62590 29980 62600 29990
rect 67510 29990 67590 30000
rect 67510 29980 67520 29990
rect 62590 29930 67520 29980
rect 67580 29980 67590 29990
rect 72500 29990 72580 30000
rect 72500 29980 72510 29990
rect 67580 29930 72510 29980
rect 72570 29980 72580 29990
rect 77490 29990 77570 30000
rect 77490 29980 77500 29990
rect 72570 29930 77500 29980
rect 77560 29980 77570 29990
rect 82210 29990 82290 30000
rect 82210 29980 82220 29990
rect 77560 29930 82220 29980
rect 82280 29980 82290 29990
rect 82280 29930 84650 29980
rect -5250 29920 84650 29930
rect -5370 29850 -5290 29860
rect -5370 29790 -5360 29850
rect -5300 29790 -5290 29850
rect -5370 29780 -5290 29790
rect 3710 29060 3790 29070
rect 3710 29000 3720 29060
rect 3780 29000 3790 29060
rect 3710 28990 3790 29000
rect 8700 29060 8780 29070
rect 8700 29000 8710 29060
rect 8770 29000 8780 29060
rect 8700 28990 8780 29000
rect 13690 29060 13770 29070
rect 13690 29000 13700 29060
rect 13760 29000 13770 29060
rect 13690 28990 13770 29000
rect 18680 29060 18760 29070
rect 18680 29000 18690 29060
rect 18750 29000 18760 29060
rect 18680 28990 18760 29000
rect 23670 29060 23750 29070
rect 23670 29000 23680 29060
rect 23740 29000 23750 29060
rect 23670 28990 23750 29000
rect 28660 29060 28740 29070
rect 28660 29000 28670 29060
rect 28730 29000 28740 29060
rect 28660 28990 28740 29000
rect 33650 29060 33730 29070
rect 33650 29000 33660 29060
rect 33720 29000 33730 29060
rect 33650 28990 33730 29000
rect 38640 29060 38720 29070
rect 38640 29000 38650 29060
rect 38710 29000 38720 29060
rect 38640 28990 38720 29000
rect 43630 29060 43710 29070
rect 43630 29000 43640 29060
rect 43700 29000 43710 29060
rect 43630 28990 43710 29000
rect 48620 29060 48700 29070
rect 48620 29000 48630 29060
rect 48690 29000 48700 29060
rect 48620 28990 48700 29000
rect 53610 29060 53690 29070
rect 53610 29000 53620 29060
rect 53680 29000 53690 29060
rect 53610 28990 53690 29000
rect 58600 29060 58680 29070
rect 58600 29000 58610 29060
rect 58670 29000 58680 29060
rect 58600 28990 58680 29000
rect 63590 29060 63670 29070
rect 63590 29000 63600 29060
rect 63660 29000 63670 29060
rect 63590 28990 63670 29000
rect 68580 29060 68660 29070
rect 68580 29000 68590 29060
rect 68650 29000 68660 29060
rect 68580 28990 68660 29000
rect 73570 29060 73650 29070
rect 73570 29000 73580 29060
rect 73640 29000 73650 29060
rect 73570 28990 73650 29000
rect 78560 29060 78640 29070
rect 78560 29000 78570 29060
rect 78630 29000 78640 29060
rect 78560 28990 78640 29000
rect 83280 29060 83360 29070
rect 83280 29000 83290 29060
rect 83350 29000 83360 29060
rect 83280 28990 83360 29000
rect 0 28950 2720 28960
rect 0 28932 2650 28950
rect 0 27508 1688 28932
rect 1752 28900 2650 28932
rect 1752 27508 1772 28900
rect 2640 28890 2650 28900
rect 2710 28890 2720 28950
rect 2640 28870 2720 28890
rect 3140 28310 3280 28350
rect 3140 28240 3170 28310
rect 3250 28240 3280 28310
rect 3140 28200 3280 28240
rect 3140 28130 3170 28200
rect 3250 28130 3280 28200
rect 3140 28100 3280 28130
rect 3730 27530 3790 28990
rect 4990 28950 7710 28960
rect 4990 28932 7640 28950
rect 0 27480 1772 27508
rect 4990 27508 6678 28932
rect 6742 28900 7640 28932
rect 6742 27508 6762 28900
rect 7630 28890 7640 28900
rect 7700 28890 7710 28950
rect 7630 28870 7710 28890
rect 8130 28310 8270 28350
rect 8130 28240 8160 28310
rect 8240 28240 8270 28310
rect 8130 28200 8270 28240
rect 8130 28130 8160 28200
rect 8240 28130 8270 28200
rect 8130 28100 8270 28130
rect 8720 27530 8780 28990
rect 9980 28950 12700 28960
rect 9980 28932 12630 28950
rect 4990 27480 6762 27508
rect 9980 27508 11668 28932
rect 11732 28900 12630 28932
rect 11732 27508 11752 28900
rect 12620 28890 12630 28900
rect 12690 28890 12700 28950
rect 12620 28870 12700 28890
rect 13120 28310 13260 28350
rect 13120 28240 13150 28310
rect 13230 28240 13260 28310
rect 13120 28200 13260 28240
rect 13120 28130 13150 28200
rect 13230 28130 13260 28200
rect 13120 28100 13260 28130
rect 13710 27530 13770 28990
rect 14970 28950 17690 28960
rect 14970 28932 17620 28950
rect 9980 27480 11752 27508
rect 14970 27508 16658 28932
rect 16722 28900 17620 28932
rect 16722 27508 16742 28900
rect 17610 28890 17620 28900
rect 17680 28890 17690 28950
rect 17610 28870 17690 28890
rect 18110 28310 18250 28350
rect 18110 28240 18140 28310
rect 18220 28240 18250 28310
rect 18110 28200 18250 28240
rect 18110 28130 18140 28200
rect 18220 28130 18250 28200
rect 18110 28100 18250 28130
rect 18700 27530 18760 28990
rect 19960 28950 22680 28960
rect 19960 28932 22610 28950
rect 14970 27480 16742 27508
rect 19960 27508 21648 28932
rect 21712 28900 22610 28932
rect 21712 27508 21732 28900
rect 22600 28890 22610 28900
rect 22670 28890 22680 28950
rect 22600 28870 22680 28890
rect 23100 28310 23240 28350
rect 23100 28240 23130 28310
rect 23210 28240 23240 28310
rect 23100 28200 23240 28240
rect 23100 28130 23130 28200
rect 23210 28130 23240 28200
rect 23100 28100 23240 28130
rect 23690 27530 23750 28990
rect 24950 28950 27670 28960
rect 24950 28932 27600 28950
rect 19960 27480 21732 27508
rect 24950 27508 26638 28932
rect 26702 28900 27600 28932
rect 26702 27508 26722 28900
rect 27590 28890 27600 28900
rect 27660 28890 27670 28950
rect 27590 28870 27670 28890
rect 28090 28310 28230 28350
rect 28090 28240 28120 28310
rect 28200 28240 28230 28310
rect 28090 28200 28230 28240
rect 28090 28130 28120 28200
rect 28200 28130 28230 28200
rect 28090 28100 28230 28130
rect 28680 27530 28740 28990
rect 29940 28950 32660 28960
rect 29940 28932 32590 28950
rect 24950 27480 26722 27508
rect 29940 27508 31628 28932
rect 31692 28900 32590 28932
rect 31692 27508 31712 28900
rect 32580 28890 32590 28900
rect 32650 28890 32660 28950
rect 32580 28870 32660 28890
rect 33080 28310 33220 28350
rect 33080 28240 33110 28310
rect 33190 28240 33220 28310
rect 33080 28200 33220 28240
rect 33080 28130 33110 28200
rect 33190 28130 33220 28200
rect 33080 28100 33220 28130
rect 33670 27530 33730 28990
rect 34930 28950 37650 28960
rect 34930 28932 37580 28950
rect 29940 27480 31712 27508
rect 34930 27508 36618 28932
rect 36682 28900 37580 28932
rect 36682 27508 36702 28900
rect 37570 28890 37580 28900
rect 37640 28890 37650 28950
rect 37570 28870 37650 28890
rect 38070 28310 38210 28350
rect 38070 28240 38100 28310
rect 38180 28240 38210 28310
rect 38070 28200 38210 28240
rect 38070 28130 38100 28200
rect 38180 28130 38210 28200
rect 38070 28100 38210 28130
rect 38660 27530 38720 28990
rect 39920 28950 42640 28960
rect 39920 28932 42570 28950
rect 34930 27480 36702 27508
rect 39920 27508 41608 28932
rect 41672 28900 42570 28932
rect 41672 27508 41692 28900
rect 42560 28890 42570 28900
rect 42630 28890 42640 28950
rect 42560 28870 42640 28890
rect 43060 28310 43200 28350
rect 43060 28240 43090 28310
rect 43170 28240 43200 28310
rect 43060 28200 43200 28240
rect 43060 28130 43090 28200
rect 43170 28130 43200 28200
rect 43060 28100 43200 28130
rect 43650 27530 43710 28990
rect 44910 28950 47630 28960
rect 44910 28932 47560 28950
rect 39920 27480 41692 27508
rect 44910 27508 46598 28932
rect 46662 28900 47560 28932
rect 46662 27508 46682 28900
rect 47550 28890 47560 28900
rect 47620 28890 47630 28950
rect 47550 28870 47630 28890
rect 48050 28310 48190 28350
rect 48050 28240 48080 28310
rect 48160 28240 48190 28310
rect 48050 28200 48190 28240
rect 48050 28130 48080 28200
rect 48160 28130 48190 28200
rect 48050 28100 48190 28130
rect 48640 27530 48700 28990
rect 49900 28950 52620 28960
rect 49900 28932 52550 28950
rect 44910 27480 46682 27508
rect 49900 27508 51588 28932
rect 51652 28900 52550 28932
rect 51652 27508 51672 28900
rect 52540 28890 52550 28900
rect 52610 28890 52620 28950
rect 52540 28870 52620 28890
rect 53040 28310 53180 28350
rect 53040 28240 53070 28310
rect 53150 28240 53180 28310
rect 53040 28200 53180 28240
rect 53040 28130 53070 28200
rect 53150 28130 53180 28200
rect 53040 28100 53180 28130
rect 53630 27530 53690 28990
rect 54890 28950 57610 28960
rect 54890 28932 57540 28950
rect 49900 27480 51672 27508
rect 54890 27508 56578 28932
rect 56642 28900 57540 28932
rect 56642 27508 56662 28900
rect 57530 28890 57540 28900
rect 57600 28890 57610 28950
rect 57530 28870 57610 28890
rect 58030 28310 58170 28350
rect 58030 28240 58060 28310
rect 58140 28240 58170 28310
rect 58030 28200 58170 28240
rect 58030 28130 58060 28200
rect 58140 28130 58170 28200
rect 58030 28100 58170 28130
rect 58620 27530 58680 28990
rect 59880 28950 62600 28960
rect 59880 28932 62530 28950
rect 54890 27480 56662 27508
rect 59880 27508 61568 28932
rect 61632 28900 62530 28932
rect 61632 27508 61652 28900
rect 62520 28890 62530 28900
rect 62590 28890 62600 28950
rect 62520 28870 62600 28890
rect 63020 28310 63160 28350
rect 63020 28240 63050 28310
rect 63130 28240 63160 28310
rect 63020 28200 63160 28240
rect 63020 28130 63050 28200
rect 63130 28130 63160 28200
rect 63020 28100 63160 28130
rect 63610 27530 63670 28990
rect 64870 28950 67590 28960
rect 64870 28932 67520 28950
rect 59880 27480 61652 27508
rect 64870 27508 66558 28932
rect 66622 28900 67520 28932
rect 66622 27508 66642 28900
rect 67510 28890 67520 28900
rect 67580 28890 67590 28950
rect 67510 28870 67590 28890
rect 68010 28310 68150 28350
rect 68010 28240 68040 28310
rect 68120 28240 68150 28310
rect 68010 28200 68150 28240
rect 68010 28130 68040 28200
rect 68120 28130 68150 28200
rect 68010 28100 68150 28130
rect 68600 27530 68660 28990
rect 69860 28950 72580 28960
rect 69860 28932 72510 28950
rect 64870 27480 66642 27508
rect 69860 27508 71548 28932
rect 71612 28900 72510 28932
rect 71612 27508 71632 28900
rect 72500 28890 72510 28900
rect 72570 28890 72580 28950
rect 72500 28870 72580 28890
rect 73000 28310 73140 28350
rect 73000 28240 73030 28310
rect 73110 28240 73140 28310
rect 73000 28200 73140 28240
rect 73000 28130 73030 28200
rect 73110 28130 73140 28200
rect 73000 28100 73140 28130
rect 73590 27530 73650 28990
rect 74850 28950 77570 28960
rect 74850 28932 77500 28950
rect 69860 27480 71632 27508
rect 74850 27508 76538 28932
rect 76602 28900 77500 28932
rect 76602 27508 76622 28900
rect 77490 28890 77500 28900
rect 77560 28890 77570 28950
rect 77490 28870 77570 28890
rect 77990 28310 78130 28350
rect 77990 28240 78020 28310
rect 78100 28240 78130 28310
rect 77990 28200 78130 28240
rect 77990 28130 78020 28200
rect 78100 28130 78130 28200
rect 77990 28100 78130 28130
rect 78580 27530 78640 28990
rect 79570 28950 82290 28960
rect 79570 28932 82220 28950
rect 74850 27480 76622 27508
rect 79570 27508 81258 28932
rect 81322 28900 82220 28932
rect 81322 27508 81342 28900
rect 82210 28890 82220 28900
rect 82280 28890 82290 28950
rect 82210 28870 82290 28890
rect 82710 28310 82850 28350
rect 82710 28240 82740 28310
rect 82820 28240 82850 28310
rect 82710 28200 82850 28240
rect 82710 28130 82740 28200
rect 82820 28130 82850 28200
rect 82710 28100 82850 28130
rect 79570 27480 81342 27508
rect 83300 27500 83360 28990
rect 83270 27490 83360 27500
rect 3730 27460 3790 27470
rect 8720 27460 8780 27470
rect 13710 27460 13770 27470
rect 18700 27460 18760 27470
rect 23690 27460 23750 27470
rect 28680 27460 28740 27470
rect 33670 27460 33730 27470
rect 38660 27460 38720 27470
rect 43650 27460 43710 27470
rect 48640 27460 48700 27470
rect 53630 27460 53690 27470
rect 58620 27460 58680 27470
rect 63610 27460 63670 27470
rect 68600 27460 68660 27470
rect 73590 27460 73650 27470
rect 78580 27460 78640 27470
rect 3780 27420 3790 27460
rect 8770 27420 8780 27460
rect 13760 27420 13770 27460
rect 18750 27420 18760 27460
rect 23740 27420 23750 27460
rect 28730 27420 28740 27460
rect 33720 27420 33730 27460
rect 38710 27420 38720 27460
rect 43700 27420 43710 27460
rect 48690 27420 48700 27460
rect 53680 27420 53690 27460
rect 58670 27420 58680 27460
rect 63660 27420 63670 27460
rect 68650 27420 68660 27460
rect 73640 27420 73650 27460
rect 78630 27420 78640 27460
rect 83270 27430 83280 27490
rect 83350 27430 83360 27490
rect 83270 27420 83360 27430
rect 83280 27350 83360 27360
rect 83280 27290 83290 27350
rect 83350 27290 83360 27350
rect 83280 27280 83360 27290
rect 79570 27240 82290 27250
rect 79570 27222 82220 27240
rect 79570 25798 81258 27222
rect 81322 27190 82220 27222
rect 81322 25798 81342 27190
rect 82210 27180 82220 27190
rect 82280 27180 82290 27240
rect 82210 27160 82290 27180
rect 82710 26600 82850 26640
rect 82710 26530 82740 26600
rect 82820 26530 82850 26600
rect 82710 26490 82850 26530
rect 82710 26420 82740 26490
rect 82820 26420 82850 26490
rect 82710 26390 82850 26420
rect 79570 25770 81342 25798
rect 83300 25790 83360 27280
rect 83270 25780 83360 25790
rect 83270 25720 83280 25780
rect 83350 25720 83360 25780
rect 83270 25710 83360 25720
rect 83280 25640 83360 25650
rect 83280 25580 83290 25640
rect 83350 25580 83360 25640
rect 83280 25570 83360 25580
rect 79570 25530 82290 25540
rect 79570 25512 82220 25530
rect 79570 24088 81258 25512
rect 81322 25480 82220 25512
rect 81322 24088 81342 25480
rect 82210 25470 82220 25480
rect 82280 25470 82290 25530
rect 82210 25450 82290 25470
rect 82710 24890 82850 24930
rect 82710 24820 82740 24890
rect 82820 24820 82850 24890
rect 82710 24780 82850 24820
rect 82710 24710 82740 24780
rect 82820 24710 82850 24780
rect 82710 24680 82850 24710
rect 79570 24060 81342 24088
rect 83300 24080 83360 25570
rect 83270 24070 83360 24080
rect 83270 24010 83280 24070
rect 83350 24010 83360 24070
rect 83270 24000 83360 24010
rect -1010 23930 -930 23940
rect -1010 23870 -1000 23930
rect -940 23870 -930 23930
rect -1010 23860 -930 23870
rect 83280 23930 83360 23940
rect 83280 23870 83290 23930
rect 83350 23870 83360 23930
rect 83280 23860 83360 23870
rect -4720 23820 -2000 23830
rect -4720 23802 -2070 23820
rect -4720 22378 -3032 23802
rect -2968 23770 -2070 23802
rect -2968 22378 -2948 23770
rect -2080 23760 -2070 23770
rect -2010 23760 -2000 23820
rect -2080 23740 -2000 23760
rect -1580 23180 -1440 23220
rect -1580 23110 -1550 23180
rect -1470 23110 -1440 23180
rect -1580 23070 -1440 23110
rect -1580 23000 -1550 23070
rect -1470 23000 -1440 23070
rect -1580 22970 -1440 23000
rect -4720 22350 -2948 22378
rect -990 22370 -930 23860
rect -1020 22360 -930 22370
rect -1020 22300 -1010 22360
rect -940 22300 -930 22360
rect 79570 23820 82290 23830
rect 79570 23802 82220 23820
rect 79570 22378 81258 23802
rect 81322 23770 82220 23802
rect 81322 22378 81342 23770
rect 82210 23760 82220 23770
rect 82280 23760 82290 23820
rect 82210 23740 82290 23760
rect 82710 23180 82850 23220
rect 82710 23110 82740 23180
rect 82820 23110 82850 23180
rect 82710 23070 82850 23110
rect 82710 23000 82740 23070
rect 82820 23000 82850 23070
rect 82710 22970 82850 23000
rect 79570 22350 81342 22378
rect 83300 22370 83360 23860
rect 83270 22360 83360 22370
rect -1020 22290 -930 22300
rect 83270 22300 83280 22360
rect 83350 22300 83360 22360
rect 83270 22290 83360 22300
rect -1010 22220 -930 22230
rect -1010 22160 -1000 22220
rect -940 22160 -930 22220
rect -1010 22150 -930 22160
rect 83280 22220 83360 22230
rect 83280 22160 83290 22220
rect 83350 22160 83360 22220
rect 83280 22150 83360 22160
rect -4720 22110 -2000 22120
rect -4720 22092 -2070 22110
rect -4720 20668 -3032 22092
rect -2968 22060 -2070 22092
rect -2968 20668 -2948 22060
rect -2080 22050 -2070 22060
rect -2010 22050 -2000 22110
rect -2080 22030 -2000 22050
rect -1580 21470 -1440 21510
rect -1580 21400 -1550 21470
rect -1470 21400 -1440 21470
rect -1580 21360 -1440 21400
rect -1580 21290 -1550 21360
rect -1470 21290 -1440 21360
rect -1580 21260 -1440 21290
rect -4720 20640 -2948 20668
rect -990 20660 -930 22150
rect -1020 20650 -930 20660
rect -1020 20590 -1010 20650
rect -940 20590 -930 20650
rect 79570 22110 82290 22120
rect 79570 22092 82220 22110
rect 79570 20668 81258 22092
rect 81322 22060 82220 22092
rect 81322 20668 81342 22060
rect 82210 22050 82220 22060
rect 82280 22050 82290 22110
rect 82210 22030 82290 22050
rect 82710 21470 82850 21510
rect 82710 21400 82740 21470
rect 82820 21400 82850 21470
rect 82710 21360 82850 21400
rect 82710 21290 82740 21360
rect 82820 21290 82850 21360
rect 82710 21260 82850 21290
rect 79570 20640 81342 20668
rect 83300 20660 83360 22150
rect 83270 20650 83360 20660
rect -1020 20580 -930 20590
rect 83270 20590 83280 20650
rect 83350 20590 83360 20650
rect 83270 20580 83360 20590
rect -1010 20510 -930 20520
rect -1010 20450 -1000 20510
rect -940 20450 -930 20510
rect -1010 20440 -930 20450
rect 83280 20510 83360 20520
rect 83280 20450 83290 20510
rect 83350 20450 83360 20510
rect 83280 20440 83360 20450
rect -4720 20400 -2000 20410
rect -4720 20382 -2070 20400
rect -4720 18958 -3032 20382
rect -2968 20350 -2070 20382
rect -2968 18958 -2948 20350
rect -2080 20340 -2070 20350
rect -2010 20340 -2000 20400
rect -2080 20320 -2000 20340
rect -1580 19760 -1440 19800
rect -1580 19690 -1550 19760
rect -1470 19690 -1440 19760
rect -1580 19650 -1440 19690
rect -1580 19580 -1550 19650
rect -1470 19580 -1440 19650
rect -1580 19550 -1440 19580
rect -4720 18930 -2948 18958
rect -990 18950 -930 20440
rect -1020 18940 -930 18950
rect -1020 18880 -1010 18940
rect -940 18880 -930 18940
rect 79570 20400 82290 20410
rect 79570 20382 82220 20400
rect 79570 18958 81258 20382
rect 81322 20350 82220 20382
rect 81322 18958 81342 20350
rect 82210 20340 82220 20350
rect 82280 20340 82290 20400
rect 82210 20320 82290 20340
rect 82710 19760 82850 19800
rect 82710 19690 82740 19760
rect 82820 19690 82850 19760
rect 82710 19650 82850 19690
rect 82710 19580 82740 19650
rect 82820 19580 82850 19650
rect 82710 19550 82850 19580
rect 79570 18930 81342 18958
rect 83300 18950 83360 20440
rect 83270 18940 83360 18950
rect -1020 18870 -930 18880
rect 83270 18880 83280 18940
rect 83350 18880 83360 18940
rect 83270 18870 83360 18880
rect -1010 18800 -930 18810
rect -1010 18740 -1000 18800
rect -940 18740 -930 18800
rect -1010 18730 -930 18740
rect 83280 18800 83360 18810
rect 83280 18740 83290 18800
rect 83350 18740 83360 18800
rect 83280 18730 83360 18740
rect -4720 18690 -2000 18700
rect -4720 18672 -2070 18690
rect -4720 17248 -3032 18672
rect -2968 18640 -2070 18672
rect -2968 17248 -2948 18640
rect -2080 18630 -2070 18640
rect -2010 18630 -2000 18690
rect -2080 18610 -2000 18630
rect -1580 18050 -1440 18090
rect -1580 17980 -1550 18050
rect -1470 17980 -1440 18050
rect -1580 17940 -1440 17980
rect -1580 17870 -1550 17940
rect -1470 17870 -1440 17940
rect -1580 17840 -1440 17870
rect -4720 17220 -2948 17248
rect -990 17240 -930 18730
rect -1020 17230 -930 17240
rect -1020 17170 -1010 17230
rect -940 17170 -930 17230
rect 79570 18690 82290 18700
rect 79570 18672 82220 18690
rect 79570 17248 81258 18672
rect 81322 18640 82220 18672
rect 81322 17248 81342 18640
rect 82210 18630 82220 18640
rect 82280 18630 82290 18690
rect 82210 18610 82290 18630
rect 82710 18050 82850 18090
rect 82710 17980 82740 18050
rect 82820 17980 82850 18050
rect 82710 17940 82850 17980
rect 82710 17870 82740 17940
rect 82820 17870 82850 17940
rect 82710 17840 82850 17870
rect 79570 17220 81342 17248
rect 83300 17240 83360 18730
rect 83270 17230 83360 17240
rect -1020 17160 -930 17170
rect 83270 17170 83280 17230
rect 83350 17170 83360 17230
rect 83270 17160 83360 17170
rect -1010 17090 -930 17100
rect -1010 17030 -1000 17090
rect -940 17030 -930 17090
rect -1010 17020 -930 17030
rect 83280 17090 83360 17100
rect 83280 17030 83290 17090
rect 83350 17030 83360 17090
rect 83280 17020 83360 17030
rect -4720 16980 -2000 16990
rect -4720 16962 -2070 16980
rect -4720 15538 -3032 16962
rect -2968 16930 -2070 16962
rect -2968 15538 -2948 16930
rect -2080 16920 -2070 16930
rect -2010 16920 -2000 16980
rect -2080 16900 -2000 16920
rect -1580 16340 -1440 16380
rect -1580 16270 -1550 16340
rect -1470 16270 -1440 16340
rect -1580 16230 -1440 16270
rect -1580 16160 -1550 16230
rect -1470 16160 -1440 16230
rect -1580 16130 -1440 16160
rect -4720 15510 -2948 15538
rect -990 15530 -930 17020
rect -1020 15520 -930 15530
rect -1020 15460 -1010 15520
rect -940 15460 -930 15520
rect 79570 16980 82290 16990
rect 79570 16962 82220 16980
rect 79570 15538 81258 16962
rect 81322 16930 82220 16962
rect 81322 15538 81342 16930
rect 82210 16920 82220 16930
rect 82280 16920 82290 16980
rect 82210 16900 82290 16920
rect 82710 16340 82850 16380
rect 82710 16270 82740 16340
rect 82820 16270 82850 16340
rect 82710 16230 82850 16270
rect 82710 16160 82740 16230
rect 82820 16160 82850 16230
rect 82710 16130 82850 16160
rect 79570 15510 81342 15538
rect 83300 15530 83360 17020
rect 83270 15520 83360 15530
rect -1020 15450 -930 15460
rect 83270 15460 83280 15520
rect 83350 15460 83360 15520
rect 83270 15450 83360 15460
rect -1010 15380 -930 15390
rect -1010 15320 -1000 15380
rect -940 15320 -930 15380
rect -1010 15310 -930 15320
rect 83280 15380 83360 15390
rect 83280 15320 83290 15380
rect 83350 15320 83360 15380
rect 83280 15310 83360 15320
rect -4720 15270 -2000 15280
rect -4720 15252 -2070 15270
rect -4720 13828 -3032 15252
rect -2968 15220 -2070 15252
rect -2968 13828 -2948 15220
rect -2080 15210 -2070 15220
rect -2010 15210 -2000 15270
rect -2080 15190 -2000 15210
rect -1580 14630 -1440 14670
rect -1580 14560 -1550 14630
rect -1470 14560 -1440 14630
rect -1580 14520 -1440 14560
rect -1580 14450 -1550 14520
rect -1470 14450 -1440 14520
rect -1580 14420 -1440 14450
rect -4720 13800 -2948 13828
rect -990 13820 -930 15310
rect -1020 13810 -930 13820
rect -1020 13750 -1010 13810
rect -940 13750 -930 13810
rect 79570 15270 82290 15280
rect 79570 15252 82220 15270
rect 79570 13828 81258 15252
rect 81322 15220 82220 15252
rect 81322 13828 81342 15220
rect 82210 15210 82220 15220
rect 82280 15210 82290 15270
rect 82210 15190 82290 15210
rect 82710 14630 82850 14670
rect 82710 14560 82740 14630
rect 82820 14560 82850 14630
rect 82710 14520 82850 14560
rect 82710 14450 82740 14520
rect 82820 14450 82850 14520
rect 82710 14420 82850 14450
rect 79570 13800 81342 13828
rect 83300 13820 83360 15310
rect 83270 13810 83360 13820
rect -1020 13740 -930 13750
rect 83270 13750 83280 13810
rect 83350 13750 83360 13810
rect 83270 13740 83360 13750
rect -1010 13670 -930 13680
rect -1010 13610 -1000 13670
rect -940 13610 -930 13670
rect -1010 13600 -930 13610
rect 83280 13670 83360 13680
rect 83280 13610 83290 13670
rect 83350 13610 83360 13670
rect 83280 13600 83360 13610
rect -4720 13560 -2000 13570
rect -4720 13542 -2070 13560
rect -4720 12118 -3032 13542
rect -2968 13510 -2070 13542
rect -2968 12118 -2948 13510
rect -2080 13500 -2070 13510
rect -2010 13500 -2000 13560
rect -2080 13480 -2000 13500
rect -1580 12920 -1440 12960
rect -1580 12850 -1550 12920
rect -1470 12850 -1440 12920
rect -1580 12810 -1440 12850
rect -1580 12740 -1550 12810
rect -1470 12740 -1440 12810
rect -1580 12710 -1440 12740
rect -4720 12090 -2948 12118
rect -990 12110 -930 13600
rect -1020 12100 -930 12110
rect -1020 12040 -1010 12100
rect -940 12040 -930 12100
rect 79570 13560 82290 13570
rect 79570 13542 82220 13560
rect 79570 12118 81258 13542
rect 81322 13510 82220 13542
rect 81322 12118 81342 13510
rect 82210 13500 82220 13510
rect 82280 13500 82290 13560
rect 82210 13480 82290 13500
rect 82710 12920 82850 12960
rect 82710 12850 82740 12920
rect 82820 12850 82850 12920
rect 82710 12810 82850 12850
rect 82710 12740 82740 12810
rect 82820 12740 82850 12810
rect 82710 12710 82850 12740
rect 79570 12090 81342 12118
rect 83300 12110 83360 13600
rect 83270 12100 83360 12110
rect -1020 12030 -930 12040
rect 83270 12040 83280 12100
rect 83350 12040 83360 12100
rect 83270 12030 83360 12040
rect -1010 11960 -930 11970
rect -1010 11900 -1000 11960
rect -940 11900 -930 11960
rect -1010 11890 -930 11900
rect 83280 11960 83360 11970
rect 83280 11900 83290 11960
rect 83350 11900 83360 11960
rect 83280 11890 83360 11900
rect -4720 11850 -2000 11860
rect -4720 11832 -2070 11850
rect -4720 10408 -3032 11832
rect -2968 11800 -2070 11832
rect -2968 10408 -2948 11800
rect -2080 11790 -2070 11800
rect -2010 11790 -2000 11850
rect -2080 11770 -2000 11790
rect -1580 11210 -1440 11250
rect -1580 11140 -1550 11210
rect -1470 11140 -1440 11210
rect -1580 11100 -1440 11140
rect -1580 11030 -1550 11100
rect -1470 11030 -1440 11100
rect -1580 11000 -1440 11030
rect -4720 10380 -2948 10408
rect -990 10400 -930 11890
rect -1020 10390 -930 10400
rect -1020 10330 -1010 10390
rect -940 10330 -930 10390
rect 79570 11850 82290 11860
rect 79570 11832 82220 11850
rect 79570 10408 81258 11832
rect 81322 11800 82220 11832
rect 81322 10408 81342 11800
rect 82210 11790 82220 11800
rect 82280 11790 82290 11850
rect 82210 11770 82290 11790
rect 82710 11210 82850 11250
rect 82710 11140 82740 11210
rect 82820 11140 82850 11210
rect 82710 11100 82850 11140
rect 82710 11030 82740 11100
rect 82820 11030 82850 11100
rect 82710 11000 82850 11030
rect 79570 10380 81342 10408
rect 83300 10400 83360 11890
rect 83270 10390 83360 10400
rect -1020 10320 -930 10330
rect 83270 10330 83280 10390
rect 83350 10330 83360 10390
rect 83270 10320 83360 10330
rect -1010 10250 -930 10260
rect -1010 10190 -1000 10250
rect -940 10190 -930 10250
rect -1010 10180 -930 10190
rect 83280 10250 83360 10260
rect 83280 10190 83290 10250
rect 83350 10190 83360 10250
rect 83280 10180 83360 10190
rect -4720 10140 -2000 10150
rect -4720 10122 -2070 10140
rect -4720 8698 -3032 10122
rect -2968 10090 -2070 10122
rect -2968 8698 -2948 10090
rect -2080 10080 -2070 10090
rect -2010 10080 -2000 10140
rect -2080 10060 -2000 10080
rect -1580 9500 -1440 9540
rect -1580 9430 -1550 9500
rect -1470 9430 -1440 9500
rect -1580 9390 -1440 9430
rect -1580 9320 -1550 9390
rect -1470 9320 -1440 9390
rect -1580 9290 -1440 9320
rect -4720 8670 -2948 8698
rect -990 8690 -930 10180
rect -1020 8680 -930 8690
rect -1020 8620 -1010 8680
rect -940 8620 -930 8680
rect 79570 10140 82290 10150
rect 79570 10122 82220 10140
rect 79570 8698 81258 10122
rect 81322 10090 82220 10122
rect 81322 8698 81342 10090
rect 82210 10080 82220 10090
rect 82280 10080 82290 10140
rect 82210 10060 82290 10080
rect 82710 9500 82850 9540
rect 82710 9430 82740 9500
rect 82820 9430 82850 9500
rect 82710 9390 82850 9430
rect 82710 9320 82740 9390
rect 82820 9320 82850 9390
rect 82710 9290 82850 9320
rect 79570 8670 81342 8698
rect 83300 8690 83360 10180
rect 83270 8680 83360 8690
rect -1020 8610 -930 8620
rect 83270 8620 83280 8680
rect 83350 8620 83360 8680
rect 83270 8610 83360 8620
rect -1010 8540 -930 8550
rect -1010 8480 -1000 8540
rect -940 8480 -930 8540
rect -1010 8470 -930 8480
rect 83280 8540 83360 8550
rect 83280 8480 83290 8540
rect 83350 8480 83360 8540
rect 83280 8470 83360 8480
rect -4720 8430 -2000 8440
rect -4720 8412 -2070 8430
rect -4720 6988 -3032 8412
rect -2968 8380 -2070 8412
rect -2968 6988 -2948 8380
rect -2080 8370 -2070 8380
rect -2010 8370 -2000 8430
rect -2080 8350 -2000 8370
rect -1580 7790 -1440 7830
rect -1580 7720 -1550 7790
rect -1470 7720 -1440 7790
rect -1580 7680 -1440 7720
rect -1580 7610 -1550 7680
rect -1470 7610 -1440 7680
rect -1580 7580 -1440 7610
rect -4720 6960 -2948 6988
rect -990 6980 -930 8470
rect -1020 6970 -930 6980
rect -1020 6910 -1010 6970
rect -940 6910 -930 6970
rect 79570 8430 82290 8440
rect 79570 8412 82220 8430
rect 79570 6988 81258 8412
rect 81322 8380 82220 8412
rect 81322 6988 81342 8380
rect 82210 8370 82220 8380
rect 82280 8370 82290 8430
rect 82210 8350 82290 8370
rect 82710 7790 82850 7830
rect 82710 7720 82740 7790
rect 82820 7720 82850 7790
rect 82710 7680 82850 7720
rect 82710 7610 82740 7680
rect 82820 7610 82850 7680
rect 82710 7580 82850 7610
rect 79570 6960 81342 6988
rect 83300 6980 83360 8470
rect 83270 6970 83360 6980
rect -1020 6900 -930 6910
rect 83270 6910 83280 6970
rect 83350 6910 83360 6970
rect 83270 6900 83360 6910
rect -1010 6830 -930 6840
rect -1010 6770 -1000 6830
rect -940 6770 -930 6830
rect -1010 6760 -930 6770
rect 83280 6830 83360 6840
rect 83280 6770 83290 6830
rect 83350 6770 83360 6830
rect 83280 6760 83360 6770
rect -4720 6720 -2000 6730
rect -4720 6702 -2070 6720
rect -4720 5278 -3032 6702
rect -2968 6670 -2070 6702
rect -2968 5278 -2948 6670
rect -2080 6660 -2070 6670
rect -2010 6660 -2000 6720
rect -2080 6640 -2000 6660
rect -1580 6080 -1440 6120
rect -1580 6010 -1550 6080
rect -1470 6010 -1440 6080
rect -1580 5970 -1440 6010
rect -1580 5900 -1550 5970
rect -1470 5900 -1440 5970
rect -1580 5870 -1440 5900
rect -4720 5250 -2948 5278
rect -990 5270 -930 6760
rect -1020 5260 -930 5270
rect -1020 5200 -1010 5260
rect -940 5200 -930 5260
rect 79570 6720 82290 6730
rect 79570 6702 82220 6720
rect 79570 5278 81258 6702
rect 81322 6670 82220 6702
rect 81322 5278 81342 6670
rect 82210 6660 82220 6670
rect 82280 6660 82290 6720
rect 82210 6640 82290 6660
rect 82710 6080 82850 6120
rect 82710 6010 82740 6080
rect 82820 6010 82850 6080
rect 82710 5970 82850 6010
rect 82710 5900 82740 5970
rect 82820 5900 82850 5970
rect 82710 5870 82850 5900
rect 79570 5250 81342 5278
rect 83300 5270 83360 6760
rect 83270 5260 83360 5270
rect -1020 5190 -930 5200
rect 83270 5200 83280 5260
rect 83350 5200 83360 5260
rect 83270 5190 83360 5200
rect -1010 5120 -930 5130
rect -1010 5060 -1000 5120
rect -940 5060 -930 5120
rect -1010 5050 -930 5060
rect 83280 5120 83360 5130
rect 83280 5060 83290 5120
rect 83350 5060 83360 5120
rect 83280 5050 83360 5060
rect -4720 5010 -2000 5020
rect -4720 4992 -2070 5010
rect -4720 3568 -3032 4992
rect -2968 4960 -2070 4992
rect -2968 3568 -2948 4960
rect -2080 4950 -2070 4960
rect -2010 4950 -2000 5010
rect -2080 4930 -2000 4950
rect -1580 4370 -1440 4410
rect -1580 4300 -1550 4370
rect -1470 4300 -1440 4370
rect -1580 4260 -1440 4300
rect -1580 4190 -1550 4260
rect -1470 4190 -1440 4260
rect -1580 4160 -1440 4190
rect -4720 3540 -2948 3568
rect -990 3560 -930 5050
rect -1020 3550 -930 3560
rect -1020 3490 -1010 3550
rect -940 3490 -930 3550
rect 79570 5010 82290 5020
rect 79570 4992 82220 5010
rect 79570 3568 81258 4992
rect 81322 4960 82220 4992
rect 81322 3568 81342 4960
rect 82210 4950 82220 4960
rect 82280 4950 82290 5010
rect 82210 4930 82290 4950
rect 82710 4370 82850 4410
rect 82710 4300 82740 4370
rect 82820 4300 82850 4370
rect 82710 4260 82850 4300
rect 82710 4190 82740 4260
rect 82820 4190 82850 4260
rect 82710 4160 82850 4190
rect 79570 3540 81342 3568
rect 83300 3560 83360 5050
rect 83270 3550 83360 3560
rect -1020 3480 -930 3490
rect 83270 3490 83280 3550
rect 83350 3490 83360 3550
rect 83270 3480 83360 3490
rect -1010 3410 -930 3420
rect -1010 3350 -1000 3410
rect -940 3350 -930 3410
rect -1010 3340 -930 3350
rect 83280 3410 83360 3420
rect 83280 3350 83290 3410
rect 83350 3350 83360 3410
rect 83280 3340 83360 3350
rect -4720 3300 -2000 3310
rect -4720 3282 -2070 3300
rect -4720 1858 -3032 3282
rect -2968 3250 -2070 3282
rect -2968 1858 -2948 3250
rect -2080 3240 -2070 3250
rect -2010 3240 -2000 3300
rect -2080 3220 -2000 3240
rect -1580 2660 -1440 2700
rect -1580 2590 -1550 2660
rect -1470 2590 -1440 2660
rect -1580 2550 -1440 2590
rect -1580 2480 -1550 2550
rect -1470 2480 -1440 2550
rect -1580 2450 -1440 2480
rect -4720 1830 -2948 1858
rect -990 1850 -930 3340
rect -1020 1840 -930 1850
rect -1020 1780 -1010 1840
rect -940 1780 -930 1840
rect 79570 3300 82290 3310
rect 79570 3282 82220 3300
rect 79570 1858 81258 3282
rect 81322 3250 82220 3282
rect 81322 1858 81342 3250
rect 82210 3240 82220 3250
rect 82280 3240 82290 3300
rect 82210 3220 82290 3240
rect 82710 2660 82850 2700
rect 82710 2590 82740 2660
rect 82820 2590 82850 2660
rect 82710 2550 82850 2590
rect 82710 2480 82740 2550
rect 82820 2480 82850 2550
rect 82710 2450 82850 2480
rect 79570 1830 81342 1858
rect 83300 1850 83360 3340
rect 83270 1840 83360 1850
rect -1020 1770 -930 1780
rect 83270 1780 83280 1840
rect 83350 1780 83360 1840
rect 83270 1770 83360 1780
rect -1010 1700 -930 1710
rect -1010 1640 -1000 1700
rect -940 1640 -930 1700
rect -1010 1630 -930 1640
rect 83280 1700 83360 1710
rect 83280 1640 83290 1700
rect 83350 1640 83360 1700
rect 83280 1630 83360 1640
rect -4720 1590 -2000 1600
rect -4720 1572 -2070 1590
rect -4720 148 -3032 1572
rect -2968 1540 -2070 1572
rect -2968 148 -2948 1540
rect -2080 1530 -2070 1540
rect -2010 1530 -2000 1590
rect -2080 1510 -2000 1530
rect -1580 950 -1440 990
rect -1580 880 -1550 950
rect -1470 880 -1440 950
rect -1580 840 -1440 880
rect -1580 770 -1550 840
rect -1470 770 -1440 840
rect -1580 740 -1440 770
rect -4720 120 -2948 148
rect -2080 140 -2000 150
rect -990 140 -930 1630
rect 79570 1590 82290 1600
rect 79570 1572 82220 1590
rect -2080 80 -2070 140
rect -2010 80 -2000 140
rect -2080 70 -2000 80
rect -1020 130 -930 140
rect -1020 70 -1010 130
rect -940 70 -930 130
rect 2640 140 2720 150
rect 2640 80 2650 140
rect 2710 130 2720 140
rect 7630 140 7710 150
rect 2710 80 3940 130
rect 2640 70 3940 80
rect 7630 80 7640 140
rect 7700 130 7710 140
rect 12620 140 12700 150
rect 7700 80 8930 130
rect 7630 70 8930 80
rect 12620 80 12630 140
rect 12690 130 12700 140
rect 17610 140 17690 150
rect 12690 80 13920 130
rect 12620 70 13920 80
rect 17610 80 17620 140
rect 17680 130 17690 140
rect 22600 140 22680 150
rect 17680 80 18910 130
rect 17610 70 18910 80
rect 22600 80 22610 140
rect 22670 130 22680 140
rect 27590 140 27670 150
rect 22670 80 23900 130
rect 22600 70 23900 80
rect 27590 80 27600 140
rect 27660 130 27670 140
rect 32580 140 32660 150
rect 27660 80 28890 130
rect 27590 70 28890 80
rect 32580 80 32590 140
rect 32650 130 32660 140
rect 37570 140 37650 150
rect 32650 80 33880 130
rect 32580 70 33880 80
rect 37570 80 37580 140
rect 37640 130 37650 140
rect 42560 140 42640 150
rect 37640 80 38870 130
rect 37570 70 38870 80
rect 42560 80 42570 140
rect 42630 130 42640 140
rect 47550 140 47630 150
rect 42630 80 43860 130
rect 42560 70 43860 80
rect 47550 80 47560 140
rect 47620 130 47630 140
rect 52540 140 52620 150
rect 47620 80 48850 130
rect 47550 70 48850 80
rect 52540 80 52550 140
rect 52610 130 52620 140
rect 57530 140 57610 150
rect 52610 80 53840 130
rect 52540 70 53840 80
rect 57530 80 57540 140
rect 57600 130 57610 140
rect 62520 140 62600 150
rect 57600 80 58830 130
rect 57530 70 58830 80
rect 62520 80 62530 140
rect 62590 130 62600 140
rect 67510 140 67590 150
rect 62590 80 63820 130
rect 62520 70 63820 80
rect 67510 80 67520 140
rect 67580 130 67590 140
rect 72500 140 72580 150
rect 67580 80 68810 130
rect 67510 70 68810 80
rect 72500 80 72510 140
rect 72570 130 72580 140
rect 77490 140 77570 150
rect 72570 80 73800 130
rect 72500 70 73800 80
rect 77490 80 77500 140
rect 77560 80 77570 140
rect 79570 148 81258 1572
rect 81322 1540 82220 1572
rect 81322 148 81342 1540
rect 82210 1530 82220 1540
rect 82280 1530 82290 1590
rect 82210 1510 82290 1530
rect 82710 950 82850 990
rect 82710 880 82740 950
rect 82820 880 82850 950
rect 82710 840 82850 880
rect 82710 770 82740 840
rect 82820 770 82850 840
rect 82710 740 82850 770
rect 79570 120 81342 148
rect 82210 140 82290 150
rect 83300 140 83360 1630
rect 77490 70 77570 80
rect 82210 80 82220 140
rect 82280 80 82290 140
rect 82210 70 82290 80
rect 83270 130 83360 140
rect 83270 70 83280 130
rect 83350 70 83360 130
rect -2880 -30 -1970 70
rect -1020 60 -930 70
rect -2860 -50 -1970 -30
rect -1010 -10 -930 0
rect -1010 -70 -1000 -10
rect -940 -70 -930 -10
rect 1840 -30 2750 70
rect 3850 40 4750 70
rect 1860 -50 2750 -30
rect 3710 -10 3790 0
rect -1010 -80 -930 -70
rect 3710 -70 3720 -10
rect 3780 -70 3790 -10
rect 3850 -20 3860 40
rect 3920 -20 4750 40
rect 3850 -50 4750 -20
rect 6830 -30 7740 70
rect 8840 40 9740 70
rect 6850 -50 7740 -30
rect 8700 -10 8780 0
rect 3710 -80 3790 -70
rect 8700 -70 8710 -10
rect 8770 -70 8780 -10
rect 8840 -20 8850 40
rect 8910 -20 9740 40
rect 8840 -50 9740 -20
rect 11820 -30 12730 70
rect 13830 40 14730 70
rect 11840 -50 12730 -30
rect 13690 -10 13770 0
rect 8700 -80 8780 -70
rect 13690 -70 13700 -10
rect 13760 -70 13770 -10
rect 13830 -20 13840 40
rect 13900 -20 14730 40
rect 13830 -50 14730 -20
rect 16810 -30 17720 70
rect 18820 40 19720 70
rect 16830 -50 17720 -30
rect 18680 -10 18760 0
rect 13690 -80 13770 -70
rect 18680 -70 18690 -10
rect 18750 -70 18760 -10
rect 18820 -20 18830 40
rect 18890 -20 19720 40
rect 18820 -50 19720 -20
rect 21800 -30 22710 70
rect 23810 40 24710 70
rect 21820 -50 22710 -30
rect 23670 -10 23750 0
rect 18680 -80 18760 -70
rect 23670 -70 23680 -10
rect 23740 -70 23750 -10
rect 23810 -20 23820 40
rect 23880 -20 24710 40
rect 23810 -50 24710 -20
rect 26790 -30 27700 70
rect 28800 40 29700 70
rect 26810 -50 27700 -30
rect 28660 -10 28740 0
rect 23670 -80 23750 -70
rect 28660 -70 28670 -10
rect 28730 -70 28740 -10
rect 28800 -20 28810 40
rect 28870 -20 29700 40
rect 28800 -50 29700 -20
rect 31780 -30 32690 70
rect 33790 40 34690 70
rect 31800 -50 32690 -30
rect 33650 -10 33730 0
rect 28660 -80 28740 -70
rect 33650 -70 33660 -10
rect 33720 -70 33730 -10
rect 33790 -20 33800 40
rect 33860 -20 34690 40
rect 33790 -50 34690 -20
rect 36770 -30 37680 70
rect 38780 40 39680 70
rect 36790 -50 37680 -30
rect 38640 -10 38720 0
rect 33650 -80 33730 -70
rect 38640 -70 38650 -10
rect 38710 -70 38720 -10
rect 38780 -20 38790 40
rect 38850 -20 39680 40
rect 38780 -50 39680 -20
rect 41760 -30 42670 70
rect 43770 40 44670 70
rect 41780 -50 42670 -30
rect 43630 -10 43710 0
rect 38640 -80 38720 -70
rect 43630 -70 43640 -10
rect 43700 -70 43710 -10
rect 43770 -20 43780 40
rect 43840 -20 44670 40
rect 43770 -50 44670 -20
rect 46750 -30 47660 70
rect 48760 40 49660 70
rect 46770 -50 47660 -30
rect 48620 -10 48700 0
rect 43630 -80 43710 -70
rect 48620 -70 48630 -10
rect 48690 -70 48700 -10
rect 48760 -20 48770 40
rect 48830 -20 49660 40
rect 48760 -50 49660 -20
rect 51740 -30 52650 70
rect 53750 40 54650 70
rect 51760 -50 52650 -30
rect 53610 -10 53690 0
rect 48620 -80 48700 -70
rect 53610 -70 53620 -10
rect 53680 -70 53690 -10
rect 53750 -20 53760 40
rect 53820 -20 54650 40
rect 53750 -50 54650 -20
rect 56730 -30 57640 70
rect 58740 40 59640 70
rect 56750 -50 57640 -30
rect 58600 -10 58680 0
rect 53610 -80 53690 -70
rect 58600 -70 58610 -10
rect 58670 -70 58680 -10
rect 58740 -20 58750 40
rect 58810 -20 59640 40
rect 58740 -50 59640 -20
rect 61720 -30 62630 70
rect 63730 40 64630 70
rect 61740 -50 62630 -30
rect 63590 -10 63670 0
rect 58600 -80 58680 -70
rect 63590 -70 63600 -10
rect 63660 -70 63670 -10
rect 63730 -20 63740 40
rect 63800 -20 64630 40
rect 63730 -50 64630 -20
rect 66710 -30 67620 70
rect 68720 40 69620 70
rect 66730 -50 67620 -30
rect 68580 -10 68660 0
rect 63590 -80 63670 -70
rect 68580 -70 68590 -10
rect 68650 -70 68660 -10
rect 68720 -20 68730 40
rect 68790 -20 69620 40
rect 68720 -50 69620 -20
rect 71700 -30 72610 70
rect 73710 40 74610 70
rect 71720 -50 72610 -30
rect 73570 -10 73650 0
rect 68580 -80 68660 -70
rect 73570 -70 73580 -10
rect 73640 -70 73650 -10
rect 73710 -20 73720 40
rect 73780 -20 74610 40
rect 73710 -50 74610 -20
rect 76690 -30 77600 70
rect 76710 -50 77600 -30
rect 78560 -10 78640 0
rect 73570 -80 73650 -70
rect 78560 -70 78570 -10
rect 78630 -70 78640 -10
rect 81410 -30 82320 70
rect 83270 60 83360 70
rect 81430 -50 82320 -30
rect 83280 -10 83360 0
rect 78560 -80 78640 -70
rect 83280 -70 83290 -10
rect 83350 -70 83360 -10
rect 83280 -80 83360 -70
rect -4720 -120 -2000 -110
rect -4720 -138 -2070 -120
rect -4720 -1562 -3032 -138
rect -2968 -170 -2070 -138
rect -2968 -1562 -2948 -170
rect -2080 -180 -2070 -170
rect -2010 -180 -2000 -120
rect -2080 -200 -2000 -180
rect -1580 -760 -1440 -720
rect -1580 -830 -1550 -760
rect -1470 -830 -1440 -760
rect -1580 -870 -1440 -830
rect -1580 -940 -1550 -870
rect -1470 -940 -1440 -870
rect -1580 -970 -1440 -940
rect -4720 -1590 -2948 -1562
rect -990 -1570 -930 -80
rect -1020 -1580 -930 -1570
rect -1020 -1640 -1010 -1580
rect -940 -1640 -930 -1580
rect 0 -120 2720 -110
rect 0 -138 2650 -120
rect 0 -1562 1688 -138
rect 1752 -170 2650 -138
rect 1752 -1562 1772 -170
rect 2640 -180 2650 -170
rect 2710 -180 2720 -120
rect 2640 -200 2720 -180
rect 3140 -760 3280 -720
rect 3140 -830 3170 -760
rect 3250 -830 3280 -760
rect 3140 -870 3280 -830
rect 3140 -940 3170 -870
rect 3250 -940 3280 -870
rect 3140 -970 3280 -940
rect 0 -1590 1772 -1562
rect 3730 -1630 3790 -80
rect 4990 -120 7710 -110
rect 4990 -138 7640 -120
rect 4990 -1562 6678 -138
rect 6742 -170 7640 -138
rect 6742 -1562 6762 -170
rect 7630 -180 7640 -170
rect 7700 -180 7710 -120
rect 7630 -200 7710 -180
rect 8130 -760 8270 -720
rect 8130 -830 8160 -760
rect 8240 -830 8270 -760
rect 8130 -870 8270 -830
rect 8130 -940 8160 -870
rect 8240 -940 8270 -870
rect 8130 -970 8270 -940
rect 4990 -1590 6762 -1562
rect 8720 -1630 8780 -80
rect 9980 -120 12700 -110
rect 9980 -138 12630 -120
rect 9980 -1562 11668 -138
rect 11732 -170 12630 -138
rect 11732 -1562 11752 -170
rect 12620 -180 12630 -170
rect 12690 -180 12700 -120
rect 12620 -200 12700 -180
rect 13120 -760 13260 -720
rect 13120 -830 13150 -760
rect 13230 -830 13260 -760
rect 13120 -870 13260 -830
rect 13120 -940 13150 -870
rect 13230 -940 13260 -870
rect 13120 -970 13260 -940
rect 9980 -1590 11752 -1562
rect 13710 -1630 13770 -80
rect 14970 -120 17690 -110
rect 14970 -138 17620 -120
rect 14970 -1562 16658 -138
rect 16722 -170 17620 -138
rect 16722 -1562 16742 -170
rect 17610 -180 17620 -170
rect 17680 -180 17690 -120
rect 17610 -200 17690 -180
rect 18110 -760 18250 -720
rect 18110 -830 18140 -760
rect 18220 -830 18250 -760
rect 18110 -870 18250 -830
rect 18110 -940 18140 -870
rect 18220 -940 18250 -870
rect 18110 -970 18250 -940
rect 14970 -1590 16742 -1562
rect 18700 -1630 18760 -80
rect 19960 -120 22680 -110
rect 19960 -138 22610 -120
rect 19960 -1562 21648 -138
rect 21712 -170 22610 -138
rect 21712 -1562 21732 -170
rect 22600 -180 22610 -170
rect 22670 -180 22680 -120
rect 22600 -200 22680 -180
rect 23100 -760 23240 -720
rect 23100 -830 23130 -760
rect 23210 -830 23240 -760
rect 23100 -870 23240 -830
rect 23100 -940 23130 -870
rect 23210 -940 23240 -870
rect 23100 -970 23240 -940
rect 19960 -1590 21732 -1562
rect 23690 -1630 23750 -80
rect 24950 -120 27670 -110
rect 24950 -138 27600 -120
rect 24950 -1562 26638 -138
rect 26702 -170 27600 -138
rect 26702 -1562 26722 -170
rect 27590 -180 27600 -170
rect 27660 -180 27670 -120
rect 27590 -200 27670 -180
rect 28090 -760 28230 -720
rect 28090 -830 28120 -760
rect 28200 -830 28230 -760
rect 28090 -870 28230 -830
rect 28090 -940 28120 -870
rect 28200 -940 28230 -870
rect 28090 -970 28230 -940
rect 24950 -1590 26722 -1562
rect 28680 -1630 28740 -80
rect 29940 -120 32660 -110
rect 29940 -138 32590 -120
rect 29940 -1562 31628 -138
rect 31692 -170 32590 -138
rect 31692 -1562 31712 -170
rect 32580 -180 32590 -170
rect 32650 -180 32660 -120
rect 32580 -200 32660 -180
rect 33080 -760 33220 -720
rect 33080 -830 33110 -760
rect 33190 -830 33220 -760
rect 33080 -870 33220 -830
rect 33080 -940 33110 -870
rect 33190 -940 33220 -870
rect 33080 -970 33220 -940
rect 29940 -1590 31712 -1562
rect 33670 -1630 33730 -80
rect 34930 -120 37650 -110
rect 34930 -138 37580 -120
rect 34930 -1562 36618 -138
rect 36682 -170 37580 -138
rect 36682 -1562 36702 -170
rect 37570 -180 37580 -170
rect 37640 -180 37650 -120
rect 37570 -200 37650 -180
rect 38070 -760 38210 -720
rect 38070 -830 38100 -760
rect 38180 -830 38210 -760
rect 38070 -870 38210 -830
rect 38070 -940 38100 -870
rect 38180 -940 38210 -870
rect 38070 -970 38210 -940
rect 34930 -1590 36702 -1562
rect 38660 -1630 38720 -80
rect 39920 -120 42640 -110
rect 39920 -138 42570 -120
rect 39920 -1562 41608 -138
rect 41672 -170 42570 -138
rect 41672 -1562 41692 -170
rect 42560 -180 42570 -170
rect 42630 -180 42640 -120
rect 42560 -200 42640 -180
rect 43060 -760 43200 -720
rect 43060 -830 43090 -760
rect 43170 -830 43200 -760
rect 43060 -870 43200 -830
rect 43060 -940 43090 -870
rect 43170 -940 43200 -870
rect 43060 -970 43200 -940
rect 39920 -1590 41692 -1562
rect 43650 -1630 43710 -80
rect 44910 -120 47630 -110
rect 44910 -138 47560 -120
rect 44910 -1562 46598 -138
rect 46662 -170 47560 -138
rect 46662 -1562 46682 -170
rect 47550 -180 47560 -170
rect 47620 -180 47630 -120
rect 47550 -200 47630 -180
rect 48050 -760 48190 -720
rect 48050 -830 48080 -760
rect 48160 -830 48190 -760
rect 48050 -870 48190 -830
rect 48050 -940 48080 -870
rect 48160 -940 48190 -870
rect 48050 -970 48190 -940
rect 44910 -1590 46682 -1562
rect 48640 -1630 48700 -80
rect 49900 -120 52620 -110
rect 49900 -138 52550 -120
rect 49900 -1562 51588 -138
rect 51652 -170 52550 -138
rect 51652 -1562 51672 -170
rect 52540 -180 52550 -170
rect 52610 -180 52620 -120
rect 52540 -200 52620 -180
rect 53040 -760 53180 -720
rect 53040 -830 53070 -760
rect 53150 -830 53180 -760
rect 53040 -870 53180 -830
rect 53040 -940 53070 -870
rect 53150 -940 53180 -870
rect 53040 -970 53180 -940
rect 49900 -1590 51672 -1562
rect 53630 -1630 53690 -80
rect 54890 -120 57610 -110
rect 54890 -138 57540 -120
rect 54890 -1562 56578 -138
rect 56642 -170 57540 -138
rect 56642 -1562 56662 -170
rect 57530 -180 57540 -170
rect 57600 -180 57610 -120
rect 57530 -200 57610 -180
rect 58030 -760 58170 -720
rect 58030 -830 58060 -760
rect 58140 -830 58170 -760
rect 58030 -870 58170 -830
rect 58030 -940 58060 -870
rect 58140 -940 58170 -870
rect 58030 -970 58170 -940
rect 54890 -1590 56662 -1562
rect 58620 -1630 58680 -80
rect 59880 -120 62600 -110
rect 59880 -138 62530 -120
rect 59880 -1562 61568 -138
rect 61632 -170 62530 -138
rect 61632 -1562 61652 -170
rect 62520 -180 62530 -170
rect 62590 -180 62600 -120
rect 62520 -200 62600 -180
rect 63020 -760 63160 -720
rect 63020 -830 63050 -760
rect 63130 -830 63160 -760
rect 63020 -870 63160 -830
rect 63020 -940 63050 -870
rect 63130 -940 63160 -870
rect 63020 -970 63160 -940
rect 59880 -1590 61652 -1562
rect 63610 -1630 63670 -80
rect 64870 -120 67590 -110
rect 64870 -138 67520 -120
rect 64870 -1562 66558 -138
rect 66622 -170 67520 -138
rect 66622 -1562 66642 -170
rect 67510 -180 67520 -170
rect 67580 -180 67590 -120
rect 67510 -200 67590 -180
rect 68010 -760 68150 -720
rect 68010 -830 68040 -760
rect 68120 -830 68150 -760
rect 68010 -870 68150 -830
rect 68010 -940 68040 -870
rect 68120 -940 68150 -870
rect 68010 -970 68150 -940
rect 64870 -1590 66642 -1562
rect 68600 -1630 68660 -80
rect 69860 -120 72580 -110
rect 69860 -138 72510 -120
rect 69860 -1562 71548 -138
rect 71612 -170 72510 -138
rect 71612 -1562 71632 -170
rect 72500 -180 72510 -170
rect 72570 -180 72580 -120
rect 72500 -200 72580 -180
rect 73000 -760 73140 -720
rect 73000 -830 73030 -760
rect 73110 -830 73140 -760
rect 73000 -870 73140 -830
rect 73000 -940 73030 -870
rect 73110 -940 73140 -870
rect 73000 -970 73140 -940
rect 69860 -1590 71632 -1562
rect 73590 -1630 73650 -80
rect 74850 -120 77570 -110
rect 74850 -138 77500 -120
rect 74850 -1562 76538 -138
rect 76602 -170 77500 -138
rect 76602 -1562 76622 -170
rect 77490 -180 77500 -170
rect 77560 -180 77570 -120
rect 77490 -200 77570 -180
rect 77990 -760 78130 -720
rect 77990 -830 78020 -760
rect 78100 -830 78130 -760
rect 77990 -870 78130 -830
rect 77990 -940 78020 -870
rect 78100 -940 78130 -870
rect 77990 -970 78130 -940
rect 74850 -1590 76622 -1562
rect 78580 -1630 78640 -80
rect 79570 -120 82290 -110
rect 79570 -138 82220 -120
rect 79570 -1562 81258 -138
rect 81322 -170 82220 -138
rect 81322 -1562 81342 -170
rect 82210 -180 82220 -170
rect 82280 -180 82290 -120
rect 82210 -200 82290 -180
rect 82710 -760 82850 -720
rect 82710 -830 82740 -760
rect 82820 -830 82850 -760
rect 82710 -870 82850 -830
rect 82710 -940 82740 -870
rect 82820 -940 82850 -870
rect 82710 -970 82850 -940
rect 79570 -1590 81342 -1562
rect 83300 -1570 83360 -80
rect 83270 -1580 83360 -1570
rect -1020 -1650 -930 -1640
rect 3710 -1640 3790 -1630
rect 3710 -1700 3720 -1640
rect 3780 -1700 3790 -1640
rect 3710 -1710 3790 -1700
rect 8700 -1640 8780 -1630
rect 8700 -1700 8710 -1640
rect 8770 -1700 8780 -1640
rect 8700 -1710 8780 -1700
rect 13690 -1640 13770 -1630
rect 13690 -1700 13700 -1640
rect 13760 -1700 13770 -1640
rect 13690 -1710 13770 -1700
rect 18680 -1640 18760 -1630
rect 18680 -1700 18690 -1640
rect 18750 -1700 18760 -1640
rect 18680 -1710 18760 -1700
rect 23670 -1640 23750 -1630
rect 23670 -1700 23680 -1640
rect 23740 -1700 23750 -1640
rect 23670 -1710 23750 -1700
rect 28660 -1640 28740 -1630
rect 28660 -1700 28670 -1640
rect 28730 -1700 28740 -1640
rect 28660 -1710 28740 -1700
rect 33650 -1640 33730 -1630
rect 33650 -1700 33660 -1640
rect 33720 -1700 33730 -1640
rect 33650 -1710 33730 -1700
rect 38640 -1640 38720 -1630
rect 38640 -1700 38650 -1640
rect 38710 -1700 38720 -1640
rect 38640 -1710 38720 -1700
rect 43630 -1640 43710 -1630
rect 43630 -1700 43640 -1640
rect 43700 -1700 43710 -1640
rect 43630 -1710 43710 -1700
rect 48620 -1640 48700 -1630
rect 48620 -1700 48630 -1640
rect 48690 -1700 48700 -1640
rect 48620 -1710 48700 -1700
rect 53610 -1640 53690 -1630
rect 53610 -1700 53620 -1640
rect 53680 -1700 53690 -1640
rect 53610 -1710 53690 -1700
rect 58600 -1640 58680 -1630
rect 58600 -1700 58610 -1640
rect 58670 -1700 58680 -1640
rect 58600 -1710 58680 -1700
rect 63590 -1640 63670 -1630
rect 63590 -1700 63600 -1640
rect 63660 -1700 63670 -1640
rect 63590 -1710 63670 -1700
rect 68580 -1640 68660 -1630
rect 68580 -1700 68590 -1640
rect 68650 -1700 68660 -1640
rect 68580 -1710 68660 -1700
rect 73570 -1640 73650 -1630
rect 73570 -1700 73580 -1640
rect 73640 -1700 73650 -1640
rect 73570 -1710 73650 -1700
rect 78560 -1640 78640 -1630
rect 78560 -1700 78570 -1640
rect 78630 -1700 78640 -1640
rect 83270 -1640 83280 -1580
rect 83350 -1640 83360 -1580
rect 83270 -1650 83360 -1640
rect 78560 -1710 78640 -1700
<< via3 >>
rect -5520 30120 -5440 30130
rect -5520 30060 -5510 30120
rect -5510 30060 -5450 30120
rect -5450 30060 -5440 30120
rect -5520 30050 -5440 30060
rect 1688 27508 1752 28932
rect 3170 28240 3180 28310
rect 3180 28240 3250 28310
rect 3170 28130 3180 28200
rect 3180 28130 3250 28200
rect 6678 27508 6742 28932
rect 8160 28240 8170 28310
rect 8170 28240 8240 28310
rect 8160 28130 8170 28200
rect 8170 28130 8240 28200
rect 11668 27508 11732 28932
rect 13150 28240 13160 28310
rect 13160 28240 13230 28310
rect 13150 28130 13160 28200
rect 13160 28130 13230 28200
rect 16658 27508 16722 28932
rect 18140 28240 18150 28310
rect 18150 28240 18220 28310
rect 18140 28130 18150 28200
rect 18150 28130 18220 28200
rect 21648 27508 21712 28932
rect 23130 28240 23140 28310
rect 23140 28240 23210 28310
rect 23130 28130 23140 28200
rect 23140 28130 23210 28200
rect 26638 27508 26702 28932
rect 28120 28240 28130 28310
rect 28130 28240 28200 28310
rect 28120 28130 28130 28200
rect 28130 28130 28200 28200
rect 31628 27508 31692 28932
rect 33110 28240 33120 28310
rect 33120 28240 33190 28310
rect 33110 28130 33120 28200
rect 33120 28130 33190 28200
rect 36618 27508 36682 28932
rect 38100 28240 38110 28310
rect 38110 28240 38180 28310
rect 38100 28130 38110 28200
rect 38110 28130 38180 28200
rect 41608 27508 41672 28932
rect 43090 28240 43100 28310
rect 43100 28240 43170 28310
rect 43090 28130 43100 28200
rect 43100 28130 43170 28200
rect 46598 27508 46662 28932
rect 48080 28240 48090 28310
rect 48090 28240 48160 28310
rect 48080 28130 48090 28200
rect 48090 28130 48160 28200
rect 51588 27508 51652 28932
rect 53070 28240 53080 28310
rect 53080 28240 53150 28310
rect 53070 28130 53080 28200
rect 53080 28130 53150 28200
rect 56578 27508 56642 28932
rect 58060 28240 58070 28310
rect 58070 28240 58140 28310
rect 58060 28130 58070 28200
rect 58070 28130 58140 28200
rect 61568 27508 61632 28932
rect 63050 28240 63060 28310
rect 63060 28240 63130 28310
rect 63050 28130 63060 28200
rect 63060 28130 63130 28200
rect 66558 27508 66622 28932
rect 68040 28240 68050 28310
rect 68050 28240 68120 28310
rect 68040 28130 68050 28200
rect 68050 28130 68120 28200
rect 71548 27508 71612 28932
rect 73030 28240 73040 28310
rect 73040 28240 73110 28310
rect 73030 28130 73040 28200
rect 73040 28130 73110 28200
rect 76538 27508 76602 28932
rect 78020 28240 78030 28310
rect 78030 28240 78100 28310
rect 78020 28130 78030 28200
rect 78030 28130 78100 28200
rect 81258 27508 81322 28932
rect 82740 28240 82750 28310
rect 82750 28240 82820 28310
rect 82740 28130 82750 28200
rect 82750 28130 82820 28200
rect 81258 25798 81322 27222
rect 82740 26530 82750 26600
rect 82750 26530 82820 26600
rect 82740 26420 82750 26490
rect 82750 26420 82820 26490
rect 81258 24088 81322 25512
rect 82740 24820 82750 24890
rect 82750 24820 82820 24890
rect 82740 24710 82750 24780
rect 82750 24710 82820 24780
rect -3032 22378 -2968 23802
rect -1550 23110 -1540 23180
rect -1540 23110 -1470 23180
rect -1550 23000 -1540 23070
rect -1540 23000 -1470 23070
rect 81258 22378 81322 23802
rect 82740 23110 82750 23180
rect 82750 23110 82820 23180
rect 82740 23000 82750 23070
rect 82750 23000 82820 23070
rect -3032 20668 -2968 22092
rect -1550 21400 -1540 21470
rect -1540 21400 -1470 21470
rect -1550 21290 -1540 21360
rect -1540 21290 -1470 21360
rect 81258 20668 81322 22092
rect 82740 21400 82750 21470
rect 82750 21400 82820 21470
rect 82740 21290 82750 21360
rect 82750 21290 82820 21360
rect -3032 18958 -2968 20382
rect -1550 19690 -1540 19760
rect -1540 19690 -1470 19760
rect -1550 19580 -1540 19650
rect -1540 19580 -1470 19650
rect 81258 18958 81322 20382
rect 82740 19690 82750 19760
rect 82750 19690 82820 19760
rect 82740 19580 82750 19650
rect 82750 19580 82820 19650
rect -3032 17248 -2968 18672
rect -1550 17980 -1540 18050
rect -1540 17980 -1470 18050
rect -1550 17870 -1540 17940
rect -1540 17870 -1470 17940
rect 81258 17248 81322 18672
rect 82740 17980 82750 18050
rect 82750 17980 82820 18050
rect 82740 17870 82750 17940
rect 82750 17870 82820 17940
rect -3032 15538 -2968 16962
rect -1550 16270 -1540 16340
rect -1540 16270 -1470 16340
rect -1550 16160 -1540 16230
rect -1540 16160 -1470 16230
rect 81258 15538 81322 16962
rect 82740 16270 82750 16340
rect 82750 16270 82820 16340
rect 82740 16160 82750 16230
rect 82750 16160 82820 16230
rect -3032 13828 -2968 15252
rect -1550 14560 -1540 14630
rect -1540 14560 -1470 14630
rect -1550 14450 -1540 14520
rect -1540 14450 -1470 14520
rect 81258 13828 81322 15252
rect 82740 14560 82750 14630
rect 82750 14560 82820 14630
rect 82740 14450 82750 14520
rect 82750 14450 82820 14520
rect -3032 12118 -2968 13542
rect -1550 12850 -1540 12920
rect -1540 12850 -1470 12920
rect -1550 12740 -1540 12810
rect -1540 12740 -1470 12810
rect 81258 12118 81322 13542
rect 82740 12850 82750 12920
rect 82750 12850 82820 12920
rect 82740 12740 82750 12810
rect 82750 12740 82820 12810
rect -3032 10408 -2968 11832
rect -1550 11140 -1540 11210
rect -1540 11140 -1470 11210
rect -1550 11030 -1540 11100
rect -1540 11030 -1470 11100
rect 81258 10408 81322 11832
rect 82740 11140 82750 11210
rect 82750 11140 82820 11210
rect 82740 11030 82750 11100
rect 82750 11030 82820 11100
rect -3032 8698 -2968 10122
rect -1550 9430 -1540 9500
rect -1540 9430 -1470 9500
rect -1550 9320 -1540 9390
rect -1540 9320 -1470 9390
rect 81258 8698 81322 10122
rect 82740 9430 82750 9500
rect 82750 9430 82820 9500
rect 82740 9320 82750 9390
rect 82750 9320 82820 9390
rect -3032 6988 -2968 8412
rect -1550 7720 -1540 7790
rect -1540 7720 -1470 7790
rect -1550 7610 -1540 7680
rect -1540 7610 -1470 7680
rect 81258 6988 81322 8412
rect 82740 7720 82750 7790
rect 82750 7720 82820 7790
rect 82740 7610 82750 7680
rect 82750 7610 82820 7680
rect -3032 5278 -2968 6702
rect -1550 6010 -1540 6080
rect -1540 6010 -1470 6080
rect -1550 5900 -1540 5970
rect -1540 5900 -1470 5970
rect 81258 5278 81322 6702
rect 82740 6010 82750 6080
rect 82750 6010 82820 6080
rect 82740 5900 82750 5970
rect 82750 5900 82820 5970
rect -3032 3568 -2968 4992
rect -1550 4300 -1540 4370
rect -1540 4300 -1470 4370
rect -1550 4190 -1540 4260
rect -1540 4190 -1470 4260
rect 81258 3568 81322 4992
rect 82740 4300 82750 4370
rect 82750 4300 82820 4370
rect 82740 4190 82750 4260
rect 82750 4190 82820 4260
rect -3032 1858 -2968 3282
rect -1550 2590 -1540 2660
rect -1540 2590 -1470 2660
rect -1550 2480 -1540 2550
rect -1540 2480 -1470 2550
rect 81258 1858 81322 3282
rect 82740 2590 82750 2660
rect 82750 2590 82820 2660
rect 82740 2480 82750 2550
rect 82750 2480 82820 2550
rect -3032 148 -2968 1572
rect -1550 880 -1540 950
rect -1540 880 -1470 950
rect -1550 770 -1540 840
rect -1540 770 -1470 840
rect 81258 148 81322 1572
rect 82740 880 82750 950
rect 82750 880 82820 950
rect 82740 770 82750 840
rect 82750 770 82820 840
rect -3032 -1562 -2968 -138
rect -1550 -830 -1540 -760
rect -1540 -830 -1470 -760
rect -1550 -940 -1540 -870
rect -1540 -940 -1470 -870
rect 1688 -1562 1752 -138
rect 3170 -830 3180 -760
rect 3180 -830 3250 -760
rect 3170 -940 3180 -870
rect 3180 -940 3250 -870
rect 6678 -1562 6742 -138
rect 8160 -830 8170 -760
rect 8170 -830 8240 -760
rect 8160 -940 8170 -870
rect 8170 -940 8240 -870
rect 11668 -1562 11732 -138
rect 13150 -830 13160 -760
rect 13160 -830 13230 -760
rect 13150 -940 13160 -870
rect 13160 -940 13230 -870
rect 16658 -1562 16722 -138
rect 18140 -830 18150 -760
rect 18150 -830 18220 -760
rect 18140 -940 18150 -870
rect 18150 -940 18220 -870
rect 21648 -1562 21712 -138
rect 23130 -830 23140 -760
rect 23140 -830 23210 -760
rect 23130 -940 23140 -870
rect 23140 -940 23210 -870
rect 26638 -1562 26702 -138
rect 28120 -830 28130 -760
rect 28130 -830 28200 -760
rect 28120 -940 28130 -870
rect 28130 -940 28200 -870
rect 31628 -1562 31692 -138
rect 33110 -830 33120 -760
rect 33120 -830 33190 -760
rect 33110 -940 33120 -870
rect 33120 -940 33190 -870
rect 36618 -1562 36682 -138
rect 38100 -830 38110 -760
rect 38110 -830 38180 -760
rect 38100 -940 38110 -870
rect 38110 -940 38180 -870
rect 41608 -1562 41672 -138
rect 43090 -830 43100 -760
rect 43100 -830 43170 -760
rect 43090 -940 43100 -870
rect 43100 -940 43170 -870
rect 46598 -1562 46662 -138
rect 48080 -830 48090 -760
rect 48090 -830 48160 -760
rect 48080 -940 48090 -870
rect 48090 -940 48160 -870
rect 51588 -1562 51652 -138
rect 53070 -830 53080 -760
rect 53080 -830 53150 -760
rect 53070 -940 53080 -870
rect 53080 -940 53150 -870
rect 56578 -1562 56642 -138
rect 58060 -830 58070 -760
rect 58070 -830 58140 -760
rect 58060 -940 58070 -870
rect 58070 -940 58140 -870
rect 61568 -1562 61632 -138
rect 63050 -830 63060 -760
rect 63060 -830 63130 -760
rect 63050 -940 63060 -870
rect 63060 -940 63130 -870
rect 66558 -1562 66622 -138
rect 68040 -830 68050 -760
rect 68050 -830 68120 -760
rect 68040 -940 68050 -870
rect 68050 -940 68120 -870
rect 71548 -1562 71612 -138
rect 73030 -830 73040 -760
rect 73040 -830 73110 -760
rect 73030 -940 73040 -870
rect 73040 -940 73110 -870
rect 76538 -1562 76602 -138
rect 78020 -830 78030 -760
rect 78030 -830 78100 -760
rect 78020 -940 78030 -870
rect 78030 -940 78100 -870
rect 81258 -1562 81322 -138
rect 82740 -830 82750 -760
rect 82750 -830 82820 -760
rect 82740 -940 82750 -870
rect 82750 -940 82820 -870
<< mimcap >>
rect 40 28880 1440 28920
rect 40 27560 80 28880
rect 1400 27560 1440 28880
rect 40 27520 1440 27560
rect 5030 28880 6430 28920
rect 5030 27560 5070 28880
rect 6390 27560 6430 28880
rect 5030 27520 6430 27560
rect 10020 28880 11420 28920
rect 10020 27560 10060 28880
rect 11380 27560 11420 28880
rect 10020 27520 11420 27560
rect 15010 28880 16410 28920
rect 15010 27560 15050 28880
rect 16370 27560 16410 28880
rect 15010 27520 16410 27560
rect 20000 28880 21400 28920
rect 20000 27560 20040 28880
rect 21360 27560 21400 28880
rect 20000 27520 21400 27560
rect 24990 28880 26390 28920
rect 24990 27560 25030 28880
rect 26350 27560 26390 28880
rect 24990 27520 26390 27560
rect 29980 28880 31380 28920
rect 29980 27560 30020 28880
rect 31340 27560 31380 28880
rect 29980 27520 31380 27560
rect 34970 28880 36370 28920
rect 34970 27560 35010 28880
rect 36330 27560 36370 28880
rect 34970 27520 36370 27560
rect 39960 28880 41360 28920
rect 39960 27560 40000 28880
rect 41320 27560 41360 28880
rect 39960 27520 41360 27560
rect 44950 28880 46350 28920
rect 44950 27560 44990 28880
rect 46310 27560 46350 28880
rect 44950 27520 46350 27560
rect 49940 28880 51340 28920
rect 49940 27560 49980 28880
rect 51300 27560 51340 28880
rect 49940 27520 51340 27560
rect 54930 28880 56330 28920
rect 54930 27560 54970 28880
rect 56290 27560 56330 28880
rect 54930 27520 56330 27560
rect 59920 28880 61320 28920
rect 59920 27560 59960 28880
rect 61280 27560 61320 28880
rect 59920 27520 61320 27560
rect 64910 28880 66310 28920
rect 64910 27560 64950 28880
rect 66270 27560 66310 28880
rect 64910 27520 66310 27560
rect 69900 28880 71300 28920
rect 69900 27560 69940 28880
rect 71260 27560 71300 28880
rect 69900 27520 71300 27560
rect 74890 28880 76290 28920
rect 74890 27560 74930 28880
rect 76250 27560 76290 28880
rect 74890 27520 76290 27560
rect 79610 28880 81010 28920
rect 79610 27560 79650 28880
rect 80970 27560 81010 28880
rect 79610 27520 81010 27560
rect 79610 27170 81010 27210
rect 79610 25850 79650 27170
rect 80970 25850 81010 27170
rect 79610 25810 81010 25850
rect 79610 25460 81010 25500
rect 79610 24140 79650 25460
rect 80970 24140 81010 25460
rect 79610 24100 81010 24140
rect -4680 23750 -3280 23790
rect -4680 22430 -4640 23750
rect -3320 22430 -3280 23750
rect -4680 22390 -3280 22430
rect 79610 23750 81010 23790
rect 79610 22430 79650 23750
rect 80970 22430 81010 23750
rect 79610 22390 81010 22430
rect -4680 22040 -3280 22080
rect -4680 20720 -4640 22040
rect -3320 20720 -3280 22040
rect -4680 20680 -3280 20720
rect 79610 22040 81010 22080
rect 79610 20720 79650 22040
rect 80970 20720 81010 22040
rect 79610 20680 81010 20720
rect -4680 20330 -3280 20370
rect -4680 19010 -4640 20330
rect -3320 19010 -3280 20330
rect -4680 18970 -3280 19010
rect 79610 20330 81010 20370
rect 79610 19010 79650 20330
rect 80970 19010 81010 20330
rect 79610 18970 81010 19010
rect -4680 18620 -3280 18660
rect -4680 17300 -4640 18620
rect -3320 17300 -3280 18620
rect -4680 17260 -3280 17300
rect 79610 18620 81010 18660
rect 79610 17300 79650 18620
rect 80970 17300 81010 18620
rect 79610 17260 81010 17300
rect -4680 16910 -3280 16950
rect -4680 15590 -4640 16910
rect -3320 15590 -3280 16910
rect -4680 15550 -3280 15590
rect 79610 16910 81010 16950
rect 79610 15590 79650 16910
rect 80970 15590 81010 16910
rect 79610 15550 81010 15590
rect -4680 15200 -3280 15240
rect -4680 13880 -4640 15200
rect -3320 13880 -3280 15200
rect -4680 13840 -3280 13880
rect 79610 15200 81010 15240
rect 79610 13880 79650 15200
rect 80970 13880 81010 15200
rect 79610 13840 81010 13880
rect -4680 13490 -3280 13530
rect -4680 12170 -4640 13490
rect -3320 12170 -3280 13490
rect -4680 12130 -3280 12170
rect 79610 13490 81010 13530
rect 79610 12170 79650 13490
rect 80970 12170 81010 13490
rect 79610 12130 81010 12170
rect -4680 11780 -3280 11820
rect -4680 10460 -4640 11780
rect -3320 10460 -3280 11780
rect -4680 10420 -3280 10460
rect 79610 11780 81010 11820
rect 79610 10460 79650 11780
rect 80970 10460 81010 11780
rect 79610 10420 81010 10460
rect -4680 10070 -3280 10110
rect -4680 8750 -4640 10070
rect -3320 8750 -3280 10070
rect -4680 8710 -3280 8750
rect 79610 10070 81010 10110
rect 79610 8750 79650 10070
rect 80970 8750 81010 10070
rect 79610 8710 81010 8750
rect -4680 8360 -3280 8400
rect -4680 7040 -4640 8360
rect -3320 7040 -3280 8360
rect -4680 7000 -3280 7040
rect 79610 8360 81010 8400
rect 79610 7040 79650 8360
rect 80970 7040 81010 8360
rect 79610 7000 81010 7040
rect -4680 6650 -3280 6690
rect -4680 5330 -4640 6650
rect -3320 5330 -3280 6650
rect -4680 5290 -3280 5330
rect 79610 6650 81010 6690
rect 79610 5330 79650 6650
rect 80970 5330 81010 6650
rect 79610 5290 81010 5330
rect -4680 4940 -3280 4980
rect -4680 3620 -4640 4940
rect -3320 3620 -3280 4940
rect -4680 3580 -3280 3620
rect 79610 4940 81010 4980
rect 79610 3620 79650 4940
rect 80970 3620 81010 4940
rect 79610 3580 81010 3620
rect -4680 3230 -3280 3270
rect -4680 1910 -4640 3230
rect -3320 1910 -3280 3230
rect -4680 1870 -3280 1910
rect 79610 3230 81010 3270
rect 79610 1910 79650 3230
rect 80970 1910 81010 3230
rect 79610 1870 81010 1910
rect -4680 1520 -3280 1560
rect -4680 200 -4640 1520
rect -3320 200 -3280 1520
rect -4680 160 -3280 200
rect 79610 1520 81010 1560
rect 79610 200 79650 1520
rect 80970 200 81010 1520
rect 79610 160 81010 200
rect -4680 -190 -3280 -150
rect -4680 -1510 -4640 -190
rect -3320 -1510 -3280 -190
rect -4680 -1550 -3280 -1510
rect 40 -190 1440 -150
rect 40 -1510 80 -190
rect 1400 -1510 1440 -190
rect 40 -1550 1440 -1510
rect 5030 -190 6430 -150
rect 5030 -1510 5070 -190
rect 6390 -1510 6430 -190
rect 5030 -1550 6430 -1510
rect 10020 -190 11420 -150
rect 10020 -1510 10060 -190
rect 11380 -1510 11420 -190
rect 10020 -1550 11420 -1510
rect 15010 -190 16410 -150
rect 15010 -1510 15050 -190
rect 16370 -1510 16410 -190
rect 15010 -1550 16410 -1510
rect 20000 -190 21400 -150
rect 20000 -1510 20040 -190
rect 21360 -1510 21400 -190
rect 20000 -1550 21400 -1510
rect 24990 -190 26390 -150
rect 24990 -1510 25030 -190
rect 26350 -1510 26390 -190
rect 24990 -1550 26390 -1510
rect 29980 -190 31380 -150
rect 29980 -1510 30020 -190
rect 31340 -1510 31380 -190
rect 29980 -1550 31380 -1510
rect 34970 -190 36370 -150
rect 34970 -1510 35010 -190
rect 36330 -1510 36370 -190
rect 34970 -1550 36370 -1510
rect 39960 -190 41360 -150
rect 39960 -1510 40000 -190
rect 41320 -1510 41360 -190
rect 39960 -1550 41360 -1510
rect 44950 -190 46350 -150
rect 44950 -1510 44990 -190
rect 46310 -1510 46350 -190
rect 44950 -1550 46350 -1510
rect 49940 -190 51340 -150
rect 49940 -1510 49980 -190
rect 51300 -1510 51340 -190
rect 49940 -1550 51340 -1510
rect 54930 -190 56330 -150
rect 54930 -1510 54970 -190
rect 56290 -1510 56330 -190
rect 54930 -1550 56330 -1510
rect 59920 -190 61320 -150
rect 59920 -1510 59960 -190
rect 61280 -1510 61320 -190
rect 59920 -1550 61320 -1510
rect 64910 -190 66310 -150
rect 64910 -1510 64950 -190
rect 66270 -1510 66310 -190
rect 64910 -1550 66310 -1510
rect 69900 -190 71300 -150
rect 69900 -1510 69940 -190
rect 71260 -1510 71300 -190
rect 69900 -1550 71300 -1510
rect 74890 -190 76290 -150
rect 74890 -1510 74930 -190
rect 76250 -1510 76290 -190
rect 74890 -1550 76290 -1510
rect 79610 -190 81010 -150
rect 79610 -1510 79650 -190
rect 80970 -1510 81010 -190
rect 79610 -1550 81010 -1510
<< mimcapcontact >>
rect 80 27560 1400 28880
rect 5070 27560 6390 28880
rect 10060 27560 11380 28880
rect 15050 27560 16370 28880
rect 20040 27560 21360 28880
rect 25030 27560 26350 28880
rect 30020 27560 31340 28880
rect 35010 27560 36330 28880
rect 40000 27560 41320 28880
rect 44990 27560 46310 28880
rect 49980 27560 51300 28880
rect 54970 27560 56290 28880
rect 59960 27560 61280 28880
rect 64950 27560 66270 28880
rect 69940 27560 71260 28880
rect 74930 27560 76250 28880
rect 79650 27560 80970 28880
rect 79650 25850 80970 27170
rect 79650 24140 80970 25460
rect -4640 22430 -3320 23750
rect 79650 22430 80970 23750
rect -4640 20720 -3320 22040
rect 79650 20720 80970 22040
rect -4640 19010 -3320 20330
rect 79650 19010 80970 20330
rect -4640 17300 -3320 18620
rect 79650 17300 80970 18620
rect -4640 15590 -3320 16910
rect 79650 15590 80970 16910
rect -4640 13880 -3320 15200
rect 79650 13880 80970 15200
rect -4640 12170 -3320 13490
rect 79650 12170 80970 13490
rect -4640 10460 -3320 11780
rect 79650 10460 80970 11780
rect -4640 8750 -3320 10070
rect 79650 8750 80970 10070
rect -4640 7040 -3320 8360
rect 79650 7040 80970 8360
rect -4640 5330 -3320 6650
rect 79650 5330 80970 6650
rect -4640 3620 -3320 4940
rect 79650 3620 80970 4940
rect -4640 1910 -3320 3230
rect 79650 1910 80970 3230
rect -4640 200 -3320 1520
rect 79650 200 80970 1520
rect -4640 -1510 -3320 -190
rect 80 -1510 1400 -190
rect 5070 -1510 6390 -190
rect 10060 -1510 11380 -190
rect 15050 -1510 16370 -190
rect 20040 -1510 21360 -190
rect 25030 -1510 26350 -190
rect 30020 -1510 31340 -190
rect 35010 -1510 36330 -190
rect 40000 -1510 41320 -190
rect 44990 -1510 46310 -190
rect 49980 -1510 51300 -190
rect 54970 -1510 56290 -190
rect 59960 -1510 61280 -190
rect 64950 -1510 66270 -190
rect 69940 -1510 71260 -190
rect 74930 -1510 76250 -190
rect 79650 -1510 80970 -190
<< metal4 >>
rect -5530 30130 -5430 30140
rect -5530 30050 -5520 30130
rect -5440 30050 -5430 30130
rect -6370 29990 -5430 30050
rect -6370 29900 -6300 29990
rect -5690 29550 -5590 29610
rect 1672 28932 1768 28948
rect 79 28880 1401 28881
rect 1672 28880 1688 28932
rect 79 27560 80 28880
rect 1400 28820 1688 28880
rect 1400 27560 1401 28820
rect 79 27559 1401 27560
rect 1672 27508 1688 28820
rect 1752 28250 1768 28932
rect 6662 28932 6758 28948
rect 5069 28880 6391 28881
rect 6662 28880 6678 28932
rect 3140 28310 3280 28350
rect 3140 28250 3170 28310
rect 1752 28240 3170 28250
rect 3250 28240 3280 28310
rect 1752 28200 3280 28240
rect 1752 28190 3170 28200
rect 1752 27508 1768 28190
rect 3140 28130 3170 28190
rect 3250 28130 3280 28200
rect 3140 28100 3280 28130
rect 5069 27560 5070 28880
rect 6390 28820 6678 28880
rect 6390 27560 6391 28820
rect 5069 27559 6391 27560
rect 1672 27492 1768 27508
rect 6662 27508 6678 28820
rect 6742 28250 6758 28932
rect 11652 28932 11748 28948
rect 10059 28880 11381 28881
rect 11652 28880 11668 28932
rect 8130 28310 8270 28350
rect 8130 28250 8160 28310
rect 6742 28240 8160 28250
rect 8240 28240 8270 28310
rect 6742 28200 8270 28240
rect 6742 28190 8160 28200
rect 6742 27508 6758 28190
rect 8130 28130 8160 28190
rect 8240 28130 8270 28200
rect 8130 28100 8270 28130
rect 10059 27560 10060 28880
rect 11380 28820 11668 28880
rect 11380 27560 11381 28820
rect 10059 27559 11381 27560
rect 6662 27492 6758 27508
rect 11652 27508 11668 28820
rect 11732 28250 11748 28932
rect 16642 28932 16738 28948
rect 15049 28880 16371 28881
rect 16642 28880 16658 28932
rect 13120 28310 13260 28350
rect 13120 28250 13150 28310
rect 11732 28240 13150 28250
rect 13230 28240 13260 28310
rect 11732 28200 13260 28240
rect 11732 28190 13150 28200
rect 11732 27508 11748 28190
rect 13120 28130 13150 28190
rect 13230 28130 13260 28200
rect 13120 28100 13260 28130
rect 15049 27560 15050 28880
rect 16370 28820 16658 28880
rect 16370 27560 16371 28820
rect 15049 27559 16371 27560
rect 11652 27492 11748 27508
rect 16642 27508 16658 28820
rect 16722 28250 16738 28932
rect 21632 28932 21728 28948
rect 20039 28880 21361 28881
rect 21632 28880 21648 28932
rect 18110 28310 18250 28350
rect 18110 28250 18140 28310
rect 16722 28240 18140 28250
rect 18220 28240 18250 28310
rect 16722 28200 18250 28240
rect 16722 28190 18140 28200
rect 16722 27508 16738 28190
rect 18110 28130 18140 28190
rect 18220 28130 18250 28200
rect 18110 28100 18250 28130
rect 20039 27560 20040 28880
rect 21360 28820 21648 28880
rect 21360 27560 21361 28820
rect 20039 27559 21361 27560
rect 16642 27492 16738 27508
rect 21632 27508 21648 28820
rect 21712 28250 21728 28932
rect 26622 28932 26718 28948
rect 25029 28880 26351 28881
rect 26622 28880 26638 28932
rect 23100 28310 23240 28350
rect 23100 28250 23130 28310
rect 21712 28240 23130 28250
rect 23210 28240 23240 28310
rect 21712 28200 23240 28240
rect 21712 28190 23130 28200
rect 21712 27508 21728 28190
rect 23100 28130 23130 28190
rect 23210 28130 23240 28200
rect 23100 28100 23240 28130
rect 25029 27560 25030 28880
rect 26350 28820 26638 28880
rect 26350 27560 26351 28820
rect 25029 27559 26351 27560
rect 21632 27492 21728 27508
rect 26622 27508 26638 28820
rect 26702 28250 26718 28932
rect 31612 28932 31708 28948
rect 30019 28880 31341 28881
rect 31612 28880 31628 28932
rect 28090 28310 28230 28350
rect 28090 28250 28120 28310
rect 26702 28240 28120 28250
rect 28200 28240 28230 28310
rect 26702 28200 28230 28240
rect 26702 28190 28120 28200
rect 26702 27508 26718 28190
rect 28090 28130 28120 28190
rect 28200 28130 28230 28200
rect 28090 28100 28230 28130
rect 30019 27560 30020 28880
rect 31340 28820 31628 28880
rect 31340 27560 31341 28820
rect 30019 27559 31341 27560
rect 26622 27492 26718 27508
rect 31612 27508 31628 28820
rect 31692 28250 31708 28932
rect 36602 28932 36698 28948
rect 35009 28880 36331 28881
rect 36602 28880 36618 28932
rect 33080 28310 33220 28350
rect 33080 28250 33110 28310
rect 31692 28240 33110 28250
rect 33190 28240 33220 28310
rect 31692 28200 33220 28240
rect 31692 28190 33110 28200
rect 31692 27508 31708 28190
rect 33080 28130 33110 28190
rect 33190 28130 33220 28200
rect 33080 28100 33220 28130
rect 35009 27560 35010 28880
rect 36330 28820 36618 28880
rect 36330 27560 36331 28820
rect 35009 27559 36331 27560
rect 31612 27492 31708 27508
rect 36602 27508 36618 28820
rect 36682 28250 36698 28932
rect 41592 28932 41688 28948
rect 39999 28880 41321 28881
rect 41592 28880 41608 28932
rect 38070 28310 38210 28350
rect 38070 28250 38100 28310
rect 36682 28240 38100 28250
rect 38180 28240 38210 28310
rect 36682 28200 38210 28240
rect 36682 28190 38100 28200
rect 36682 27508 36698 28190
rect 38070 28130 38100 28190
rect 38180 28130 38210 28200
rect 38070 28100 38210 28130
rect 39999 27560 40000 28880
rect 41320 28820 41608 28880
rect 41320 27560 41321 28820
rect 39999 27559 41321 27560
rect 36602 27492 36698 27508
rect 41592 27508 41608 28820
rect 41672 28250 41688 28932
rect 46582 28932 46678 28948
rect 44989 28880 46311 28881
rect 46582 28880 46598 28932
rect 43060 28310 43200 28350
rect 43060 28250 43090 28310
rect 41672 28240 43090 28250
rect 43170 28240 43200 28310
rect 41672 28200 43200 28240
rect 41672 28190 43090 28200
rect 41672 27508 41688 28190
rect 43060 28130 43090 28190
rect 43170 28130 43200 28200
rect 43060 28100 43200 28130
rect 44989 27560 44990 28880
rect 46310 28820 46598 28880
rect 46310 27560 46311 28820
rect 44989 27559 46311 27560
rect 41592 27492 41688 27508
rect 46582 27508 46598 28820
rect 46662 28250 46678 28932
rect 51572 28932 51668 28948
rect 49979 28880 51301 28881
rect 51572 28880 51588 28932
rect 48050 28310 48190 28350
rect 48050 28250 48080 28310
rect 46662 28240 48080 28250
rect 48160 28240 48190 28310
rect 46662 28200 48190 28240
rect 46662 28190 48080 28200
rect 46662 27508 46678 28190
rect 48050 28130 48080 28190
rect 48160 28130 48190 28200
rect 48050 28100 48190 28130
rect 49979 27560 49980 28880
rect 51300 28820 51588 28880
rect 51300 27560 51301 28820
rect 49979 27559 51301 27560
rect 46582 27492 46678 27508
rect 51572 27508 51588 28820
rect 51652 28250 51668 28932
rect 56562 28932 56658 28948
rect 54969 28880 56291 28881
rect 56562 28880 56578 28932
rect 53040 28310 53180 28350
rect 53040 28250 53070 28310
rect 51652 28240 53070 28250
rect 53150 28240 53180 28310
rect 51652 28200 53180 28240
rect 51652 28190 53070 28200
rect 51652 27508 51668 28190
rect 53040 28130 53070 28190
rect 53150 28130 53180 28200
rect 53040 28100 53180 28130
rect 54969 27560 54970 28880
rect 56290 28820 56578 28880
rect 56290 27560 56291 28820
rect 54969 27559 56291 27560
rect 51572 27492 51668 27508
rect 56562 27508 56578 28820
rect 56642 28250 56658 28932
rect 61552 28932 61648 28948
rect 59959 28880 61281 28881
rect 61552 28880 61568 28932
rect 58030 28310 58170 28350
rect 58030 28250 58060 28310
rect 56642 28240 58060 28250
rect 58140 28240 58170 28310
rect 56642 28200 58170 28240
rect 56642 28190 58060 28200
rect 56642 27508 56658 28190
rect 58030 28130 58060 28190
rect 58140 28130 58170 28200
rect 58030 28100 58170 28130
rect 59959 27560 59960 28880
rect 61280 28820 61568 28880
rect 61280 27560 61281 28820
rect 59959 27559 61281 27560
rect 56562 27492 56658 27508
rect 61552 27508 61568 28820
rect 61632 28250 61648 28932
rect 66542 28932 66638 28948
rect 64949 28880 66271 28881
rect 66542 28880 66558 28932
rect 63020 28310 63160 28350
rect 63020 28250 63050 28310
rect 61632 28240 63050 28250
rect 63130 28240 63160 28310
rect 61632 28200 63160 28240
rect 61632 28190 63050 28200
rect 61632 27508 61648 28190
rect 63020 28130 63050 28190
rect 63130 28130 63160 28200
rect 63020 28100 63160 28130
rect 64949 27560 64950 28880
rect 66270 28820 66558 28880
rect 66270 27560 66271 28820
rect 64949 27559 66271 27560
rect 61552 27492 61648 27508
rect 66542 27508 66558 28820
rect 66622 28250 66638 28932
rect 71532 28932 71628 28948
rect 69939 28880 71261 28881
rect 71532 28880 71548 28932
rect 68010 28310 68150 28350
rect 68010 28250 68040 28310
rect 66622 28240 68040 28250
rect 68120 28240 68150 28310
rect 66622 28200 68150 28240
rect 66622 28190 68040 28200
rect 66622 27508 66638 28190
rect 68010 28130 68040 28190
rect 68120 28130 68150 28200
rect 68010 28100 68150 28130
rect 69939 27560 69940 28880
rect 71260 28820 71548 28880
rect 71260 27560 71261 28820
rect 69939 27559 71261 27560
rect 66542 27492 66638 27508
rect 71532 27508 71548 28820
rect 71612 28250 71628 28932
rect 76522 28932 76618 28948
rect 74929 28880 76251 28881
rect 76522 28880 76538 28932
rect 73000 28310 73140 28350
rect 73000 28250 73030 28310
rect 71612 28240 73030 28250
rect 73110 28240 73140 28310
rect 71612 28200 73140 28240
rect 71612 28190 73030 28200
rect 71612 27508 71628 28190
rect 73000 28130 73030 28190
rect 73110 28130 73140 28200
rect 73000 28100 73140 28130
rect 74929 27560 74930 28880
rect 76250 28820 76538 28880
rect 76250 27560 76251 28820
rect 74929 27559 76251 27560
rect 71532 27492 71628 27508
rect 76522 27508 76538 28820
rect 76602 28250 76618 28932
rect 81242 28932 81338 28948
rect 79649 28880 80971 28881
rect 81242 28880 81258 28932
rect 77990 28310 78130 28350
rect 77990 28250 78020 28310
rect 76602 28240 78020 28250
rect 78100 28240 78130 28310
rect 76602 28200 78130 28240
rect 76602 28190 78020 28200
rect 76602 27508 76618 28190
rect 77990 28130 78020 28190
rect 78100 28130 78130 28200
rect 77990 28100 78130 28130
rect 79649 27560 79650 28880
rect 80970 28820 81258 28880
rect 80970 27560 80971 28820
rect 79649 27559 80971 27560
rect 76522 27492 76618 27508
rect 81242 27508 81258 28820
rect 81322 28250 81338 28932
rect 82710 28310 82850 28350
rect 82710 28250 82740 28310
rect 81322 28240 82740 28250
rect 82820 28240 82850 28310
rect 81322 28200 82850 28240
rect 81322 28190 82740 28200
rect 81322 27508 81338 28190
rect 82710 28130 82740 28190
rect 82820 28130 82850 28200
rect 82710 28100 82850 28130
rect 81242 27492 81338 27508
rect 81242 27222 81338 27238
rect 79649 27170 80971 27171
rect 81242 27170 81258 27222
rect 79649 25850 79650 27170
rect 80970 27110 81258 27170
rect 80970 25850 80971 27110
rect 79649 25849 80971 25850
rect 81242 25798 81258 27110
rect 81322 26540 81338 27222
rect 82710 26600 82850 26640
rect 82710 26540 82740 26600
rect 81322 26530 82740 26540
rect 82820 26530 82850 26600
rect 81322 26490 82850 26530
rect 81322 26480 82740 26490
rect 81322 25798 81338 26480
rect 82710 26420 82740 26480
rect 82820 26420 82850 26490
rect 82710 26390 82850 26420
rect 81242 25782 81338 25798
rect 81242 25512 81338 25528
rect 79649 25460 80971 25461
rect 81242 25460 81258 25512
rect 79649 24140 79650 25460
rect 80970 25400 81258 25460
rect 80970 24140 80971 25400
rect 79649 24139 80971 24140
rect 81242 24088 81258 25400
rect 81322 24830 81338 25512
rect 82710 24890 82850 24930
rect 82710 24830 82740 24890
rect 81322 24820 82740 24830
rect 82820 24820 82850 24890
rect 81322 24780 82850 24820
rect 81322 24770 82740 24780
rect 81322 24088 81338 24770
rect 82710 24710 82740 24770
rect 82820 24710 82850 24780
rect 82710 24680 82850 24710
rect 81242 24072 81338 24088
rect -3048 23802 -2952 23818
rect -4641 23750 -3319 23751
rect -3048 23750 -3032 23802
rect -4641 22430 -4640 23750
rect -3320 23690 -3032 23750
rect -3320 22430 -3319 23690
rect -4641 22429 -3319 22430
rect -3048 22378 -3032 23690
rect -2968 23120 -2952 23802
rect 81242 23802 81338 23818
rect 79649 23750 80971 23751
rect 81242 23750 81258 23802
rect -1580 23180 -1440 23220
rect -1580 23120 -1550 23180
rect -2968 23110 -1550 23120
rect -1470 23110 -1440 23180
rect -2968 23070 -1440 23110
rect -2968 23060 -1550 23070
rect -2968 22378 -2952 23060
rect -1580 23000 -1550 23060
rect -1470 23000 -1440 23070
rect -1580 22970 -1440 23000
rect 79649 22430 79650 23750
rect 80970 23690 81258 23750
rect 80970 22430 80971 23690
rect 79649 22429 80971 22430
rect -3048 22362 -2952 22378
rect 81242 22378 81258 23690
rect 81322 23120 81338 23802
rect 82710 23180 82850 23220
rect 82710 23120 82740 23180
rect 81322 23110 82740 23120
rect 82820 23110 82850 23180
rect 81322 23070 82850 23110
rect 81322 23060 82740 23070
rect 81322 22378 81338 23060
rect 82710 23000 82740 23060
rect 82820 23000 82850 23070
rect 82710 22970 82850 23000
rect 81242 22362 81338 22378
rect -3048 22092 -2952 22108
rect -4641 22040 -3319 22041
rect -3048 22040 -3032 22092
rect -4641 20720 -4640 22040
rect -3320 21980 -3032 22040
rect -3320 20720 -3319 21980
rect -4641 20719 -3319 20720
rect -3048 20668 -3032 21980
rect -2968 21410 -2952 22092
rect 81242 22092 81338 22108
rect 79649 22040 80971 22041
rect 81242 22040 81258 22092
rect -1580 21470 -1440 21510
rect -1580 21410 -1550 21470
rect -2968 21400 -1550 21410
rect -1470 21400 -1440 21470
rect -2968 21360 -1440 21400
rect -2968 21350 -1550 21360
rect -2968 20668 -2952 21350
rect -1580 21290 -1550 21350
rect -1470 21290 -1440 21360
rect -1580 21260 -1440 21290
rect 79649 20720 79650 22040
rect 80970 21980 81258 22040
rect 80970 20720 80971 21980
rect 79649 20719 80971 20720
rect -3048 20652 -2952 20668
rect 81242 20668 81258 21980
rect 81322 21410 81338 22092
rect 82710 21470 82850 21510
rect 82710 21410 82740 21470
rect 81322 21400 82740 21410
rect 82820 21400 82850 21470
rect 81322 21360 82850 21400
rect 81322 21350 82740 21360
rect 81322 20668 81338 21350
rect 82710 21290 82740 21350
rect 82820 21290 82850 21360
rect 82710 21260 82850 21290
rect 81242 20652 81338 20668
rect -3048 20382 -2952 20398
rect -4641 20330 -3319 20331
rect -3048 20330 -3032 20382
rect -4641 19010 -4640 20330
rect -3320 20270 -3032 20330
rect -3320 19010 -3319 20270
rect -4641 19009 -3319 19010
rect -3048 18958 -3032 20270
rect -2968 19700 -2952 20382
rect 81242 20382 81338 20398
rect 79649 20330 80971 20331
rect 81242 20330 81258 20382
rect -1580 19760 -1440 19800
rect -1580 19700 -1550 19760
rect -2968 19690 -1550 19700
rect -1470 19690 -1440 19760
rect -2968 19650 -1440 19690
rect -2968 19640 -1550 19650
rect -2968 18958 -2952 19640
rect -1580 19580 -1550 19640
rect -1470 19580 -1440 19650
rect -1580 19550 -1440 19580
rect 79649 19010 79650 20330
rect 80970 20270 81258 20330
rect 80970 19010 80971 20270
rect 79649 19009 80971 19010
rect -3048 18942 -2952 18958
rect 81242 18958 81258 20270
rect 81322 19700 81338 20382
rect 82710 19760 82850 19800
rect 82710 19700 82740 19760
rect 81322 19690 82740 19700
rect 82820 19690 82850 19760
rect 81322 19650 82850 19690
rect 81322 19640 82740 19650
rect 81322 18958 81338 19640
rect 82710 19580 82740 19640
rect 82820 19580 82850 19650
rect 82710 19550 82850 19580
rect 81242 18942 81338 18958
rect -3048 18672 -2952 18688
rect -4641 18620 -3319 18621
rect -3048 18620 -3032 18672
rect -4641 17300 -4640 18620
rect -3320 18560 -3032 18620
rect -3320 17300 -3319 18560
rect -4641 17299 -3319 17300
rect -3048 17248 -3032 18560
rect -2968 17990 -2952 18672
rect 81242 18672 81338 18688
rect 79649 18620 80971 18621
rect 81242 18620 81258 18672
rect -1580 18050 -1440 18090
rect -1580 17990 -1550 18050
rect -2968 17980 -1550 17990
rect -1470 17980 -1440 18050
rect -2968 17940 -1440 17980
rect -2968 17930 -1550 17940
rect -2968 17248 -2952 17930
rect -1580 17870 -1550 17930
rect -1470 17870 -1440 17940
rect -1580 17840 -1440 17870
rect 79649 17300 79650 18620
rect 80970 18560 81258 18620
rect 80970 17300 80971 18560
rect 79649 17299 80971 17300
rect -3048 17232 -2952 17248
rect 81242 17248 81258 18560
rect 81322 17990 81338 18672
rect 82710 18050 82850 18090
rect 82710 17990 82740 18050
rect 81322 17980 82740 17990
rect 82820 17980 82850 18050
rect 81322 17940 82850 17980
rect 81322 17930 82740 17940
rect 81322 17248 81338 17930
rect 82710 17870 82740 17930
rect 82820 17870 82850 17940
rect 82710 17840 82850 17870
rect 81242 17232 81338 17248
rect -3048 16962 -2952 16978
rect -4641 16910 -3319 16911
rect -3048 16910 -3032 16962
rect -4641 15590 -4640 16910
rect -3320 16850 -3032 16910
rect -3320 15590 -3319 16850
rect -4641 15589 -3319 15590
rect -3048 15538 -3032 16850
rect -2968 16280 -2952 16962
rect 81242 16962 81338 16978
rect 79649 16910 80971 16911
rect 81242 16910 81258 16962
rect -1580 16340 -1440 16380
rect -1580 16280 -1550 16340
rect -2968 16270 -1550 16280
rect -1470 16270 -1440 16340
rect -2968 16230 -1440 16270
rect -2968 16220 -1550 16230
rect -2968 15538 -2952 16220
rect -1580 16160 -1550 16220
rect -1470 16160 -1440 16230
rect -1580 16130 -1440 16160
rect 79649 15590 79650 16910
rect 80970 16850 81258 16910
rect 80970 15590 80971 16850
rect 79649 15589 80971 15590
rect -3048 15522 -2952 15538
rect 81242 15538 81258 16850
rect 81322 16280 81338 16962
rect 82710 16340 82850 16380
rect 82710 16280 82740 16340
rect 81322 16270 82740 16280
rect 82820 16270 82850 16340
rect 81322 16230 82850 16270
rect 81322 16220 82740 16230
rect 81322 15538 81338 16220
rect 82710 16160 82740 16220
rect 82820 16160 82850 16230
rect 82710 16130 82850 16160
rect 81242 15522 81338 15538
rect -3048 15252 -2952 15268
rect -4641 15200 -3319 15201
rect -3048 15200 -3032 15252
rect -4641 13880 -4640 15200
rect -3320 15140 -3032 15200
rect -3320 13880 -3319 15140
rect -4641 13879 -3319 13880
rect -3048 13828 -3032 15140
rect -2968 14570 -2952 15252
rect 81242 15252 81338 15268
rect 79649 15200 80971 15201
rect 81242 15200 81258 15252
rect -1580 14630 -1440 14670
rect -1580 14570 -1550 14630
rect -2968 14560 -1550 14570
rect -1470 14560 -1440 14630
rect -2968 14520 -1440 14560
rect -2968 14510 -1550 14520
rect -2968 13828 -2952 14510
rect -1580 14450 -1550 14510
rect -1470 14450 -1440 14520
rect -1580 14420 -1440 14450
rect 79649 13880 79650 15200
rect 80970 15140 81258 15200
rect 80970 13880 80971 15140
rect 79649 13879 80971 13880
rect -3048 13812 -2952 13828
rect 81242 13828 81258 15140
rect 81322 14570 81338 15252
rect 82710 14630 82850 14670
rect 82710 14570 82740 14630
rect 81322 14560 82740 14570
rect 82820 14560 82850 14630
rect 81322 14520 82850 14560
rect 81322 14510 82740 14520
rect 81322 13828 81338 14510
rect 82710 14450 82740 14510
rect 82820 14450 82850 14520
rect 82710 14420 82850 14450
rect 81242 13812 81338 13828
rect -3048 13542 -2952 13558
rect -4641 13490 -3319 13491
rect -3048 13490 -3032 13542
rect -4641 12170 -4640 13490
rect -3320 13430 -3032 13490
rect -3320 12170 -3319 13430
rect -4641 12169 -3319 12170
rect -3048 12118 -3032 13430
rect -2968 12860 -2952 13542
rect 81242 13542 81338 13558
rect 79649 13490 80971 13491
rect 81242 13490 81258 13542
rect -1580 12920 -1440 12960
rect -1580 12860 -1550 12920
rect -2968 12850 -1550 12860
rect -1470 12850 -1440 12920
rect -2968 12810 -1440 12850
rect -2968 12800 -1550 12810
rect -2968 12118 -2952 12800
rect -1580 12740 -1550 12800
rect -1470 12740 -1440 12810
rect -1580 12710 -1440 12740
rect 79649 12170 79650 13490
rect 80970 13430 81258 13490
rect 80970 12170 80971 13430
rect 79649 12169 80971 12170
rect -3048 12102 -2952 12118
rect 81242 12118 81258 13430
rect 81322 12860 81338 13542
rect 82710 12920 82850 12960
rect 82710 12860 82740 12920
rect 81322 12850 82740 12860
rect 82820 12850 82850 12920
rect 81322 12810 82850 12850
rect 81322 12800 82740 12810
rect 81322 12118 81338 12800
rect 82710 12740 82740 12800
rect 82820 12740 82850 12810
rect 82710 12710 82850 12740
rect 81242 12102 81338 12118
rect -3048 11832 -2952 11848
rect -4641 11780 -3319 11781
rect -3048 11780 -3032 11832
rect -4641 10460 -4640 11780
rect -3320 11720 -3032 11780
rect -3320 10460 -3319 11720
rect -4641 10459 -3319 10460
rect -3048 10408 -3032 11720
rect -2968 11150 -2952 11832
rect 81242 11832 81338 11848
rect 79649 11780 80971 11781
rect 81242 11780 81258 11832
rect -1580 11210 -1440 11250
rect -1580 11150 -1550 11210
rect -2968 11140 -1550 11150
rect -1470 11140 -1440 11210
rect -2968 11100 -1440 11140
rect -2968 11090 -1550 11100
rect -2968 10408 -2952 11090
rect -1580 11030 -1550 11090
rect -1470 11030 -1440 11100
rect -1580 11000 -1440 11030
rect 79649 10460 79650 11780
rect 80970 11720 81258 11780
rect 80970 10460 80971 11720
rect 79649 10459 80971 10460
rect -3048 10392 -2952 10408
rect 81242 10408 81258 11720
rect 81322 11150 81338 11832
rect 82710 11210 82850 11250
rect 82710 11150 82740 11210
rect 81322 11140 82740 11150
rect 82820 11140 82850 11210
rect 81322 11100 82850 11140
rect 81322 11090 82740 11100
rect 81322 10408 81338 11090
rect 82710 11030 82740 11090
rect 82820 11030 82850 11100
rect 82710 11000 82850 11030
rect 81242 10392 81338 10408
rect -3048 10122 -2952 10138
rect -4641 10070 -3319 10071
rect -3048 10070 -3032 10122
rect -4641 8750 -4640 10070
rect -3320 10010 -3032 10070
rect -3320 8750 -3319 10010
rect -4641 8749 -3319 8750
rect -3048 8698 -3032 10010
rect -2968 9440 -2952 10122
rect 81242 10122 81338 10138
rect 79649 10070 80971 10071
rect 81242 10070 81258 10122
rect -1580 9500 -1440 9540
rect -1580 9440 -1550 9500
rect -2968 9430 -1550 9440
rect -1470 9430 -1440 9500
rect -2968 9390 -1440 9430
rect -2968 9380 -1550 9390
rect -2968 8698 -2952 9380
rect -1580 9320 -1550 9380
rect -1470 9320 -1440 9390
rect -1580 9290 -1440 9320
rect 79649 8750 79650 10070
rect 80970 10010 81258 10070
rect 80970 8750 80971 10010
rect 79649 8749 80971 8750
rect -3048 8682 -2952 8698
rect 81242 8698 81258 10010
rect 81322 9440 81338 10122
rect 82710 9500 82850 9540
rect 82710 9440 82740 9500
rect 81322 9430 82740 9440
rect 82820 9430 82850 9500
rect 81322 9390 82850 9430
rect 81322 9380 82740 9390
rect 81322 8698 81338 9380
rect 82710 9320 82740 9380
rect 82820 9320 82850 9390
rect 82710 9290 82850 9320
rect 81242 8682 81338 8698
rect -3048 8412 -2952 8428
rect -4641 8360 -3319 8361
rect -3048 8360 -3032 8412
rect -4641 7040 -4640 8360
rect -3320 8300 -3032 8360
rect -3320 7040 -3319 8300
rect -4641 7039 -3319 7040
rect -3048 6988 -3032 8300
rect -2968 7730 -2952 8412
rect 81242 8412 81338 8428
rect 79649 8360 80971 8361
rect 81242 8360 81258 8412
rect -1580 7790 -1440 7830
rect -1580 7730 -1550 7790
rect -2968 7720 -1550 7730
rect -1470 7720 -1440 7790
rect -2968 7680 -1440 7720
rect -2968 7670 -1550 7680
rect -2968 6988 -2952 7670
rect -1580 7610 -1550 7670
rect -1470 7610 -1440 7680
rect -1580 7580 -1440 7610
rect 79649 7040 79650 8360
rect 80970 8300 81258 8360
rect 80970 7040 80971 8300
rect 79649 7039 80971 7040
rect -3048 6972 -2952 6988
rect 81242 6988 81258 8300
rect 81322 7730 81338 8412
rect 82710 7790 82850 7830
rect 82710 7730 82740 7790
rect 81322 7720 82740 7730
rect 82820 7720 82850 7790
rect 81322 7680 82850 7720
rect 81322 7670 82740 7680
rect 81322 6988 81338 7670
rect 82710 7610 82740 7670
rect 82820 7610 82850 7680
rect 82710 7580 82850 7610
rect 81242 6972 81338 6988
rect -3048 6702 -2952 6718
rect -4641 6650 -3319 6651
rect -3048 6650 -3032 6702
rect -4641 5330 -4640 6650
rect -3320 6590 -3032 6650
rect -3320 5330 -3319 6590
rect -4641 5329 -3319 5330
rect -3048 5278 -3032 6590
rect -2968 6020 -2952 6702
rect 81242 6702 81338 6718
rect 79649 6650 80971 6651
rect 81242 6650 81258 6702
rect -1580 6080 -1440 6120
rect -1580 6020 -1550 6080
rect -2968 6010 -1550 6020
rect -1470 6010 -1440 6080
rect -2968 5970 -1440 6010
rect -2968 5960 -1550 5970
rect -2968 5278 -2952 5960
rect -1580 5900 -1550 5960
rect -1470 5900 -1440 5970
rect -1580 5870 -1440 5900
rect 79649 5330 79650 6650
rect 80970 6590 81258 6650
rect 80970 5330 80971 6590
rect 79649 5329 80971 5330
rect -3048 5262 -2952 5278
rect 81242 5278 81258 6590
rect 81322 6020 81338 6702
rect 82710 6080 82850 6120
rect 82710 6020 82740 6080
rect 81322 6010 82740 6020
rect 82820 6010 82850 6080
rect 81322 5970 82850 6010
rect 81322 5960 82740 5970
rect 81322 5278 81338 5960
rect 82710 5900 82740 5960
rect 82820 5900 82850 5970
rect 82710 5870 82850 5900
rect 81242 5262 81338 5278
rect -3048 4992 -2952 5008
rect -4641 4940 -3319 4941
rect -3048 4940 -3032 4992
rect -4641 3620 -4640 4940
rect -3320 4880 -3032 4940
rect -3320 3620 -3319 4880
rect -4641 3619 -3319 3620
rect -3048 3568 -3032 4880
rect -2968 4310 -2952 4992
rect 81242 4992 81338 5008
rect 79649 4940 80971 4941
rect 81242 4940 81258 4992
rect -1580 4370 -1440 4410
rect -1580 4310 -1550 4370
rect -2968 4300 -1550 4310
rect -1470 4300 -1440 4370
rect -2968 4260 -1440 4300
rect -2968 4250 -1550 4260
rect -2968 3568 -2952 4250
rect -1580 4190 -1550 4250
rect -1470 4190 -1440 4260
rect -1580 4160 -1440 4190
rect 79649 3620 79650 4940
rect 80970 4880 81258 4940
rect 80970 3620 80971 4880
rect 79649 3619 80971 3620
rect -3048 3552 -2952 3568
rect 81242 3568 81258 4880
rect 81322 4310 81338 4992
rect 82710 4370 82850 4410
rect 82710 4310 82740 4370
rect 81322 4300 82740 4310
rect 82820 4300 82850 4370
rect 81322 4260 82850 4300
rect 81322 4250 82740 4260
rect 81322 3568 81338 4250
rect 82710 4190 82740 4250
rect 82820 4190 82850 4260
rect 82710 4160 82850 4190
rect 81242 3552 81338 3568
rect -3048 3282 -2952 3298
rect -4641 3230 -3319 3231
rect -3048 3230 -3032 3282
rect -4641 1910 -4640 3230
rect -3320 3170 -3032 3230
rect -3320 1910 -3319 3170
rect -4641 1909 -3319 1910
rect -3048 1858 -3032 3170
rect -2968 2600 -2952 3282
rect 81242 3282 81338 3298
rect 79649 3230 80971 3231
rect 81242 3230 81258 3282
rect -1580 2660 -1440 2700
rect -1580 2600 -1550 2660
rect -2968 2590 -1550 2600
rect -1470 2590 -1440 2660
rect -2968 2550 -1440 2590
rect -2968 2540 -1550 2550
rect -2968 1858 -2952 2540
rect -1580 2480 -1550 2540
rect -1470 2480 -1440 2550
rect -1580 2450 -1440 2480
rect 79649 1910 79650 3230
rect 80970 3170 81258 3230
rect 80970 1910 80971 3170
rect 79649 1909 80971 1910
rect -3048 1842 -2952 1858
rect 81242 1858 81258 3170
rect 81322 2600 81338 3282
rect 82710 2660 82850 2700
rect 82710 2600 82740 2660
rect 81322 2590 82740 2600
rect 82820 2590 82850 2660
rect 81322 2550 82850 2590
rect 81322 2540 82740 2550
rect 81322 1858 81338 2540
rect 82710 2480 82740 2540
rect 82820 2480 82850 2550
rect 82710 2450 82850 2480
rect 81242 1842 81338 1858
rect -3048 1572 -2952 1588
rect -4641 1520 -3319 1521
rect -3048 1520 -3032 1572
rect -4641 200 -4640 1520
rect -3320 1460 -3032 1520
rect -3320 200 -3319 1460
rect -4641 199 -3319 200
rect -3048 148 -3032 1460
rect -2968 890 -2952 1572
rect 81242 1572 81338 1588
rect 79649 1520 80971 1521
rect 81242 1520 81258 1572
rect -1580 950 -1440 990
rect -1580 890 -1550 950
rect -2968 880 -1550 890
rect -1470 880 -1440 950
rect -2968 840 -1440 880
rect -2968 830 -1550 840
rect -2968 148 -2952 830
rect -1580 770 -1550 830
rect -1470 770 -1440 840
rect -1580 740 -1440 770
rect 79649 200 79650 1520
rect 80970 1460 81258 1520
rect 80970 200 80971 1460
rect 79649 199 80971 200
rect -3048 132 -2952 148
rect 81242 148 81258 1460
rect 81322 890 81338 1572
rect 82710 950 82850 990
rect 82710 890 82740 950
rect 81322 880 82740 890
rect 82820 880 82850 950
rect 81322 840 82850 880
rect 81322 830 82740 840
rect 81322 148 81338 830
rect 82710 770 82740 830
rect 82820 770 82850 840
rect 82710 740 82850 770
rect 81242 132 81338 148
rect 80 40 140 100
rect 5070 40 5130 100
rect 10060 40 10120 100
rect 15050 40 15110 100
rect 20040 40 20100 100
rect 25030 40 25090 100
rect 30020 40 30080 100
rect 35010 40 35070 100
rect 40000 40 40060 100
rect 44990 40 45050 100
rect 49980 40 50040 100
rect 54970 40 55030 100
rect 59960 40 60020 100
rect 64950 40 65010 100
rect 69940 40 70000 100
rect 74930 40 74990 100
rect -4720 -20 78640 40
rect 78580 -70 78640 -20
rect 79510 -20 84330 40
rect 79510 -70 79570 -20
rect -3048 -138 -2952 -122
rect -4641 -190 -3319 -189
rect -3048 -190 -3032 -138
rect -4641 -1510 -4640 -190
rect -3320 -250 -3032 -190
rect -3320 -1510 -3319 -250
rect -4641 -1511 -3319 -1510
rect -3048 -1562 -3032 -250
rect -2968 -820 -2952 -138
rect 1672 -138 1768 -122
rect 79 -190 1401 -189
rect 1672 -190 1688 -138
rect -1580 -760 -1440 -720
rect -1580 -820 -1550 -760
rect -2968 -830 -1550 -820
rect -1470 -830 -1440 -760
rect -2968 -870 -1440 -830
rect -2968 -880 -1550 -870
rect -2968 -1562 -2952 -880
rect -1580 -940 -1550 -880
rect -1470 -940 -1440 -870
rect -1580 -970 -1440 -940
rect 79 -1510 80 -190
rect 1400 -250 1688 -190
rect 1400 -1510 1401 -250
rect 79 -1511 1401 -1510
rect -3048 -1578 -2952 -1562
rect 1672 -1562 1688 -250
rect 1752 -820 1768 -138
rect 6662 -138 6758 -122
rect 5069 -190 6391 -189
rect 6662 -190 6678 -138
rect 3140 -760 3280 -720
rect 3140 -820 3170 -760
rect 1752 -830 3170 -820
rect 3250 -830 3280 -760
rect 1752 -870 3280 -830
rect 1752 -880 3170 -870
rect 1752 -1562 1768 -880
rect 3140 -940 3170 -880
rect 3250 -940 3280 -870
rect 3140 -970 3280 -940
rect 5069 -1510 5070 -190
rect 6390 -250 6678 -190
rect 6390 -1510 6391 -250
rect 5069 -1511 6391 -1510
rect 1672 -1578 1768 -1562
rect 6662 -1562 6678 -250
rect 6742 -820 6758 -138
rect 11652 -138 11748 -122
rect 10059 -190 11381 -189
rect 11652 -190 11668 -138
rect 8130 -760 8270 -720
rect 8130 -820 8160 -760
rect 6742 -830 8160 -820
rect 8240 -830 8270 -760
rect 6742 -870 8270 -830
rect 6742 -880 8160 -870
rect 6742 -1562 6758 -880
rect 8130 -940 8160 -880
rect 8240 -940 8270 -870
rect 8130 -970 8270 -940
rect 10059 -1510 10060 -190
rect 11380 -250 11668 -190
rect 11380 -1510 11381 -250
rect 10059 -1511 11381 -1510
rect 6662 -1578 6758 -1562
rect 11652 -1562 11668 -250
rect 11732 -820 11748 -138
rect 16642 -138 16738 -122
rect 15049 -190 16371 -189
rect 16642 -190 16658 -138
rect 13120 -760 13260 -720
rect 13120 -820 13150 -760
rect 11732 -830 13150 -820
rect 13230 -830 13260 -760
rect 11732 -870 13260 -830
rect 11732 -880 13150 -870
rect 11732 -1562 11748 -880
rect 13120 -940 13150 -880
rect 13230 -940 13260 -870
rect 13120 -970 13260 -940
rect 15049 -1510 15050 -190
rect 16370 -250 16658 -190
rect 16370 -1510 16371 -250
rect 15049 -1511 16371 -1510
rect 11652 -1578 11748 -1562
rect 16642 -1562 16658 -250
rect 16722 -820 16738 -138
rect 21632 -138 21728 -122
rect 20039 -190 21361 -189
rect 21632 -190 21648 -138
rect 18110 -760 18250 -720
rect 18110 -820 18140 -760
rect 16722 -830 18140 -820
rect 18220 -830 18250 -760
rect 16722 -870 18250 -830
rect 16722 -880 18140 -870
rect 16722 -1562 16738 -880
rect 18110 -940 18140 -880
rect 18220 -940 18250 -870
rect 18110 -970 18250 -940
rect 20039 -1510 20040 -190
rect 21360 -250 21648 -190
rect 21360 -1510 21361 -250
rect 20039 -1511 21361 -1510
rect 16642 -1578 16738 -1562
rect 21632 -1562 21648 -250
rect 21712 -820 21728 -138
rect 26622 -138 26718 -122
rect 25029 -190 26351 -189
rect 26622 -190 26638 -138
rect 23100 -760 23240 -720
rect 23100 -820 23130 -760
rect 21712 -830 23130 -820
rect 23210 -830 23240 -760
rect 21712 -870 23240 -830
rect 21712 -880 23130 -870
rect 21712 -1562 21728 -880
rect 23100 -940 23130 -880
rect 23210 -940 23240 -870
rect 23100 -970 23240 -940
rect 25029 -1510 25030 -190
rect 26350 -250 26638 -190
rect 26350 -1510 26351 -250
rect 25029 -1511 26351 -1510
rect 21632 -1578 21728 -1562
rect 26622 -1562 26638 -250
rect 26702 -820 26718 -138
rect 31612 -138 31708 -122
rect 30019 -190 31341 -189
rect 31612 -190 31628 -138
rect 28090 -760 28230 -720
rect 28090 -820 28120 -760
rect 26702 -830 28120 -820
rect 28200 -830 28230 -760
rect 26702 -870 28230 -830
rect 26702 -880 28120 -870
rect 26702 -1562 26718 -880
rect 28090 -940 28120 -880
rect 28200 -940 28230 -870
rect 28090 -970 28230 -940
rect 30019 -1510 30020 -190
rect 31340 -250 31628 -190
rect 31340 -1510 31341 -250
rect 30019 -1511 31341 -1510
rect 26622 -1578 26718 -1562
rect 31612 -1562 31628 -250
rect 31692 -820 31708 -138
rect 36602 -138 36698 -122
rect 35009 -190 36331 -189
rect 36602 -190 36618 -138
rect 33080 -760 33220 -720
rect 33080 -820 33110 -760
rect 31692 -830 33110 -820
rect 33190 -830 33220 -760
rect 31692 -870 33220 -830
rect 31692 -880 33110 -870
rect 31692 -1562 31708 -880
rect 33080 -940 33110 -880
rect 33190 -940 33220 -870
rect 33080 -970 33220 -940
rect 35009 -1510 35010 -190
rect 36330 -250 36618 -190
rect 36330 -1510 36331 -250
rect 35009 -1511 36331 -1510
rect 31612 -1578 31708 -1562
rect 36602 -1562 36618 -250
rect 36682 -820 36698 -138
rect 41592 -138 41688 -122
rect 39999 -190 41321 -189
rect 41592 -190 41608 -138
rect 38070 -760 38210 -720
rect 38070 -820 38100 -760
rect 36682 -830 38100 -820
rect 38180 -830 38210 -760
rect 36682 -870 38210 -830
rect 36682 -880 38100 -870
rect 36682 -1562 36698 -880
rect 38070 -940 38100 -880
rect 38180 -940 38210 -870
rect 38070 -970 38210 -940
rect 39999 -1510 40000 -190
rect 41320 -250 41608 -190
rect 41320 -1510 41321 -250
rect 39999 -1511 41321 -1510
rect 36602 -1578 36698 -1562
rect 41592 -1562 41608 -250
rect 41672 -820 41688 -138
rect 46582 -138 46678 -122
rect 44989 -190 46311 -189
rect 46582 -190 46598 -138
rect 43060 -760 43200 -720
rect 43060 -820 43090 -760
rect 41672 -830 43090 -820
rect 43170 -830 43200 -760
rect 41672 -870 43200 -830
rect 41672 -880 43090 -870
rect 41672 -1562 41688 -880
rect 43060 -940 43090 -880
rect 43170 -940 43200 -870
rect 43060 -970 43200 -940
rect 44989 -1510 44990 -190
rect 46310 -250 46598 -190
rect 46310 -1510 46311 -250
rect 44989 -1511 46311 -1510
rect 41592 -1578 41688 -1562
rect 46582 -1562 46598 -250
rect 46662 -820 46678 -138
rect 51572 -138 51668 -122
rect 49979 -190 51301 -189
rect 51572 -190 51588 -138
rect 48050 -760 48190 -720
rect 48050 -820 48080 -760
rect 46662 -830 48080 -820
rect 48160 -830 48190 -760
rect 46662 -870 48190 -830
rect 46662 -880 48080 -870
rect 46662 -1562 46678 -880
rect 48050 -940 48080 -880
rect 48160 -940 48190 -870
rect 48050 -970 48190 -940
rect 49979 -1510 49980 -190
rect 51300 -250 51588 -190
rect 51300 -1510 51301 -250
rect 49979 -1511 51301 -1510
rect 46582 -1578 46678 -1562
rect 51572 -1562 51588 -250
rect 51652 -820 51668 -138
rect 56562 -138 56658 -122
rect 54969 -190 56291 -189
rect 56562 -190 56578 -138
rect 53040 -760 53180 -720
rect 53040 -820 53070 -760
rect 51652 -830 53070 -820
rect 53150 -830 53180 -760
rect 51652 -870 53180 -830
rect 51652 -880 53070 -870
rect 51652 -1562 51668 -880
rect 53040 -940 53070 -880
rect 53150 -940 53180 -870
rect 53040 -970 53180 -940
rect 54969 -1510 54970 -190
rect 56290 -250 56578 -190
rect 56290 -1510 56291 -250
rect 54969 -1511 56291 -1510
rect 51572 -1578 51668 -1562
rect 56562 -1562 56578 -250
rect 56642 -820 56658 -138
rect 61552 -138 61648 -122
rect 59959 -190 61281 -189
rect 61552 -190 61568 -138
rect 58030 -760 58170 -720
rect 58030 -820 58060 -760
rect 56642 -830 58060 -820
rect 58140 -830 58170 -760
rect 56642 -870 58170 -830
rect 56642 -880 58060 -870
rect 56642 -1562 56658 -880
rect 58030 -940 58060 -880
rect 58140 -940 58170 -870
rect 58030 -970 58170 -940
rect 59959 -1510 59960 -190
rect 61280 -250 61568 -190
rect 61280 -1510 61281 -250
rect 59959 -1511 61281 -1510
rect 56562 -1578 56658 -1562
rect 61552 -1562 61568 -250
rect 61632 -820 61648 -138
rect 66542 -138 66638 -122
rect 64949 -190 66271 -189
rect 66542 -190 66558 -138
rect 63020 -760 63160 -720
rect 63020 -820 63050 -760
rect 61632 -830 63050 -820
rect 63130 -830 63160 -760
rect 61632 -870 63160 -830
rect 61632 -880 63050 -870
rect 61632 -1562 61648 -880
rect 63020 -940 63050 -880
rect 63130 -940 63160 -870
rect 63020 -970 63160 -940
rect 64949 -1510 64950 -190
rect 66270 -250 66558 -190
rect 66270 -1510 66271 -250
rect 64949 -1511 66271 -1510
rect 61552 -1578 61648 -1562
rect 66542 -1562 66558 -250
rect 66622 -820 66638 -138
rect 71532 -138 71628 -122
rect 69939 -190 71261 -189
rect 71532 -190 71548 -138
rect 68010 -760 68150 -720
rect 68010 -820 68040 -760
rect 66622 -830 68040 -820
rect 68120 -830 68150 -760
rect 66622 -870 68150 -830
rect 66622 -880 68040 -870
rect 66622 -1562 66638 -880
rect 68010 -940 68040 -880
rect 68120 -940 68150 -870
rect 68010 -970 68150 -940
rect 69939 -1510 69940 -190
rect 71260 -250 71548 -190
rect 71260 -1510 71261 -250
rect 69939 -1511 71261 -1510
rect 66542 -1578 66638 -1562
rect 71532 -1562 71548 -250
rect 71612 -820 71628 -138
rect 76522 -138 76618 -122
rect 78580 -130 79570 -70
rect 74929 -190 76251 -189
rect 76522 -190 76538 -138
rect 73000 -760 73140 -720
rect 73000 -820 73030 -760
rect 71612 -830 73030 -820
rect 73110 -830 73140 -760
rect 71612 -870 73140 -830
rect 71612 -880 73030 -870
rect 71612 -1562 71628 -880
rect 73000 -940 73030 -880
rect 73110 -940 73140 -870
rect 73000 -970 73140 -940
rect 74929 -1510 74930 -190
rect 76250 -250 76538 -190
rect 76250 -1510 76251 -250
rect 74929 -1511 76251 -1510
rect 71532 -1578 71628 -1562
rect 76522 -1562 76538 -250
rect 76602 -820 76618 -138
rect 81242 -138 81338 -122
rect 79649 -190 80971 -189
rect 81242 -190 81258 -138
rect 77990 -760 78130 -720
rect 77990 -820 78020 -760
rect 76602 -830 78020 -820
rect 78100 -830 78130 -760
rect 76602 -870 78130 -830
rect 76602 -880 78020 -870
rect 76602 -1562 76618 -880
rect 77990 -940 78020 -880
rect 78100 -940 78130 -870
rect 77990 -970 78130 -940
rect 79649 -1510 79650 -190
rect 80970 -250 81258 -190
rect 80970 -1510 80971 -250
rect 79649 -1511 80971 -1510
rect 76522 -1578 76618 -1562
rect 81242 -1562 81258 -250
rect 81322 -820 81338 -138
rect 82710 -760 82850 -720
rect 82710 -820 82740 -760
rect 81322 -830 82740 -820
rect 82820 -830 82850 -760
rect 81322 -870 82850 -830
rect 81322 -880 82740 -870
rect 81322 -1562 81338 -880
rect 82710 -940 82740 -880
rect 82820 -940 82850 -870
rect 82710 -970 82850 -940
rect 81242 -1578 81338 -1562
use dum_vert  cap_dum_0 ~/dac_layout
timestamp 1730644682
transform 0 1 18560 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  cap_dum_1
timestamp 1730644682
transform 0 1 43510 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  cap_dum_2
timestamp 1730644682
transform 0 1 48500 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  cap_dum_3
timestamp 1730644682
transform 0 1 53490 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  cap_dum_4
timestamp 1730644682
transform 0 1 58480 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  cap_dum_5
timestamp 1730644682
transform 0 1 63470 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  cap_dum_6
timestamp 1730644682
transform 0 1 68460 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  cap_dum_7
timestamp 1730644682
transform 0 1 73450 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  cap_dum_8
timestamp 1730644682
transform 0 1 78440 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  cap_dum_10
timestamp 1730644682
transform 0 1 8580 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  cap_dum_11
timestamp 1730644682
transform 0 1 13570 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  cap_dum_12
timestamp 1730644682
transform 0 1 38520 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  cap_dum_13
timestamp 1730644682
transform 0 1 23550 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  cap_dum_14
timestamp 1730644682
transform 0 1 28540 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  cap_dum_15
timestamp 1730644682
transform 0 1 33530 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  cap_dum_16
timestamp 1730644682
transform 0 1 -1130 -1 0 25920
box 270 -3590 1980 1130
use dum_vert  dum_vert_0
timestamp 1730644682
transform 0 1 3590 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  dum_vert_1
timestamp 1730644682
transform 0 1 -1130 -1 0 29340
box 270 -3590 1980 1130
use dum_vert  dum_vert_2
timestamp 1730644682
transform 0 1 -1130 -1 0 27630
box 270 -3590 1980 1130
use end  end_0 ~/dac_layout
timestamp 1729689530
transform 0 1 0 -1 0 27360
box 0 0 27360 4720
use end  end_1
timestamp 1729689530
transform 0 1 4990 -1 0 27360
box 0 0 27360 4720
use end  end_2
timestamp 1729689530
transform 0 1 69860 -1 0 27360
box 0 0 27360 4720
use end  end_3
timestamp 1729689530
transform 0 1 74850 -1 0 27360
box 0 0 27360 4720
use mid_2  mid_2_0 ~/dac_layout
timestamp 1729709358
transform 1 0 34930 0 1 13680
box 0 -13680 9800 13680
use mid_2to4_  mid_2to4__0 ~/dac_layout
timestamp 1729683266
transform 0 1 29940 -1 0 27360
box 0 0 27360 4720
use mid_2to4_  mid_2to4__1
timestamp 1729683266
transform 0 1 44910 -1 0 27360
box 0 0 27360 4720
use mid_4to8  mid_4to8_0 ~/dac_layout
timestamp 1729685583
transform 0 1 19960 -1 0 27360
box 0 0 27360 4720
use mid_4to8  mid_4to8_1
timestamp 1729685583
transform 0 1 24950 -1 0 27360
box 0 0 27360 4720
use mid_4to8  mid_4to8_2
timestamp 1729685583
transform 0 1 49900 -1 0 27360
box 0 0 27360 4720
use mid_4to8  mid_4to8_3
timestamp 1729685583
transform 0 1 54890 -1 0 27360
box 0 0 27360 4720
use mid_6to8  mid_6to8_0 ~/dac_layout
timestamp 1729688460
transform 0 1 9980 -1 0 27360
box 0 0 27360 4720
use mid_6to8  mid_6to8_1
timestamp 1729688460
transform 0 1 14970 -1 0 27360
box 0 0 27360 4720
use mid_6to8  mid_6to8_2
timestamp 1729688460
transform 0 1 59880 -1 0 27360
box 0 0 27360 4720
use mid_6to8  mid_6to8_3
timestamp 1729688460
transform 0 1 64870 -1 0 27360
box 0 0 27360 4720
use smpl_switch  smpl_switch_1 ~/dac_layout
timestamp 1730647371
transform 1 0 -5980 0 -1 30210
box -800 -190 1230 30230
<< labels >>
flabel metal1 18630 28046 18632 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 18568 28352 18570 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 13640 28046 13642 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 13578 28352 13580 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 8650 28046 8652 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 8588 28352 8590 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 3660 28046 3662 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 3598 28352 3600 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 38590 28046 38592 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 38528 28352 38530 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 33600 28046 33602 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 33538 28352 33540 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 28610 28046 28612 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 28548 28352 28550 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 23620 28046 23622 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 23558 28352 23560 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 58550 28046 58552 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 58488 28352 58490 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 53560 28046 53562 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 53498 28352 53500 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 48570 28046 48572 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 48508 28352 48510 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 43580 28046 43582 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 43518 28352 43520 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 78510 28046 78512 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 78448 28352 78450 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 73520 28046 73522 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 73458 28352 73460 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 68530 28046 68532 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 68468 28352 68470 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 63540 28046 63542 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 63478 28352 63480 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 17620 28510 17680 28570 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel via1 17730 28350 17790 28410 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel via1 17730 28040 17790 28100 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel metal1 17620 28200 17680 28260 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel metal4 15090 28790 15150 28850 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 18630 28046 18632 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 18568 28352 18570 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 18152 27968 18212 28028 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 18152 28418 18212 28478 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 18690 28190 18750 28240 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 18690 28510 18750 28570 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 12630 28510 12690 28570 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel via1 12740 28350 12800 28410 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel via1 12740 28040 12800 28100 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel metal1 12630 28200 12690 28260 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel metal4 10100 28790 10160 28850 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 13640 28046 13642 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 13578 28352 13580 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 13162 27968 13222 28028 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 13162 28418 13222 28478 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 13700 28190 13760 28240 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 13700 28510 13760 28570 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 7640 28510 7700 28570 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel via1 7750 28350 7810 28410 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel via1 7750 28040 7810 28100 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel metal1 7640 28200 7700 28260 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel metal4 5110 28790 5170 28850 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 8650 28046 8652 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 8588 28352 8590 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 8172 27968 8232 28028 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 8172 28418 8232 28478 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 8710 28190 8770 28240 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 8710 28510 8770 28570 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 2650 28510 2710 28570 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel via1 2760 28350 2820 28410 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel via1 2760 28040 2820 28100 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel metal1 2650 28200 2710 28260 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel metal4 120 28790 180 28850 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 3660 28046 3662 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 3598 28352 3600 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 3182 27968 3242 28028 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 3182 28418 3242 28478 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 3720 28190 3780 28240 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 3720 28510 3780 28570 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 37580 28510 37640 28570 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel via1 37690 28350 37750 28410 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel via1 37690 28040 37750 28100 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel metal1 37580 28200 37640 28260 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel metal4 35050 28790 35110 28850 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 38590 28046 38592 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 38528 28352 38530 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 38112 27968 38172 28028 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 38112 28418 38172 28478 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 38650 28190 38710 28240 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 38650 28510 38710 28570 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 32590 28510 32650 28570 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel via1 32700 28350 32760 28410 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel via1 32700 28040 32760 28100 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel metal1 32590 28200 32650 28260 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel metal4 30060 28790 30120 28850 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 33600 28046 33602 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 33538 28352 33540 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 33122 27968 33182 28028 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 33122 28418 33182 28478 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 33660 28190 33720 28240 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 33660 28510 33720 28570 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 27600 28510 27660 28570 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel via1 27710 28350 27770 28410 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel via1 27710 28040 27770 28100 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel metal1 27600 28200 27660 28260 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel metal4 25070 28790 25130 28850 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 28610 28046 28612 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 28548 28352 28550 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 28132 27968 28192 28028 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 28132 28418 28192 28478 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 28670 28190 28730 28240 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 28670 28510 28730 28570 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 22610 28510 22670 28570 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel via1 22720 28350 22780 28410 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel via1 22720 28040 22780 28100 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel metal1 22610 28200 22670 28260 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel metal4 20080 28790 20140 28850 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 23620 28046 23622 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 23558 28352 23560 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 23142 27968 23202 28028 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 23142 28418 23202 28478 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 23680 28190 23740 28240 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 23680 28510 23740 28570 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 57540 28510 57600 28570 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel via1 57650 28350 57710 28410 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel via1 57650 28040 57710 28100 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel metal1 57540 28200 57600 28260 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel metal4 55010 28790 55070 28850 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 58550 28046 58552 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 58488 28352 58490 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 58072 27968 58132 28028 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 58072 28418 58132 28478 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 58610 28190 58670 28240 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 58610 28510 58670 28570 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 52550 28510 52610 28570 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel via1 52660 28350 52720 28410 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel via1 52660 28040 52720 28100 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel metal1 52550 28200 52610 28260 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel metal4 50020 28790 50080 28850 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 53560 28046 53562 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 53498 28352 53500 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 53082 27968 53142 28028 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 53082 28418 53142 28478 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 53620 28190 53680 28240 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 53620 28510 53680 28570 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 47560 28510 47620 28570 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel via1 47670 28350 47730 28410 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel via1 47670 28040 47730 28100 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel metal1 47560 28200 47620 28260 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel metal4 45030 28790 45090 28850 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 48570 28046 48572 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 48508 28352 48510 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 48092 27968 48152 28028 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 48092 28418 48152 28478 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 48630 28190 48690 28240 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 48630 28510 48690 28570 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 42570 28510 42630 28570 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel via1 42680 28350 42740 28410 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel via1 42680 28040 42740 28100 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel metal1 42570 28200 42630 28260 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel metal4 40040 28790 40100 28850 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 43580 28046 43582 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 43518 28352 43520 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 43102 27968 43162 28028 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 43102 28418 43162 28478 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 43640 28190 43700 28240 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 43640 28510 43700 28570 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 77500 28510 77560 28570 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel via1 77610 28350 77670 28410 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel via1 77610 28040 77670 28100 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel metal1 77500 28200 77560 28260 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel metal4 74970 28790 75030 28850 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 78510 28046 78512 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 78448 28352 78450 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 78032 27968 78092 28028 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 78032 28418 78092 28478 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 78570 28190 78630 28240 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 78570 28510 78630 28570 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 72510 28510 72570 28570 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel via1 72620 28350 72680 28410 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel via1 72620 28040 72680 28100 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel metal1 72510 28200 72570 28260 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel metal4 69980 28790 70040 28850 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 73520 28046 73522 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 73458 28352 73460 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 73042 27968 73102 28028 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 73042 28418 73102 28478 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 73580 28190 73640 28240 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 73580 28510 73640 28570 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 67520 28510 67580 28570 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel via1 67630 28350 67690 28410 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel via1 67630 28040 67690 28100 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel metal1 67520 28200 67580 28260 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel metal4 64990 28790 65050 28850 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 68530 28046 68532 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 68468 28352 68470 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 68052 27968 68112 28028 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 68052 28418 68112 28478 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 68590 28190 68650 28240 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 68590 28510 68650 28570 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 62530 28510 62590 28570 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel via1 62640 28350 62700 28410 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel via1 62640 28040 62700 28100 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel metal1 62530 28200 62590 28260 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel metal4 60000 28790 60060 28850 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 63540 28046 63542 28106 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal1 63478 28352 63480 28412 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 63062 27968 63122 28028 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 63062 28418 63122 28478 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 63600 28190 63660 28240 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 63600 28510 63660 28570 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 63600 -560 63660 -500 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 63600 -880 63660 -830 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 63062 -652 63122 -592 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 63062 -1102 63122 -1042 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 63478 -718 63480 -658 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 63540 -1024 63542 -964 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal4 60000 -280 60060 -220 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 62530 -870 62590 -810 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel via1 62640 -1030 62700 -970 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel via1 62640 -720 62700 -660 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel metal1 62530 -560 62590 -500 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel metal1 68590 -560 68650 -500 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 68590 -880 68650 -830 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 68052 -652 68112 -592 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 68052 -1102 68112 -1042 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 68468 -718 68470 -658 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 68530 -1024 68532 -964 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal4 64990 -280 65050 -220 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 67520 -870 67580 -810 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel via1 67630 -1030 67690 -970 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel via1 67630 -720 67690 -660 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel metal1 67520 -560 67580 -500 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel metal1 73580 -560 73640 -500 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 73580 -880 73640 -830 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 73042 -652 73102 -592 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 73042 -1102 73102 -1042 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 73458 -718 73460 -658 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 73520 -1024 73522 -964 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal4 69980 -280 70040 -220 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 72510 -870 72570 -810 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel via1 72620 -1030 72680 -970 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel via1 72620 -720 72680 -660 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel metal1 72510 -560 72570 -500 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel metal1 78570 -560 78630 -500 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 78570 -880 78630 -830 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 78032 -652 78092 -592 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 78032 -1102 78092 -1042 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 78448 -718 78450 -658 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 78510 -1024 78512 -964 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal4 74970 -280 75030 -220 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 77500 -870 77560 -810 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel via1 77610 -1030 77670 -970 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel via1 77610 -720 77670 -660 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel metal1 77500 -560 77560 -500 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel metal1 43640 -560 43700 -500 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 43640 -880 43700 -830 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 43102 -652 43162 -592 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 43102 -1102 43162 -1042 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 43518 -718 43520 -658 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 43580 -1024 43582 -964 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal4 40040 -280 40100 -220 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 42570 -870 42630 -810 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel via1 42680 -1030 42740 -970 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel via1 42680 -720 42740 -660 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel metal1 42570 -560 42630 -500 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel metal1 48630 -560 48690 -500 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 48630 -880 48690 -830 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 48092 -652 48152 -592 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 48092 -1102 48152 -1042 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 48508 -718 48510 -658 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 48570 -1024 48572 -964 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal4 45030 -280 45090 -220 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 47560 -870 47620 -810 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel via1 47670 -1030 47730 -970 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel via1 47670 -720 47730 -660 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel metal1 47560 -560 47620 -500 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel metal1 53620 -560 53680 -500 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 53620 -880 53680 -830 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 53082 -652 53142 -592 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 53082 -1102 53142 -1042 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 53498 -718 53500 -658 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 53560 -1024 53562 -964 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal4 50020 -280 50080 -220 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 52550 -870 52610 -810 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel via1 52660 -1030 52720 -970 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel via1 52660 -720 52720 -660 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel metal1 52550 -560 52610 -500 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel metal1 58610 -560 58670 -500 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 58610 -880 58670 -830 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 58072 -652 58132 -592 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 58072 -1102 58132 -1042 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 58488 -718 58490 -658 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 58550 -1024 58552 -964 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal4 55010 -280 55070 -220 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 57540 -870 57600 -810 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel via1 57650 -1030 57710 -970 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel via1 57650 -720 57710 -660 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel metal1 57540 -560 57600 -500 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel metal1 23680 -560 23740 -500 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 23680 -880 23740 -830 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 23142 -652 23202 -592 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 23142 -1102 23202 -1042 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 23558 -718 23560 -658 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 23620 -1024 23622 -964 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal4 20080 -280 20140 -220 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 22610 -870 22670 -810 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel via1 22720 -1030 22780 -970 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel via1 22720 -720 22780 -660 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel metal1 22610 -560 22670 -500 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel metal1 28670 -560 28730 -500 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 28670 -880 28730 -830 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 28132 -652 28192 -592 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 28132 -1102 28192 -1042 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 28548 -718 28550 -658 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 28610 -1024 28612 -964 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal4 25070 -280 25130 -220 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 27600 -870 27660 -810 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel via1 27710 -1030 27770 -970 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel via1 27710 -720 27770 -660 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel metal1 27600 -560 27660 -500 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel metal1 33660 -560 33720 -500 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 33660 -880 33720 -830 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 33122 -652 33182 -592 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 33122 -1102 33182 -1042 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 33538 -718 33540 -658 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 33600 -1024 33602 -964 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal4 30060 -280 30120 -220 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 32590 -870 32650 -810 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel via1 32700 -1030 32760 -970 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel via1 32700 -720 32760 -660 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel metal1 32590 -560 32650 -500 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel metal1 38650 -560 38710 -500 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 38650 -880 38710 -830 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 38112 -652 38172 -592 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 38112 -1102 38172 -1042 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 38528 -718 38530 -658 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 38590 -1024 38592 -964 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal4 35050 -280 35110 -220 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 37580 -870 37640 -810 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel via1 37690 -1030 37750 -970 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel via1 37690 -720 37750 -660 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel metal1 37580 -560 37640 -500 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel metal1 3720 -560 3780 -500 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 3720 -880 3780 -830 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 3182 -652 3242 -592 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 3182 -1102 3242 -1042 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 3598 -718 3600 -658 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 3660 -1024 3662 -964 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal4 120 -280 180 -220 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 2650 -870 2710 -810 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel via1 2760 -1030 2820 -970 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel via1 2760 -720 2820 -660 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel metal1 2650 -560 2710 -500 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel metal1 8710 -560 8770 -500 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 8710 -880 8770 -830 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 8172 -652 8232 -592 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 8172 -1102 8232 -1042 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 8588 -718 8590 -658 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 8650 -1024 8652 -964 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal4 5110 -280 5170 -220 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 7640 -870 7700 -810 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel via1 7750 -1030 7810 -970 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel via1 7750 -720 7810 -660 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel metal1 7640 -560 7700 -500 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel metal1 13700 -560 13760 -500 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 13700 -880 13760 -830 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 13162 -652 13222 -592 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 13162 -1102 13222 -1042 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 13578 -718 13580 -658 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 13640 -1024 13642 -964 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal4 10100 -280 10160 -220 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 12630 -870 12690 -810 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel via1 12740 -1030 12800 -970 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel via1 12740 -720 12800 -660 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel metal1 12630 -560 12690 -500 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel metal1 18690 -560 18750 -500 0 FreeSans 256 90 0 0 Vdd
port 3 nsew
flabel metal1 18690 -880 18750 -830 0 FreeSans 256 90 0 0 Vdd
port 7 nsew
flabel metal1 18152 -652 18212 -592 0 FreeSans 256 90 0 0 Vin
port 5 nsew
flabel metal1 18152 -1102 18212 -1042 0 FreeSans 256 90 0 0 GND
port 9 nsew
flabel metal1 18568 -718 18570 -658 0 FreeSans 256 90 0 0 phi1_n
port 4 nsew
flabel metal1 18630 -1024 18632 -964 0 FreeSans 256 90 0 0 phi2_n
port 10 nsew
flabel metal4 15090 -280 15150 -220 0 FreeSans 256 90 0 0 com_x
port 0 nsew
flabel metal1 17620 -870 17680 -810 0 FreeSans 256 90 0 0 sub
port 1 nsew
flabel via1 17730 -1030 17790 -970 0 FreeSans 256 90 0 0 phi2
port 8 nsew
flabel via1 17730 -720 17790 -660 0 FreeSans 256 90 0 0 phi1
port 2 nsew
flabel metal1 17620 -560 17680 -500 0 FreeSans 256 90 0 0 sub
port 6 nsew
flabel metal3 -4974 29924 -4864 29974 0 FreeSans 160 0 0 0 sub
port 14 nsew
flabel metal3 -4970 30212 -4866 30266 0 FreeSans 160 0 0 0 sphi1
port 22 nsew
flabel metal3 -4976 30354 -4872 30408 0 FreeSans 160 0 0 0 sphi2
port 24 nsew
flabel metal3 -4982 30492 -4874 30542 0 FreeSans 160 0 0 0 phi10
port 26 nsew
flabel metal3 -4974 30636 -4866 30686 0 FreeSans 160 0 0 0 phi20
port 28 nsew
flabel metal3 -4972 30776 -4864 30826 0 FreeSans 160 0 0 0 phi11
port 30 nsew
flabel metal3 -4970 30914 -4862 30964 0 FreeSans 160 0 0 0 phi21
port 32 nsew
flabel metal3 -4974 31054 -4866 31104 0 FreeSans 160 0 0 0 phi12
port 34 nsew
flabel metal3 -4980 31194 -4872 31244 0 FreeSans 160 0 0 0 phi22
port 36 nsew
flabel metal3 -4968 31336 -4860 31386 0 FreeSans 160 0 0 0 phi13
port 38 nsew
flabel metal3 -4956 31474 -4848 31524 0 FreeSans 160 0 0 0 phi23
port 40 nsew
flabel metal3 -4958 31618 -4850 31668 0 FreeSans 160 0 0 0 phi14
port 42 nsew
flabel metal3 -4954 31756 -4846 31806 0 FreeSans 160 0 0 0 phi24
port 44 nsew
flabel metal3 -4954 31896 -4846 31946 0 FreeSans 160 0 0 0 phi15
port 46 nsew
flabel metal3 -4950 32032 -4842 32082 0 FreeSans 160 0 0 0 phi25
port 48 nsew
flabel metal3 -4952 32172 -4844 32222 0 FreeSans 160 0 0 0 phi16
port 50 nsew
flabel metal3 -4954 32314 -4846 32364 0 FreeSans 160 0 0 0 phi26
port 52 nsew
flabel metal3 -4950 32454 -4842 32504 0 FreeSans 160 0 0 0 phi17
port 54 nsew
flabel metal3 -4946 32594 -4838 32644 0 FreeSans 160 0 0 0 phi27
port 56 nsew
flabel metal1 -4822 29920 -4730 29944 0 FreeSans 160 0 0 0 gnd
port 58 nsew
flabel metal1 -4798 30214 -4706 30240 0 FreeSans 160 0 0 0 sphi1_n
port 64 nsew
flabel metal1 -4800 30350 -4708 30376 0 FreeSans 160 0 0 0 sphi2_n
port 66 nsew
flabel metal1 -4802 30490 -4710 30516 0 FreeSans 160 0 0 0 phi1_n0
port 68 nsew
flabel metal1 -4802 30632 -4710 30658 0 FreeSans 160 0 0 0 phi2_n0
port 70 nsew
flabel metal1 -4802 30770 -4710 30796 0 FreeSans 160 0 0 0 phi1_n1
port 72 nsew
flabel metal1 -4800 30912 -4708 30938 0 FreeSans 160 0 0 0 phi2_n1
port 74 nsew
flabel metal1 -4798 31050 -4706 31076 0 FreeSans 160 0 0 0 phi1_n2
port 76 nsew
flabel metal1 -4796 31192 -4704 31218 0 FreeSans 160 0 0 0 phi2_n2
port 78 nsew
flabel metal1 -4794 31332 -4702 31358 0 FreeSans 160 0 0 0 phi1_n3
port 80 nsew
flabel metal1 -4792 31472 -4700 31498 0 FreeSans 160 0 0 0 phi2_n3
port 82 nsew
flabel metal1 -4792 31612 -4700 31638 0 FreeSans 160 0 0 0 phi1_n4
port 84 nsew
flabel metal1 -4790 31752 -4698 31778 0 FreeSans 160 0 0 0 phi2_n4
port 86 nsew
flabel metal1 -4788 31892 -4696 31918 0 FreeSans 160 0 0 0 phi1_n5
port 88 nsew
flabel metal1 -4786 32032 -4694 32058 0 FreeSans 160 0 0 0 phi2_n5
port 90 nsew
flabel metal1 -4794 32170 -4702 32196 0 FreeSans 160 0 0 0 phi1_n6
port 92 nsew
flabel metal1 -4798 32310 -4706 32336 0 FreeSans 160 0 0 0 phi2_n6
port 94 nsew
flabel metal1 -4794 32452 -4702 32478 0 FreeSans 160 0 0 0 phi1_n7
port 96 nsew
flabel metal1 -4790 32592 -4698 32618 0 FreeSans 160 0 0 0 phi2_n7
port 98 nsew
flabel metal1 -4812 30062 -4720 30088 0 FreeSans 160 0 0 0 vin
port 60 nsew
flabel metal3 -4972 30066 -4862 30116 0 FreeSans 160 0 0 0 vdd
port 18 nsew
<< end >>
