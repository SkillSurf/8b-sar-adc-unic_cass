magic
tech sky130A
magscale 1 2
timestamp 1730665161
<< nwell >>
rect 910 0 1010 80
<< pwell >>
rect 910 -840 1010 -760
<< locali >>
rect 710 180 1190 200
rect 710 140 840 180
rect 1080 140 1190 180
rect 710 110 1190 140
rect 710 -890 1140 -860
rect 710 -930 840 -890
rect 1080 -930 1140 -890
rect 710 -950 1140 -930
<< viali >>
rect 840 140 1080 180
rect 840 -930 1080 -890
<< metal1 >>
rect 670 180 1230 200
rect 670 140 840 180
rect 1080 140 1230 180
rect 670 130 1230 140
rect 910 10 930 70
rect 990 10 1010 70
rect 900 -340 930 -220
rect 850 -350 930 -340
rect 850 -410 860 -350
rect 920 -410 930 -350
rect 850 -420 930 -410
rect 900 -540 930 -420
rect 990 -330 1020 -220
rect 990 -340 1110 -330
rect 990 -410 1030 -340
rect 1100 -410 1110 -340
rect 990 -420 1110 -410
rect 990 -540 1020 -420
rect 910 -830 930 -760
rect 990 -830 1010 -760
rect 910 -840 1010 -830
rect 670 -890 1180 -880
rect 670 -930 840 -890
rect 1080 -930 1180 -890
rect 670 -950 1180 -930
<< via1 >>
rect 930 10 990 70
rect 860 -410 920 -350
rect 1030 -410 1100 -340
rect 930 -830 990 -760
<< metal2 >>
rect 710 230 1200 260
rect 850 -340 880 230
rect 920 10 930 70
rect 990 10 1000 70
rect 850 -350 930 -340
rect 850 -410 860 -350
rect 920 -410 930 -350
rect 850 -420 930 -410
rect 960 -700 990 10
rect 1020 -340 1110 -330
rect 1020 -410 1030 -340
rect 1100 -410 1110 -340
rect 1020 -420 1110 -410
rect 960 -730 1060 -700
rect 920 -830 930 -760
rect 990 -830 1000 -760
rect 920 -840 1000 -830
rect 950 -970 980 -840
rect 1030 -970 1060 -730
<< via2 >>
rect 1030 -410 1090 -350
<< metal3 >>
rect 1020 -340 1140 -330
rect 1020 -410 1030 -340
rect 1100 -410 1140 -340
rect 1020 -420 1140 -410
<< via3 >>
rect 1030 -350 1100 -340
rect 1030 -410 1090 -350
rect 1090 -410 1100 -350
<< metal4 >>
rect 1020 -340 1140 -330
rect 1020 -410 1030 -340
rect 1100 -400 1350 -340
rect 1100 -410 1140 -400
rect 1020 -420 1140 -410
use sky130_fd_pr__pfet_01v8_NKK3FE  XM1 ~/final
timestamp 1728804544
transform 1 0 961 0 1 -96
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_5WP7M2  XM2 ~/final
timestamp 1730665161
transform 1 0 961 0 1 -661
box -211 -279 211 279
<< labels >>
flabel metal1 770 130 830 190 0 FreeSans 256 0 0 0 Vdd
port 3 nsew
flabel metal1 862 -408 922 -348 0 FreeSans 256 0 0 0 Vin
port 5 nsew
flabel metal1 770 -940 830 -880 0 FreeSans 256 0 0 0 sub
port 6 nsew
rlabel metal1 910 -840 920 -760 1 clk
port 7 n
rlabel metal1 1000 10 1010 70 1 clk_b
port 8 n
rlabel metal1 990 -410 1020 -380 1 Vout
port 9 n
<< end >>
