magic
tech sky130A
magscale 1 2
timestamp 1729222717
<< checkpaint >>
rect 16799 3404 19911 3457
rect 16799 -1737 20450 3404
rect 17338 -1790 20450 -1737
rect 31791 -2951 34903 2243
<< error_s >>
rect 2346 6153 2381 6187
rect 2347 6134 2381 6153
rect 468 5023 503 5057
rect 1061 5040 1095 5058
rect 469 5004 503 5023
rect 488 -17 503 5004
rect 522 4970 557 5004
rect 522 -17 556 4970
rect 522 -51 537 -17
rect 1025 -70 1095 5040
rect 1025 -106 1078 -70
rect 2366 -123 2381 6134
rect 2400 6100 2435 6134
rect 2400 -123 2434 6100
rect 18580 2127 18615 2161
rect 18581 2108 18615 2127
rect 3686 1573 3720 1591
rect 3686 1537 3756 1573
rect 3703 1503 3774 1537
rect 2400 -157 2415 -123
rect 3703 -176 3773 1503
rect 3703 -212 3756 -176
rect 8044 -229 8059 1537
rect 8078 -229 8112 1591
rect 12364 613 12398 667
rect 16756 649 16790 667
rect 8078 -263 8093 -229
rect 12383 -282 12398 613
rect 12417 579 12452 613
rect 12417 -282 12451 579
rect 12417 -316 12432 -282
rect 16720 -335 16790 649
rect 16720 -371 16773 -335
rect 18061 -388 18076 978
rect 18095 -388 18129 1032
rect 18095 -422 18110 -388
rect 18600 -441 18615 2108
rect 18634 2074 18669 2108
rect 18634 -441 18668 2074
rect 31695 1036 31729 1054
rect 31695 1000 31765 1036
rect 31712 966 31783 1000
rect 21016 679 21051 713
rect 21017 660 21051 679
rect 20815 611 20887 617
rect 20815 577 20827 611
rect 20815 571 20887 577
rect 19120 437 19154 455
rect 19120 401 19190 437
rect 19137 367 19208 401
rect 19858 367 19893 401
rect 20651 384 20685 402
rect 18634 -475 18649 -441
rect 19137 -494 19207 367
rect 19859 348 19893 367
rect 19137 -530 19190 -494
rect 19878 -547 19893 348
rect 19912 314 19947 348
rect 19912 -547 19946 314
rect 19912 -581 19927 -547
rect 20615 -600 20685 384
rect 20815 -517 20887 -511
rect 20815 -551 20827 -517
rect 20815 -557 20887 -551
rect 20615 -636 20668 -600
rect 21036 -653 21051 660
rect 21070 626 21105 660
rect 21070 -653 21104 626
rect 21234 558 21306 564
rect 21234 524 21246 558
rect 21234 518 21306 524
rect 24806 149 24841 183
rect 24807 130 24841 149
rect 24605 81 24677 87
rect 24605 47 24617 81
rect 24605 41 24677 47
rect 23111 -71 23169 -65
rect 23111 -105 23123 -71
rect 23111 -111 23169 -105
rect 23281 -222 23315 -204
rect 21436 -275 21470 -257
rect 23281 -258 23351 -222
rect 21436 -311 21506 -275
rect 23298 -292 23369 -258
rect 21453 -345 21524 -311
rect 21804 -345 21839 -311
rect 22227 -328 22262 -310
rect 21234 -570 21306 -564
rect 21234 -604 21246 -570
rect 21234 -610 21306 -604
rect 21070 -687 21085 -653
rect 21453 -706 21523 -345
rect 21805 -364 21839 -345
rect 22191 -333 22262 -328
rect 21635 -413 21693 -407
rect 21635 -447 21647 -413
rect 21635 -453 21693 -447
rect 21635 -623 21693 -617
rect 21635 -657 21647 -623
rect 21635 -663 21693 -657
rect 21453 -742 21506 -706
rect 21824 -759 21839 -364
rect 21858 -398 21893 -364
rect 21858 -759 21892 -398
rect 22004 -466 22062 -460
rect 22004 -500 22016 -466
rect 22004 -506 22062 -500
rect 22004 -676 22062 -670
rect 22004 -710 22016 -676
rect 22004 -716 22062 -710
rect 21858 -793 21873 -759
rect 22191 -812 22261 -333
rect 22373 -401 22431 -395
rect 23111 -399 23169 -393
rect 22373 -435 22385 -401
rect 22543 -434 22577 -416
rect 22965 -434 22999 -416
rect 22373 -441 22431 -435
rect 22543 -470 22613 -434
rect 22560 -504 22631 -470
rect 22373 -729 22431 -723
rect 22373 -763 22385 -729
rect 22373 -769 22431 -763
rect 22191 -848 22244 -812
rect 22560 -865 22630 -504
rect 22742 -572 22800 -566
rect 22742 -606 22754 -572
rect 22742 -612 22800 -606
rect 22742 -782 22800 -776
rect 22742 -816 22754 -782
rect 22742 -822 22800 -816
rect 22560 -901 22613 -865
rect 22929 -918 22999 -434
rect 23111 -433 23123 -399
rect 23111 -439 23169 -433
rect 23111 -507 23169 -501
rect 23111 -541 23123 -507
rect 23111 -547 23169 -541
rect 23111 -835 23169 -829
rect 23111 -869 23123 -835
rect 23111 -875 23169 -869
rect 22929 -954 22982 -918
rect 23298 -971 23368 -292
rect 23480 -360 23538 -354
rect 23480 -394 23492 -360
rect 23480 -400 23538 -394
rect 23650 -475 23684 -457
rect 23650 -511 23720 -475
rect 23667 -545 23738 -511
rect 23480 -570 23538 -564
rect 23480 -604 23492 -570
rect 23480 -610 23538 -604
rect 23480 -678 23538 -672
rect 23480 -712 23492 -678
rect 23480 -718 23538 -712
rect 23480 -888 23538 -882
rect 23480 -922 23492 -888
rect 23480 -928 23538 -922
rect 23298 -1007 23351 -971
rect 23667 -1024 23737 -545
rect 23849 -613 23907 -607
rect 23849 -647 23861 -613
rect 24019 -646 24053 -628
rect 24441 -646 24475 -628
rect 23849 -653 23907 -647
rect 24019 -682 24089 -646
rect 24036 -716 24107 -682
rect 23849 -941 23907 -935
rect 23849 -975 23861 -941
rect 23849 -981 23907 -975
rect 23667 -1060 23720 -1024
rect 24036 -1077 24106 -716
rect 24218 -784 24276 -778
rect 24218 -818 24230 -784
rect 24218 -824 24276 -818
rect 24218 -994 24276 -988
rect 24218 -1028 24230 -994
rect 24218 -1034 24276 -1028
rect 24036 -1113 24089 -1077
rect 24405 -1130 24475 -646
rect 24605 -1047 24677 -1041
rect 24605 -1081 24617 -1047
rect 24605 -1087 24677 -1081
rect 24405 -1166 24458 -1130
rect 24826 -1183 24841 130
rect 24860 96 24895 130
rect 24860 -1183 24894 96
rect 25024 28 25096 34
rect 25024 -6 25036 28
rect 25024 -12 25096 -6
rect 30617 -130 30651 -76
rect 25226 -705 25260 -687
rect 25226 -741 25296 -705
rect 25243 -775 25314 -741
rect 25594 -775 25629 -741
rect 25024 -1100 25096 -1094
rect 25024 -1134 25036 -1100
rect 25024 -1140 25096 -1134
rect 24860 -1217 24875 -1183
rect 25243 -1236 25313 -775
rect 25595 -794 25629 -775
rect 25425 -843 25483 -837
rect 25425 -877 25437 -843
rect 25425 -883 25483 -877
rect 25425 -1153 25483 -1147
rect 25425 -1187 25437 -1153
rect 25425 -1193 25483 -1187
rect 25243 -1272 25296 -1236
rect 25614 -1289 25629 -794
rect 25648 -828 25683 -794
rect 26331 -796 26344 -783
rect 25648 -1289 25682 -828
rect 25794 -896 25852 -890
rect 25794 -930 25806 -896
rect 25794 -936 25852 -930
rect 25996 -1117 26034 -796
rect 26295 -1117 26348 -796
rect 25794 -1206 25852 -1200
rect 25794 -1240 25806 -1206
rect 25794 -1246 25852 -1240
rect 25648 -1323 25663 -1289
rect 26297 -1395 26310 -1361
rect 26331 -1429 26344 -1327
rect 30636 -1443 30651 -130
rect 30670 -164 30705 -130
rect 30670 -1443 30704 -164
rect 30670 -1477 30685 -1443
rect 31175 -1496 31190 -130
rect 31209 -1496 31243 -76
rect 31209 -1530 31224 -1496
rect 31712 -1549 31782 966
rect 31712 -1585 31765 -1549
use sky130_fd_sc_hd__inv_1  x30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 26034 0 1 -1378
box -38 -48 314 592
use sky130_fd_pr__pfet_01v8_lvt_EHBMNA  XM1
timestamp 0
transform 1 0 3060 0 1 2979
box -696 -3191 696 3191
use sky130_fd_pr__pfet_01v8_lvt_EHBMNA  XM2
timestamp 0
transform 1 0 1721 0 1 3032
box -696 -3191 696 3191
use sky130_fd_pr__nfet_01v8_lvt_YJMECZ  XM3
timestamp 0
transform 1 0 243 0 1 2520
box -296 -2573 296 2573
use sky130_fd_pr__nfet_01v8_lvt_YJMECZ  XM4
timestamp 0
transform 1 0 782 0 1 2467
box -296 -2573 296 2573
use sky130_fd_pr__nfet_01v8_542FHV  XM5
timestamp 0
transform 1 0 10238 0 1 4691
box -2196 -5009 2196 5009
use sky130_fd_pr__nfet_01v8_WH99ML  XM6
timestamp 0
transform 1 0 5899 0 1 654
box -2196 -919 2196 919
use sky130_fd_pr__nfet_01v8_H2YH6E  XM7
timestamp 0
transform 1 0 14577 0 1 139
box -2196 -510 2196 510
use sky130_fd_pr__pfet_01v8_lvt_5LG8TG  XM8
timestamp 0
transform 1 0 17416 0 1 295
box -696 -719 696 719
use sky130_fd_pr__pfet_01v8_lvt_FHTFBK  XM9
timestamp 0
transform 1 0 18355 0 1 860
box -296 -1337 296 1337
use sky130_fd_pr__pfet_01v8_lvt_FHTFBK  XM10
timestamp 0
transform 1 0 18894 0 1 807
box -296 -1337 296 1337
use sky130_fd_pr__nfet_01v8_Q9QDRV  XM11
timestamp 0
transform 1 0 19533 0 1 -73
box -396 -510 396 510
use sky130_fd_pr__nfet_01v8_Q9QDRV  XM12
timestamp 0
transform 1 0 20272 0 1 -126
box -396 -510 396 510
use sky130_fd_pr__pfet_01v8_lvt_FMK5UC  XM13
timestamp 0
transform 1 0 20851 0 1 30
box -236 -719 236 719
use sky130_fd_pr__pfet_01v8_lvt_FMK5UC  XM14
timestamp 0
transform 1 0 21270 0 1 -23
box -236 -719 236 719
use sky130_fd_pr__pfet_01v8_lvt_FMK5UC  XM15
timestamp 0
transform 1 0 24641 0 1 -500
box -236 -719 236 719
use sky130_fd_pr__pfet_01v8_lvt_FMK5UC  XM16
timestamp 0
transform 1 0 25060 0 1 -553
box -236 -719 236 719
use sky130_fd_pr__nfet_01v8_QWUGQF  XM17
timestamp 0
transform 1 0 21664 0 1 -535
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_QWUGQF  XM18
timestamp 0
transform 1 0 22033 0 1 -588
box -211 -260 211 260
use sky130_fd_pr__pfet_01v8_J8PPQP  XM19
timestamp 0
transform 1 0 22402 0 1 -582
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_QWUGQF  XM20
timestamp 0
transform 1 0 22771 0 1 -694
box -211 -260 211 260
use sky130_fd_pr__pfet_01v8_NR67KK  XM21
timestamp 0
transform 1 0 23140 0 1 -470
box -211 -537 211 537
use sky130_fd_pr__nfet_01v8_A23HQP  XM22
timestamp 0
transform 1 0 23509 0 1 -641
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_J8PPQP  XM23
timestamp 0
transform 1 0 23878 0 1 -794
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_QWUGQF  XM24
timestamp 0
transform 1 0 24247 0 1 -906
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_lvt_TGNW9T  XM25
timestamp 0
transform 1 0 25454 0 1 -1015
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_lvt_TGNW9T  XM26
timestamp 0
transform 1 0 25823 0 1 -1068
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_WH99ML  XM27
timestamp 0
transform 1 0 28491 0 1 -560
box -2196 -919 2196 919
use sky130_fd_pr__nfet_01v8_lvt_4HYZBZ  XM28
timestamp 0
transform 1 0 30930 0 1 -813
box -296 -719 296 719
use sky130_fd_pr__nfet_01v8_lvt_NRMQA7  XM29
timestamp 0
transform 1 0 31469 0 1 2696
box -296 -4281 296 4281
use sky130_fd_pr__pfet_01v8_lvt_JHTFBT  XM30
timestamp 0
transform 1 0 32408 0 1 -301
box -696 -1337 696 1337
use sky130_fd_pr__pfet_01v8_lvt_FHTFBK  XM31
timestamp 0
transform 1 0 33347 0 1 -354
box -296 -1337 296 1337
<< end >>
