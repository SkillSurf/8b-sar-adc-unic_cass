* SPICE3 file created from dac_top.ext - technology: sky130A

X0 mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1 mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2 mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3 mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X5 mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=74.24 ps=660.48 w=1 l=0.15
X6 mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=74.24 ps=660.48 w=1 l=0.15
X7 mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=74.24 ps=660.48 w=1 l=0.15
X8 mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=74.24 ps=660.48 w=1 l=0.15
X9 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X10 mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X11 mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X12 mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X13 mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X14 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X15 mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X16 mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X17 mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X18 mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X19 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X20 mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X21 mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X22 mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X23 mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X24 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X25 mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X26 mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X27 mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X28 mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X29 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X30 mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X31 mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X32 mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X33 mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X34 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X35 mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X36 mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X37 mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X38 mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X39 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X40 mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X41 mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X42 mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X43 mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X44 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X45 mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X46 mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X47 mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X48 mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X49 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X50 mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X51 mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X52 mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X53 mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X54 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X55 mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X56 mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X57 mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X58 mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X59 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X60 mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X61 mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X62 mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X63 mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X64 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X65 mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X66 mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X67 mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X68 mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X69 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X70 mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X71 mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X72 mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X73 mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X74 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X75 mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X76 mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X77 mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X78 mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X79 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X80 mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X81 mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X82 mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X83 mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X84 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X85 mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X86 mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X87 mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X88 mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X89 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X90 mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X91 mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X92 mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X93 mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X94 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X95 mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X96 mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X97 mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X98 mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X99 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X100 mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X101 mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X102 mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X103 mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X104 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X105 mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X106 mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X107 mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X108 mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X109 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X110 mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X111 mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X112 mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X113 mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X114 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X115 mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X116 mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X117 mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X118 mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X119 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X120 mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X121 mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X122 mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X123 mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X124 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X125 mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X126 mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X127 mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X128 mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X129 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X130 mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X131 mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X132 mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X133 mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X134 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X135 mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X136 mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X137 mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X138 mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X139 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X140 mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X141 mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X142 mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X143 mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X144 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X145 mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X146 mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X147 mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X148 mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X149 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X150 mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X151 mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X152 mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X153 mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X154 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X155 mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X156 mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X157 mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X158 mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X159 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X160 mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X161 mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X162 mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X163 mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X164 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X165 mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X166 mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X167 mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X168 mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X169 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X170 mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X171 mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X172 mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X173 mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X174 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X175 mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X176 mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X177 mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X178 mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X179 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X180 mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X181 mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X182 mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X183 mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X184 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X185 mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X186 mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X187 mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X188 mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X189 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X190 mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X191 mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X192 mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X193 mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X194 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X195 mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X196 mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X197 mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X198 mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X199 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X200 mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X201 mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X202 mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X203 mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X204 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X205 mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X206 mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X207 mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X208 mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X209 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X210 mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X211 mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X212 mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X213 mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X214 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X215 mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X216 mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X217 mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X218 mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X219 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X220 mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X221 mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X222 mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X223 mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X224 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X225 mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X226 mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X227 mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X228 mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X229 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X230 mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X231 mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X232 mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X233 mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X234 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X235 mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X236 mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X237 mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X238 mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X239 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X240 mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X241 mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X242 mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X243 mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X244 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X245 mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X246 mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X247 mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X248 mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X249 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X250 mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X251 mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X252 mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X253 mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X254 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X255 mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X256 mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X257 mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X258 mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X259 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X260 mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X261 mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X262 mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X263 mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X264 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X265 mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X266 mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X267 mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X268 mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X269 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X270 mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X271 mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X272 mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X273 mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X274 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X275 mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X276 mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X277 mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X278 mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X279 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X280 mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X281 mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X282 mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X283 mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X284 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X285 mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X286 mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X287 mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X288 mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X289 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X290 mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X291 mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X292 mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X293 mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X294 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X295 mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X296 mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X297 mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X298 mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X299 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X300 mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X301 mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X302 mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X303 mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X304 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X305 mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X306 mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X307 mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X308 mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X309 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X310 mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X311 mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X312 mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X313 mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X314 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X315 mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X316 mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X317 mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X318 mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X319 end_3/8_cap_array_final_1/cap_final_7/com_x mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X320 mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X321 mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X322 mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X323 mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X324 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X325 mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X326 mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X327 mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X328 mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X329 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X330 mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X331 mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X332 mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X333 mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X334 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X335 mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X336 mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X337 mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X338 mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X339 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X340 mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X341 mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X342 mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X343 mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X344 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X345 mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X346 mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X347 mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X348 mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X349 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X350 mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X351 mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X352 mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X353 mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X354 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X355 mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X356 mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X357 mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X358 mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X359 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X360 mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X361 mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X362 mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X363 mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X364 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X365 mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X366 mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X367 mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X368 mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X369 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X370 mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X371 mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X372 mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X373 mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X374 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X375 mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X376 mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X377 mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X378 mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X379 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X380 mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X381 mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X382 mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X383 mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X384 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X385 mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X386 mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X387 mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X388 mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X389 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X390 mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X391 mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X392 mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X393 mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X394 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X395 mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X396 mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X397 mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X398 mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X399 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X400 mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X401 mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X402 mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X403 mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X404 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X405 mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X406 mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X407 mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X408 mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X409 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X410 mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X411 mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X412 mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X413 mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X414 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X415 mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X416 mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X417 mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X418 mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X419 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X420 mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X421 mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X422 mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X423 mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X424 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X425 mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X426 mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X427 mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X428 mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X429 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X430 mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X431 mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X432 mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X433 mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X434 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X435 mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X436 mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X437 mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X438 mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X439 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X440 mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X441 mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X442 mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X443 mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X444 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X445 mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X446 mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X447 mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X448 mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X449 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X450 mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X451 mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X452 mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X453 mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X454 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X455 mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X456 mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X457 mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X458 mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X459 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X460 mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X461 mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X462 mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X463 mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X464 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X465 mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X466 mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X467 mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X468 mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X469 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X470 mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X471 mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X472 mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X473 mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X474 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X475 mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X476 mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X477 mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X478 mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X479 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X480 mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X481 mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X482 mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X483 mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X484 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X485 mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X486 mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X487 mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X488 mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X489 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X490 mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X491 mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X492 mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X493 mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X494 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X495 mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X496 mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X497 mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X498 mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X499 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X500 mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X501 mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X502 mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X503 mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X504 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X505 mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X506 mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X507 mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X508 mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X509 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X510 mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X511 mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X512 mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X513 mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X514 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X515 mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X516 mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X517 mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X518 mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X519 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X520 mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X521 mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X522 mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X523 mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X524 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X525 mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X526 mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X527 mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X528 mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X529 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X530 mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X531 mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X532 mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X533 mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X534 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X535 mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X536 mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X537 mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X538 mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X539 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X540 mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X541 mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X542 mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X543 mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X544 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X545 mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X546 mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X547 mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X548 mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X549 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X550 mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X551 mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X552 mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X553 mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X554 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X555 mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X556 mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X557 mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X558 mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X559 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X560 end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X561 end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X562 end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X563 end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X564 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X565 end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X566 end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X567 end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X568 end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X569 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X570 end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X571 end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X572 end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X573 end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X574 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X575 end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X576 end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X577 end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X578 end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X579 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X580 end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X581 end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X582 end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X583 end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X584 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X585 end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X586 end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X587 end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X588 end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X589 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X590 end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X591 end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X592 end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X593 end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X594 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X595 end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X596 end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X597 end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X598 end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X599 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X600 end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X601 end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X602 end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X603 end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X604 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X605 end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X606 end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X607 end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X608 end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X609 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X610 end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X611 end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X612 end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X613 end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X614 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X615 end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X616 end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X617 end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X618 end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X619 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X620 end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X621 end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X622 end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X623 end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X624 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X625 end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X626 end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X627 end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X628 end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X629 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X630 end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X631 end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X632 end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X633 end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X634 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X635 end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X636 end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X637 end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X638 end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X639 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X640 mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X641 mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X642 mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X643 mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X644 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X645 mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X646 mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X647 mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X648 mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X649 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X650 mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X651 mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X652 mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X653 mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X654 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X655 mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X656 mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X657 mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X658 mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X659 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X660 mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X661 mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X662 mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X663 mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X664 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X665 mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X666 mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X667 mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X668 mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X669 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X670 mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X671 mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X672 mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X673 mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X674 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X675 mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X676 mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X677 mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X678 mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X679 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X680 mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X681 mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X682 mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X683 mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X684 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X685 mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X686 mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X687 mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X688 mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X689 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X690 mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X691 mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X692 mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X693 mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X694 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X695 mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X696 mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X697 mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X698 mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X699 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X700 mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X701 mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X702 mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X703 mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X704 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X705 mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X706 mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X707 mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X708 mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X709 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X710 mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X711 mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X712 mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X713 mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X714 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X715 mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X716 mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X717 mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X718 mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X719 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X720 end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X721 end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X722 end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X723 end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X724 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X725 end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X726 end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X727 end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X728 end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X729 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X730 end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X731 end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X732 end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X733 end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X734 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X735 end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X736 end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X737 end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X738 end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X739 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X740 end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X741 end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X742 end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X743 end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X744 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X745 end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X746 end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X747 end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X748 end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X749 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X750 end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X751 end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X752 end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X753 end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X754 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X755 end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X756 end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X757 end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X758 end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X759 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X760 end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X761 end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X762 end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X763 end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X764 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X765 end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X766 end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X767 end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X768 end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X769 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X770 end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X771 end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X772 end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X773 end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X774 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X775 end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X776 end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X777 end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X778 end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X779 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X780 end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X781 end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X782 end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X783 end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X784 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X785 end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X786 end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X787 end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X788 end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X789 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X790 end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X791 end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X792 end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X793 end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X794 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X795 end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X796 end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X797 end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X798 end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X799 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X800 mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X801 mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X802 mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X803 mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X804 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X805 mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X806 mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X807 mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X808 mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X809 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X810 mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X811 mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X812 mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X813 mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X814 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X815 mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X816 mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X817 mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X818 mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X819 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X820 mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X821 mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X822 mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X823 mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X824 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X825 mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X826 mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X827 mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X828 mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X829 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X830 mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X831 mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X832 mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X833 mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X834 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X835 mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X836 mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X837 mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X838 mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X839 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X840 mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X841 mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X842 mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X843 mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X844 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X845 mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X846 mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X847 mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X848 mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X849 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X850 mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X851 mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X852 mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X853 mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X854 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X855 mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X856 mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X857 mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X858 mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X859 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X860 mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X861 mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X862 mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X863 mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X864 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X865 mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X866 mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X867 mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X868 mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X869 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X870 mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X871 mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X872 mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X873 mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X874 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X875 mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X876 mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X877 mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X878 mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X879 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X880 end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X881 end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X882 end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X883 end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X884 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X885 end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X886 end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X887 end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X888 end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X889 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X890 end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X891 end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X892 end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X893 end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X894 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X895 end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X896 end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X897 end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X898 end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X899 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X900 end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X901 end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X902 end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X903 end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X904 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X905 end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X906 end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X907 end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X908 end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X909 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X910 end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X911 end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X912 end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X913 end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X914 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X915 end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X916 end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X917 end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X918 end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X919 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X920 end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X921 end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X922 end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X923 end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X924 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X925 end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X926 end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X927 end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X928 end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X929 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X930 end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X931 end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X932 end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X933 end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X934 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X935 end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X936 end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X937 end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X938 end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X939 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X940 end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X941 end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X942 end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X943 end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X944 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X945 end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X946 end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X947 end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X948 end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X949 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X950 end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X951 end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X952 end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X953 end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X954 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X955 end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X956 end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X957 end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X958 end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X959 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X960 end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X961 end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X962 end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X963 end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X964 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X965 end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X966 end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X967 end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X968 end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X969 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X970 end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X971 end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X972 end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X973 end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X974 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X975 end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X976 end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X977 end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X978 end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X979 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X980 end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X981 end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X982 end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X983 end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X984 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X985 end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X986 end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X987 end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X988 end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X989 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X990 end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X991 end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X992 end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X993 end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X994 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X995 end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X996 end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X997 end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X998 end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X999 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1000 end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1001 end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1002 end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1003 end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1004 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1005 end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1006 end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1007 end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1008 end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1009 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1010 end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1011 end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1012 end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1013 end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1014 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1015 end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1016 end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1017 end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1018 end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1019 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1020 end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1021 end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1022 end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1023 end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1024 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1025 end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1026 end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1027 end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1028 end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1029 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1030 end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1031 end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1032 end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1033 end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1034 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1035 end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1036 end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1037 end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1038 end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1039 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1040 mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1041 mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1042 mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1043 mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1044 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1045 mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1046 mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1047 mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1048 mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1049 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1050 mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1051 mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1052 mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1053 mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1054 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1055 mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1056 mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1057 mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1058 mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1059 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1060 mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1061 mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1062 mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1063 mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1064 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1065 mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1066 mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1067 mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1068 mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1069 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1070 mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1071 mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1072 mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1073 mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1074 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1075 mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1076 mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1077 mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1078 mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1079 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1080 mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1081 mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1082 mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1083 mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1084 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1085 mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1086 mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1087 mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1088 mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1089 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1090 mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1091 mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1092 mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1093 mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1094 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1095 mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1096 mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1097 mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1098 mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1099 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1100 mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1101 mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1102 mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1103 mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1104 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1105 mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1106 mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1107 mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1108 mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1109 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1110 mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1111 mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1112 mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1113 mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1114 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1115 mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1116 mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1117 mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1118 mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1119 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1120 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1121 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1122 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1123 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1124 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1125 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1126 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1127 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1128 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1129 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1130 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1131 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1132 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1133 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1134 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1135 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1136 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1137 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1138 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1139 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1140 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1141 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1142 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1143 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1144 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1145 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1146 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1147 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1148 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1149 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1150 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1151 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1152 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1153 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1154 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1155 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1156 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1157 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1158 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1159 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1160 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1161 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1162 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1163 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1164 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1165 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1166 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1167 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1168 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1169 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1170 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1171 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1172 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1173 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1174 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1175 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1176 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1177 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1178 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1179 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1180 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1181 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1182 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1183 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1184 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1185 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1186 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1187 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1188 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1189 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1190 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1191 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1192 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1193 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1194 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1195 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1196 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1197 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1198 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1199 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1200 mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_0/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1201 mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_0/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1202 mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_0/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1203 mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_0/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1204 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1205 mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1206 mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1207 mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1208 mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1209 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1210 mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1211 mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1212 mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1213 mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1214 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1215 mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1216 mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1217 mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1218 mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1219 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1220 mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1221 mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1222 mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1223 mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1224 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1225 mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1226 mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1227 mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1228 mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1229 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1230 mid_2_0/m4_2410_n9430# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1231 mid_2_0/m4_2410_n9430# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1232 mid_2_0/m4_2410_n9430# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1233 mid_2_0/m4_2410_n9430# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1234 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/m4_2410_n9430# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1235 mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1236 mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1237 mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1238 mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1239 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1240 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1241 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1242 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1243 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1244 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1245 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1246 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1247 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1248 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1249 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1250 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1251 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1252 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1253 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_2/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1254 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1255 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1256 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1257 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1258 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1259 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1260 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1261 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1262 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1263 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1264 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1265 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1266 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1267 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1268 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1269 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1270 mid_2_0/mid_2_low_0/m4_2410_n9430# mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1271 mid_2_0/mid_2_low_0/m4_2410_n9430# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1272 mid_2_0/mid_2_low_0/m4_2410_n9430# mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1273 mid_2_0/mid_2_low_0/m4_2410_n9430# mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1274 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/m4_2410_n9430# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1275 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1276 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X1277 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/Vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1278 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1279 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
C0 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# 5.002839f
C1 mid_2_0/8_cap_array_final_0/cap_final_3/phi2 mid_2_0/8_cap_array_final_0/cap_final_2/phi1 2.68972f
C2 mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vdd 4.686877f
C3 mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C4 end_3/8_cap_array_final_1/cap_final_7/Vdd mid_2_0/8_cap_array_final_0/cap_final_0/phi1 37.061146f
C5 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# 5.002838f
C6 mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n 42.41612f
C7 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# 5.002838f
C8 mid_4to8_1/8_cap_array_final_1/m1_n130_1750# mid_4to8_1/8_cap_array_final_1/m1_n130_1630# 8.59886f
C9 mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C10 mid_2_0/8_cap_array_final_0/cap_final_0/phi1_n mid_2_0/8_cap_array_final_0/cap_final_0/phi2_n 25.578663f
C11 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# 5.002494f
C12 mid_6to8_1/8_cap_array_final_1/m1_n130_3980# mid_6to8_1/8_cap_array_final_1/m1_n130_4100# 8.59886f
C13 end_0/8_cap_array_final_1/m1_n130_1870# end_0/8_cap_array_final_1/m1_n130_1750# 8.59886f
C14 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# 5.002838f
C15 mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n mid_2_0/8_cap_array_final_0/cap_final_6/phi1 4.235847f
C16 mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C17 mid_4to8_0/8_cap_array_final_1/m1_n130_1750# mid_4to8_0/8_cap_array_final_1/m1_n130_1630# 8.59886f
C18 mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C19 mid_2to4__1/8_cap_array_final_1/m1_n130_1630# mid_2_0/8_cap_array_final_0/cap_final_2/phi2 8.62096f
C20 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# 5.002838f
C21 mid_4to8_0/8_cap_array_final_1/m1_n130_4340# mid_4to8_0/8_cap_array_final_1/m1_n130_4220# 8.59886f
C22 mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C23 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# 5.002838f
C24 mid_6to8_3/8_cap_array_final_1/m1_n130_3980# mid_6to8_3/8_cap_array_final_1/m1_n130_4100# 8.59886f
C25 end_3/8_cap_array_final_1/m1_n130_1870# end_3/8_cap_array_final_1/m1_n130_1750# 8.59886f
C26 end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/phi1 2.178203f
C27 mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C28 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# 5.002839f
C29 mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C30 mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C31 mid_6to8_0/8_cap_array_final_1/m1_n130_4340# mid_6to8_0/8_cap_array_final_1/m1_n130_4220# 8.59886f
C32 mid_2_0/8_cap_array_final_0/cap_final_6/phi2 mid_2_0/8_cap_array_final_0/cap_final_6/phi1 83.12768f
C33 mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin 4.006585f
C34 mid_2_0/8_cap_array_final_0/cap_final_4/phi2 mid_2_0/8_cap_array_final_0/cap_final_6/phi1 39.084137f
C35 mid_2_0/8_cap_array_final_0/cap_final_6/phi2 mid_6to8_2/8_cap_array_final_1/m1_n130_2110# 8.66467f
C36 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# 5.272134f
C37 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi2_n mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi1_n 25.456757f
C38 mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/Vin 3.020648f
C39 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# 5.002838f
C40 mid_6to8_1/8_cap_array_final_1/m1_n130_2110# mid_6to8_1/8_cap_array_final_1/m1_n130_1990# 8.59886f
C41 mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C42 mid_2_0/8_cap_array_final_0/cap_final_3/phi1 mid_2_0/8_cap_array_final_0/cap_final_2/phi2 37.594597f
C43 mid_2_0/8_cap_array_final_0/cap_final_3/phi1 mid_2_0/8_cap_array_final_0/cap_final_6/phi2 6.085594f
C44 mid_2_0/8_cap_array_final_0/cap_final_3/phi1 mid_2_0/8_cap_array_final_0/cap_final_4/phi2 6.49583f
C45 mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C46 mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C47 mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C48 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# 5.002839f
C49 mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C50 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# 4.979833f
C51 mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vdd 18.423512f
C52 end_0/8_cap_array_final_1/m1_n130_1750# end_0/8_cap_array_final_1/m1_n130_1630# 8.59886f
C53 mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C54 mid_4to8_3/8_cap_array_final_1/m1_n130_4340# mid_4to8_3/8_cap_array_final_1/m1_n130_4220# 8.59886f
C55 mid_6to8_3/8_cap_array_final_1/m1_n130_2110# mid_6to8_3/8_cap_array_final_1/m1_n130_1990# 8.59886f
C56 mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n 36.905354f
C57 mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C58 mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n 7.061357f
C59 end_3/8_cap_array_final_1/cap_final_7/Vdd end_3/8_cap_array_final_1/cap_final_7/phi2_n 33.527004f
C60 mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C61 end_2/8_cap_array_final_1/m1_n130_4340# end_2/8_cap_array_final_1/m1_n130_4220# 8.59886f
C62 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# 5.002838f
C63 mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C64 mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n mid_6to8_2/8_cap_array_final_1/m1_n130_3980# 8.664217f
C65 mid_6to8_1/8_cap_array_final_1/m1_n130_4220# mid_6to8_1/8_cap_array_final_1/m1_n130_4100# 8.59886f
C66 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# 5.002838f
C67 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# 5.002839f
C68 mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/phi2_n 21.364698f
C69 mid_4to8_0/8_cap_array_final_1/m1_n130_4460# mid_4to8_0/8_cap_array_final_1/m1_n130_4340# 8.59886f
C70 end_3/8_cap_array_final_1/m1_n130_1750# end_3/8_cap_array_final_1/m1_n130_1630# 8.59886f
C71 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# 5.002839f
C72 end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/GND 5.607867f
C73 mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n 38.046253f
C74 mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C75 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1_n mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2_n 29.46952f
C76 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1_n mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1 2.693218f
C77 mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C78 mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n 18.272886f
C79 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# 5.002839f
C80 mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C81 mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C82 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# 5.002838f
C83 mid_6to8_3/8_cap_array_final_1/m1_n130_4220# mid_6to8_3/8_cap_array_final_1/m1_n130_4100# 8.59886f
C84 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2 mid_2_0/8_cap_array_final_0/cap_final_2/phi1 39.219715f
C85 mid_2_0/8_cap_array_final_0/cap_final_3/phi1 mid_2_0/8_cap_array_final_0/cap_final_3/phi2 64.9875f
C86 end_3/8_cap_array_final_1/cap_final_7/Vdd end_3/8_cap_array_final_1/cap_final_7/Vin 48.838326f
C87 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# 5.002839f
C88 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# 5.002493f
C89 mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C90 mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n 55.251537f
C91 mid_6to8_1/8_cap_array_final_1/m1_n130_1990# mid_6to8_1/8_cap_array_final_1/m1_n130_1870# 8.59886f
C92 mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin 16.566456f
C93 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi1 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi2 40.405228f
C94 mid_2_0/8_cap_array_final_0/cap_final_4/phi1 mid_2_0/8_cap_array_final_0/cap_final_6/phi1 42.98026f
C95 end_0/8_cap_array_final_1/m1_n130_4460# end_0/8_cap_array_final_1/m1_n130_4340# 8.59886f
C96 end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/cap_final_7/Vin 0.246419p
C97 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# 5.272134f
C98 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# 5.002839f
C99 mid_2_0/8_cap_array_final_0/cap_final_4/phi2 mid_2_0/8_cap_array_final_0/cap_final_6/phi2 36.94984f
C100 mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272134f
C101 mid_6to8_3/8_cap_array_final_1/m1_n130_1990# mid_6to8_3/8_cap_array_final_1/m1_n130_1870# 8.59886f
C102 end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C103 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2_n mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2 2.730069f
C104 mid_2to4__0/8_cap_array_final_1/m1_n130_1630# mid_2_0/8_cap_array_final_0/cap_final_2/phi2 8.62096f
C105 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# 5.002839f
C106 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi2 37.759907f
C107 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# 5.272134f
C108 mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C109 mid_2_0/8_cap_array_final_0/cap_final_3/phi1 mid_2_0/8_cap_array_final_0/cap_final_4/phi1 84.24828f
C110 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# 4.980177f
C111 end_3/8_cap_array_final_1/m1_n130_4460# end_3/8_cap_array_final_1/m1_n130_4340# 8.59886f
C112 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# 4.980177f
C113 mid_2_0/8_cap_array_final_0/cap_final_6/phi1 end_3/8_cap_array_final_1/cap_final_7/phi1 0.130666p
C114 mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C115 mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C116 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# 5.002839f
C117 mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C118 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# 5.002838f
C119 mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n mid_4to8_1/8_cap_array_final_1/m1_n130_4220# 8.649531f
C120 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# 5.002839f
C121 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1_n mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2_n 21.9877f
C122 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# 5.002493f
C123 end_3/8_cap_array_final_1/cap_final_7/phi2_n end_0/8_cap_array_final_1/m1_n130_3860# 8.72684f
C124 mid_2_0/8_cap_array_final_0/cap_final_3/phi1 end_3/8_cap_array_final_1/cap_final_7/phi1 2.300412f
C125 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# 5.002838f
C126 mid_2_0/8_cap_array_final_0/cap_final_2/phi2 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2 9.110595f
C127 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# 5.002838f
C128 mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C129 mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C130 mid_6to8_1/8_cap_array_final_1/m1_n130_1870# mid_6to8_1/8_cap_array_final_1/m1_n130_1750# 8.59886f
C131 mid_4to8_1/8_cap_array_final_1/m1_n130_4340# mid_4to8_1/8_cap_array_final_1/m1_n130_4460# 8.59886f
C132 mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C133 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# 5.002838f
C134 mid_2_0/8_cap_array_final_0/cap_final_3/phi2 mid_2_0/8_cap_array_final_0/cap_final_2/phi2 18.284271f
C135 mid_2_0/8_cap_array_final_0/cap_final_0/phi2_n mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2_n 9.007117f
C136 mid_2_0/8_cap_array_final_0/cap_final_3/phi2 mid_2_0/8_cap_array_final_0/cap_final_6/phi2 36.360214f
C137 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# 5.002838f
C138 mid_2_0/8_cap_array_final_0/cap_final_4/phi2 mid_2_0/8_cap_array_final_0/cap_final_3/phi2 72.199745f
C139 end_1/8_cap_array_final_1/m1_n130_2230# end_1/8_cap_array_final_1/m1_n130_2110# 8.59886f
C140 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2_n mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n 17.995602f
C141 mid_4to8_2/8_cap_array_final_1/m1_n130_1870# mid_4to8_2/8_cap_array_final_1/m1_n130_1750# 8.59886f
C142 mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C143 mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C144 end_3/8_cap_array_final_1/cap_final_7/phi1_n mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n 28.056658f
C145 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1_n mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi1_n 8.918006f
C146 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# 5.002839f
C147 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# 5.002838f
C148 mid_2_0/8_cap_array_final_0/cap_final_4/phi2 mid_4to8_3/8_cap_array_final_1/m1_n130_1870# 8.649647f
C149 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# 5.002839f
C150 mid_6to8_3/8_cap_array_final_1/m1_n130_1870# mid_6to8_3/8_cap_array_final_1/m1_n130_1750# 8.59886f
C151 mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C152 end_1/8_cap_array_final_1/m1_n130_3980# end_1/8_cap_array_final_1/m1_n130_4100# 8.59886f
C153 mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C154 mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C155 end_3/8_cap_array_final_1/cap_final_7/Vdd end_3/8_cap_array_final_1/cap_final_7/phi1 4.889181f
C156 end_3/8_cap_array_final_1/cap_final_7/phi2 mid_2_0/8_cap_array_final_0/cap_final_6/phi1 21.651308f
C157 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# 5.002839f
C158 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1_n mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n 9.312764f
C159 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi1 8.931144f
C160 mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C161 mid_2_0/8_cap_array_final_0/cap_final_4/phi1 mid_2_0/8_cap_array_final_0/cap_final_6/phi2 7.159061f
C162 mid_2_0/8_cap_array_final_0/cap_final_4/phi1 mid_2_0/8_cap_array_final_0/cap_final_4/phi2 69.67373f
C163 mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C164 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1 mid_2_0/8_cap_array_final_0/cap_final_2/phi1 18.34155f
C165 mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272135f
C166 mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C167 mid_2_0/8_cap_array_final_0/cap_final_0/phi2_n mid_2_0/8_cap_array_final_0/cap_final_0/phi2 2.638682f
C168 mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/phi1_n 2.907911f
C169 end_0/8_cap_array_final_1/m1_n130_4340# end_0/8_cap_array_final_1/m1_n130_4220# 8.59886f
C170 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# 5.002839f
C171 mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C172 mid_6to8_1/8_cap_array_final_1/m1_n130_1750# mid_6to8_1/8_cap_array_final_1/m1_n130_1630# 8.59886f
C173 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# 5.002839f
C174 mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n 22.605503f
C175 mid_2_0/8_cap_array_final_0/cap_final_4/phi2 mid_4to8_0/8_cap_array_final_1/m1_n130_1870# 8.649647f
C176 mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/phi1 43.301292f
C177 end_1/8_cap_array_final_1/m1_n130_2110# end_1/8_cap_array_final_1/m1_n130_1990# 8.59886f
C178 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# 5.002838f
C179 mid_4to8_2/8_cap_array_final_1/m1_n130_1750# mid_4to8_2/8_cap_array_final_1/m1_n130_1630# 8.59886f
C180 end_3/8_cap_array_final_1/m1_n130_4340# end_3/8_cap_array_final_1/m1_n130_4220# 8.59886f
C181 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# 5.002838f
C182 end_3/8_cap_array_final_1/cap_final_7/Vin end_3/8_cap_array_final_1/cap_final_7/phi1 6.758001f
C183 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# 5.002839f
C184 mid_6to8_3/8_cap_array_final_1/m1_n130_1750# mid_6to8_3/8_cap_array_final_1/m1_n130_1630# 8.59886f
C185 mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C186 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# 5.002838f
C187 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi1 mid_2_0/8_cap_array_final_0/cap_final_0/phi2 36.920002f
C188 mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C189 mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n 36.33864f
C190 mid_2_0/8_cap_array_final_0/cap_final_4/phi1 mid_2_0/8_cap_array_final_0/cap_final_3/phi2 43.597073f
C191 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# 5.002838f
C192 end_1/8_cap_array_final_1/m1_n130_3980# end_1/8_cap_array_final_1/m1_n130_3860# 8.59886f
C193 end_1/8_cap_array_final_1/m1_n130_4220# end_1/8_cap_array_final_1/m1_n130_4100# 8.59886f
C194 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# 5.002838f
C195 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi1_n mid_2_0/8_cap_array_final_0/cap_final_0/phi2_n 21.9664f
C196 end_3/8_cap_array_final_1/cap_final_7/phi2 end_2/8_cap_array_final_1/m1_n130_2230# 8.728628f
C197 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1_n mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n 18.339928f
C198 mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C199 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# 5.002839f
C200 mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1_n 2.193301f
C201 mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C202 mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n mid_4to8_3/8_cap_array_final_1/m1_n130_4220# 8.649531f
C203 end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/phi2_n 5.805031f
C204 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# 5.002839f
C205 mid_6to8_1/8_cap_array_final_1/m1_n130_4460# mid_6to8_1/8_cap_array_final_1/m1_n130_4340# 8.59886f
C206 mid_2_0/8_cap_array_final_0/cap_final_6/phi2 mid_6to8_1/8_cap_array_final_1/m1_n130_2110# 8.66467f
C207 mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n 72.16842f
C208 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2 mid_2_0/8_cap_array_final_0/cap_final_2/phi2 18.01004f
C209 mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n 28.517117f
C210 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# 5.002838f
C211 mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND 13.09726f
C212 end_1/8_cap_array_final_1/m1_n130_1990# end_1/8_cap_array_final_1/m1_n130_1870# 8.59886f
C213 end_3/8_cap_array_final_1/cap_final_7/phi2 mid_2_0/8_cap_array_final_0/cap_final_6/phi2 0.108955p
C214 mid_4to8_2/8_cap_array_final_1/m1_n130_4460# mid_4to8_2/8_cap_array_final_1/m1_n130_4340# 8.59886f
C215 mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C216 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# 5.002839f
C217 mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C218 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# 4.980177f
C219 end_3/8_cap_array_final_1/cap_final_7/Vdd mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n 2.116855f
C220 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi1_n mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi1 2.605365f
C221 mid_6to8_3/8_cap_array_final_1/m1_n130_4460# mid_6to8_3/8_cap_array_final_1/m1_n130_4340# 8.59886f
C222 mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C223 mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C224 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# 4.980177f
C225 mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C226 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# 5.002838f
C227 mid_2_0/8_cap_array_final_0/cap_final_4/phi1 end_3/8_cap_array_final_1/cap_final_7/phi1 3.002692f
C228 mid_2_0/8_cap_array_final_0/cap_final_0/phi1_n mid_2_0/8_cap_array_final_0/cap_final_0/phi1 2.612484f
C229 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# 5.002838f
C230 mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C231 mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n mid_6to8_1/8_cap_array_final_1/m1_n130_3980# 8.664217f
C232 mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND 6.603709f
C233 mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C234 mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C235 mid_2_0/8_cap_array_final_0/cap_final_3/phi1 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1 19.728592f
C236 mid_2_0/8_cap_array_final_0/cap_final_2/phi2 mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n 3.017917f
C237 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# 5.002839f
C238 mid_2_0/8_cap_array_final_0/cap_final_3/phi2 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2 18.108353f
C239 mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C240 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# 5.002838f
C241 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# 5.002838f
C242 mid_2_0/8_cap_array_final_0/cap_final_4/phi2 mid_4to8_2/8_cap_array_final_1/m1_n130_1870# 8.649647f
C243 end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/m1_n130_2230# 8.728628f
C244 mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C245 mid_6to8_2/8_cap_array_final_1/m1_n130_3980# mid_6to8_2/8_cap_array_final_1/m1_n130_4100# 8.59886f
C246 end_1/8_cap_array_final_1/m1_n130_1870# end_1/8_cap_array_final_1/m1_n130_1750# 8.59886f
C247 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1_n mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2_n 29.427896f
C248 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# 5.002839f
C249 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# 4.980177f
C250 mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272134f
C251 mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272134f
C252 end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C253 mid_6to8_1/8_cap_array_final_1/m1_n130_4340# mid_6to8_1/8_cap_array_final_1/m1_n130_4220# 8.59886f
C254 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# 5.002839f
C255 mid_2_0/8_cap_array_final_0/cap_final_2/phi1 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi1 9.170131f
C256 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# 5.002838f
C257 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# 5.272133f
C258 mid_4to8_2/8_cap_array_final_1/m1_n130_4340# mid_4to8_2/8_cap_array_final_1/m1_n130_4220# 8.59886f
C259 mid_6to8_2/8_cap_array_final_1/m1_n130_2110# mid_6to8_2/8_cap_array_final_1/m1_n130_1990# 8.59886f
C260 mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n 6.004341f
C261 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# 5.002838f
C262 mid_6to8_3/8_cap_array_final_1/m1_n130_4340# mid_6to8_3/8_cap_array_final_1/m1_n130_4220# 8.59886f
C263 end_3/8_cap_array_final_1/cap_final_7/phi2 end_3/8_cap_array_final_1/cap_final_7/phi1 96.23077f
C264 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# 5.002839f
C265 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1 mid_2_0/8_cap_array_final_0/cap_final_2/phi1 9.289417f
C266 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/m4_2410_n9430# 5.002839f
C267 mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C268 mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C269 mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C270 end_1/8_cap_array_final_1/m1_n130_1750# end_1/8_cap_array_final_1/m1_n130_1630# 8.59886f
C271 mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1_n 19.731527f
C272 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# 5.002838f
C273 mid_6to8_2/8_cap_array_final_1/m1_n130_4220# mid_6to8_2/8_cap_array_final_1/m1_n130_4100# 8.59886f
C274 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# 5.002838f
C275 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# 5.002838f
C276 mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C277 mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n 6.385192f
C278 end_3/8_cap_array_final_1/cap_final_7/Vin mid_2_0/8_cap_array_final_0/cap_final_0/phi1_n 22.264221f
C279 mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n 84.23691f
C280 end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/GND 12.56054f
C281 mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C282 mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi1_n 9.193998f
C283 mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n mid_4to8_2/8_cap_array_final_1/m1_n130_4220# 8.649531f
C284 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2 36.950897f
C285 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# 5.002838f
C286 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# 5.002839f
C287 mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C288 mid_2_0/8_cap_array_final_0/cap_final_3/phi2 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1 2.222702f
C289 mid_6to8_2/8_cap_array_final_1/m1_n130_1990# mid_6to8_2/8_cap_array_final_1/m1_n130_1870# 8.59886f
C290 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# 5.002838f
C291 end_3/8_cap_array_final_1/cap_final_7/Vdd mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n 16.618898f
C292 mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C293 mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n 2.654304f
C294 end_1/8_cap_array_final_1/m1_n130_4460# end_1/8_cap_array_final_1/m1_n130_4340# 8.59886f
C295 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# 5.27179f
C296 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# 5.002839f
C297 mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C298 mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n 69.256165f
C299 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# 5.002838f
C300 mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C301 mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/phi2_n 0.108858p
C302 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# 5.002839f
C303 mid_6to8_0/8_cap_array_final_1/m1_n130_3980# mid_6to8_0/8_cap_array_final_1/m1_n130_4100# 8.59886f
C304 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1 mid_2_0/8_cap_array_final_0/cap_final_0/phi1 8.929021f
C305 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# 5.002839f
C306 mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C307 mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C308 mid_2_0/8_cap_array_final_0/cap_final_2/phi2 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi2 9.05189f
C309 mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n end_3/8_cap_array_final_1/cap_final_7/Vdd 8.281558f
C310 mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vdd 8.691263f
C311 mid_2_0/8_cap_array_final_0/cap_final_6/phi2 mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n 4.41127f
C312 mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n 24.055714f
C313 end_3/8_cap_array_final_1/cap_final_7/phi2_n end_2/8_cap_array_final_1/m1_n130_3860# 8.72684f
C314 mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n 42.957775f
C315 mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/GND 3.442492f
C316 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# 5.002493f
C317 mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n end_3/8_cap_array_final_1/cap_final_7/Vin 2.262305f
C318 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# 5.002838f
C319 end_3/8_cap_array_final_1/cap_final_7/phi2 end_1/8_cap_array_final_1/m1_n130_2230# 8.728628f
C320 mid_6to8_2/8_cap_array_final_1/m1_n130_1870# mid_6to8_2/8_cap_array_final_1/m1_n130_1750# 8.59886f
C321 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# 5.002838f
C322 mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C323 mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C324 mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n mid_2_0/8_cap_array_final_0/cap_final_2/phi1 2.93221f
C325 end_2/8_cap_array_final_1/m1_n130_2230# end_2/8_cap_array_final_1/m1_n130_2110# 8.59886f
C326 mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C327 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# 5.002839f
C328 mid_2_0/8_cap_array_final_0/cap_final_6/phi2 mid_6to8_0/8_cap_array_final_1/m1_n130_2110# 8.66467f
C329 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi2_n mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n 9.046399f
C330 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# 5.002494f
C331 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# 5.002494f
C332 mid_2_0/8_cap_array_final_0/cap_final_4/phi2 mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n 3.66953f
C333 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# 5.002838f
C334 mid_2_0/8_cap_array_final_0/cap_final_0/phi1 mid_2_0/8_cap_array_final_0/cap_final_0/phi2 40.528915f
C335 end_2/8_cap_array_final_1/m1_n130_3980# end_2/8_cap_array_final_1/m1_n130_4100# 8.59886f
C336 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi2 8.979368f
C337 mid_6to8_0/8_cap_array_final_1/m1_n130_2110# mid_6to8_0/8_cap_array_final_1/m1_n130_1990# 8.59886f
C338 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C339 mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C340 mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n end_3/8_cap_array_final_1/cap_final_7/phi1_n 2.231639f
C341 mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C342 mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin 7.361336f
C343 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# 4.980177f
C344 mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C345 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# 4.980177f
C346 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# 5.272134f
C347 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2_n mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n 24.224424f
C348 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# 5.002494f
C349 mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2_n 18.107841f
C350 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# 5.002839f
C351 mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C352 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# 5.002839f
C353 end_1/8_cap_array_final_1/m1_n130_4340# end_1/8_cap_array_final_1/m1_n130_4220# 8.59886f
C354 mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C355 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2 44.305923f
C356 mid_6to8_0/8_cap_array_final_1/m1_n130_4220# mid_6to8_0/8_cap_array_final_1/m1_n130_4100# 8.59886f
C357 mid_6to8_0/8_cap_array_final_1/m1_n130_3980# mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n 8.664217f
C358 mid_6to8_2/8_cap_array_final_1/m1_n130_1750# mid_6to8_2/8_cap_array_final_1/m1_n130_1630# 8.59886f
C359 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# 5.002494f
C360 mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272134f
C361 mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C362 mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C363 end_2/8_cap_array_final_1/m1_n130_2110# end_2/8_cap_array_final_1/m1_n130_1990# 8.59886f
C364 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# 5.002838f
C365 end_3/8_cap_array_final_1/cap_final_7/phi2_n end_3/8_cap_array_final_1/m1_n130_3860# 8.72684f
C366 mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C367 mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272134f
C368 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# 5.002838f
C369 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# 5.002838f
C370 mid_2to4__1/8_cap_array_final_1/m1_n130_4460# mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n 8.620945f
C371 mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C372 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# 5.002493f
C373 mid_6to8_0/8_cap_array_final_1/m1_n130_1990# mid_6to8_0/8_cap_array_final_1/m1_n130_1870# 8.59886f
C374 mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C375 mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n 20.080708f
C376 end_3/8_cap_array_final_1/cap_final_7/Vdd end_3/8_cap_array_final_1/cap_final_7/phi1_n 51.499012f
C377 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# 5.002838f
C378 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# 5.002839f
C379 end_2/8_cap_array_final_1/m1_n130_3980# end_2/8_cap_array_final_1/m1_n130_3860# 8.59886f
C380 end_2/8_cap_array_final_1/m1_n130_4220# end_2/8_cap_array_final_1/m1_n130_4100# 8.59886f
C381 mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n 50.32686f
C382 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# 5.002839f
C383 mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C384 mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/phi1_n 0.130461p
C385 mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C386 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# 5.002839f
C387 mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n mid_2_0/8_cap_array_final_0/cap_final_4/phi1 3.570629f
C388 end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/phi2_n 83.35017f
C389 mid_6to8_2/8_cap_array_final_1/m1_n130_4460# mid_6to8_2/8_cap_array_final_1/m1_n130_4340# 8.59886f
C390 mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C391 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2_n 2.752844f
C392 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2 44.41014f
C393 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# 5.272134f
C394 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# 5.002839f
C395 mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C396 mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C397 mid_4to8_1/8_cap_array_final_1/m1_n130_4340# mid_4to8_1/8_cap_array_final_1/m1_n130_4220# 8.59886f
C398 end_2/8_cap_array_final_1/m1_n130_1990# end_2/8_cap_array_final_1/m1_n130_1870# 8.59886f
C399 mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C400 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# 5.002838f
C401 mid_4to8_1/8_cap_array_final_1/m1_n130_1870# mid_2_0/8_cap_array_final_0/cap_final_4/phi2 8.649647f
C402 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# 5.002494f
C403 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1_n mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi2_n 22.7839f
C404 end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/Vin 46.440384f
C405 mid_6to8_0/8_cap_array_final_1/m1_n130_1870# mid_6to8_0/8_cap_array_final_1/m1_n130_1750# 8.59886f
C406 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# 5.002839f
C407 mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C408 mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C409 end_0/8_cap_array_final_1/m1_n130_2230# end_0/8_cap_array_final_1/m1_n130_2110# 8.59886f
C410 mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C411 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# 5.002494f
C412 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# 5.002838f
C413 mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n mid_4to8_0/8_cap_array_final_1/m1_n130_4220# 8.649531f
C414 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# 5.002838f
C415 end_3/8_cap_array_final_1/cap_final_7/Vdd end_3/8_cap_array_final_1/cap_final_7/com_x 2.626611f
C416 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2 mid_2_0/8_cap_array_final_0/cap_final_0/phi2 9.010565f
C417 end_3/8_cap_array_final_1/cap_final_7/Vdd mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n 2.178562f
C418 end_0/8_cap_array_final_1/m1_n130_3980# end_0/8_cap_array_final_1/m1_n130_4100# 8.59886f
C419 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# 5.002838f
C420 mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C421 mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n end_3/8_cap_array_final_1/cap_final_7/Vdd 4.265811f
C422 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# 5.002494f
C423 end_3/8_cap_array_final_1/m1_n130_2230# end_3/8_cap_array_final_1/m1_n130_2110# 8.59886f
C424 mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C425 mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C426 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi2_n mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi2 2.615672f
C427 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# 5.002493f
C428 mid_4to8_3/8_cap_array_final_1/m1_n130_1870# mid_4to8_3/8_cap_array_final_1/m1_n130_1750# 8.59886f
C429 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# 5.002838f
C430 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# 5.002838f
C431 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# 5.002839f
C432 end_3/8_cap_array_final_1/m1_n130_3980# end_3/8_cap_array_final_1/m1_n130_4100# 8.59886f
C433 mid_2_0/8_cap_array_final_0/cap_final_3/phi1 mid_2_0/8_cap_array_final_0/cap_final_2/phi1 20.084393f
C434 end_2/8_cap_array_final_1/m1_n130_1870# end_2/8_cap_array_final_1/m1_n130_1750# 8.59886f
C435 mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C436 mid_2to4__0/8_cap_array_final_1/m1_n130_4460# mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n 8.620945f
C437 mid_2_0/8_cap_array_final_0/cap_final_6/phi2 mid_6to8_3/8_cap_array_final_1/m1_n130_2110# 8.66467f
C438 mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C439 mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C440 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# 5.272134f
C441 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# 5.272133f
C442 mid_6to8_0/8_cap_array_final_1/m1_n130_1750# mid_6to8_0/8_cap_array_final_1/m1_n130_1630# 8.59886f
C443 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# 5.002838f
C444 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# 5.002839f
C445 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# 5.002839f
C446 end_3/8_cap_array_final_1/cap_final_7/Vdd end_3/8_cap_array_final_1/cap_final_7/GND 0.288759p
C447 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# 5.002838f
C448 mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C449 end_3/8_cap_array_final_1/cap_final_7/com_x end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# 5.002839f
C450 mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C451 end_0/8_cap_array_final_1/m1_n130_2110# end_0/8_cap_array_final_1/m1_n130_1990# 8.59886f
C452 mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n end_3/8_cap_array_final_1/cap_final_7/GND 3.445286f
C453 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# 5.002838f
C454 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# 5.002839f
C455 mid_6to8_2/8_cap_array_final_1/m1_n130_4340# mid_6to8_2/8_cap_array_final_1/m1_n130_4220# 8.59886f
C456 mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C457 end_3/8_cap_array_final_1/cap_final_7/com_x end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# 5.002493f
C458 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/m4_2410_n9430# 5.002838f
C459 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# 5.002839f
C460 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# 5.002839f
C461 end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/phi2_n 27.94766f
C462 end_3/8_cap_array_final_1/m1_n130_2110# end_3/8_cap_array_final_1/m1_n130_1990# 8.59886f
C463 mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C464 mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C465 mid_4to8_3/8_cap_array_final_1/m1_n130_1750# mid_4to8_3/8_cap_array_final_1/m1_n130_1630# 8.59886f
C466 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# 5.002838f
C467 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1_n mid_2_0/8_cap_array_final_0/cap_final_0/phi1_n 8.91752f
C468 end_3/8_cap_array_final_1/cap_final_7/phi2_n end_1/8_cap_array_final_1/m1_n130_3860# 8.72684f
C469 end_3/8_cap_array_final_1/cap_final_7/phi1_n end_3/8_cap_array_final_1/cap_final_7/phi1 24.894503f
C470 mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n mid_6to8_3/8_cap_array_final_1/m1_n130_3980# 8.664217f
C471 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# 5.002838f
C472 mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C473 end_0/8_cap_array_final_1/m1_n130_3980# end_0/8_cap_array_final_1/m1_n130_3860# 8.59886f
C474 end_0/8_cap_array_final_1/m1_n130_4220# end_0/8_cap_array_final_1/m1_n130_4100# 8.59886f
C475 mid_2_0/8_cap_array_final_0/cap_final_6/phi2 end_3/8_cap_array_final_1/cap_final_7/GND 2.737761f
C476 end_3/8_cap_array_final_1/cap_final_7/phi2 end_0/8_cap_array_final_1/m1_n130_2230# 8.728628f
C477 end_2/8_cap_array_final_1/m1_n130_1750# end_2/8_cap_array_final_1/m1_n130_1630# 8.59886f
C478 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# 5.002838f
C479 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# 5.002838f
C480 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# 5.002838f
C481 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# 5.002839f
C482 end_3/8_cap_array_final_1/cap_final_7/GND end_3/8_cap_array_final_1/cap_final_7/Vin 0.234498p
C483 mid_2_0/8_cap_array_final_0/cap_final_3/phi2 mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n 3.331975f
C484 mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C485 end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C486 mid_6to8_0/8_cap_array_final_1/m1_n130_4460# mid_6to8_0/8_cap_array_final_1/m1_n130_4340# 8.59886f
C487 mid_2_0/8_cap_array_final_0/cap_final_2/phi2 mid_2_0/8_cap_array_final_0/cap_final_2/phi1 52.873554f
C488 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# 5.002838f
C489 end_3/8_cap_array_final_1/m1_n130_3980# end_3/8_cap_array_final_1/m1_n130_3860# 8.59886f
C490 end_3/8_cap_array_final_1/m1_n130_4220# end_3/8_cap_array_final_1/m1_n130_4100# 8.59886f
C491 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# 5.002839f
C492 mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C493 mid_4to8_1/8_cap_array_final_1/m1_n130_1870# mid_4to8_1/8_cap_array_final_1/m1_n130_1750# 8.59886f
C494 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# 5.002839f
C495 end_3/8_cap_array_final_1/cap_final_7/com_x end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# 5.002838f
C496 mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C497 end_3/8_cap_array_final_1/cap_final_7/com_x mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# 5.002838f
C498 end_0/8_cap_array_final_1/m1_n130_1990# end_0/8_cap_array_final_1/m1_n130_1870# 8.59886f
C499 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi2_n mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2_n 8.973002f
C500 mid_2_0/8_cap_array_final_0/cap_final_3/phi1 mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n 3.266874f
C501 mid_4to8_0/8_cap_array_final_1/m1_n130_1870# mid_4to8_0/8_cap_array_final_1/m1_n130_1750# 8.59886f
C502 end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 4.980177f
C503 mid_2_0/8_cap_array_final_0/cap_final_3/phi1 mid_2_0/8_cap_array_final_0/cap_final_6/phi1 42.41868f
C504 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1_n mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1 2.727184f
C505 mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C506 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# 5.002839f
C507 mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C508 mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C509 mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.272134f
C510 mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002839f
C511 end_3/8_cap_array_final_1/m1_n130_1990# end_3/8_cap_array_final_1/m1_n130_1870# 8.59886f
C512 mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2_n 9.101527f
C513 mid_4to8_3/8_cap_array_final_1/m1_n130_4460# mid_4to8_3/8_cap_array_final_1/m1_n130_4340# 8.59886f
C514 end_3/8_cap_array_final_1/cap_final_7/com_x end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# 5.002839f
C515 end_2/8_cap_array_final_1/m1_n130_4460# end_2/8_cap_array_final_1/m1_n130_4340# 8.59886f
C516 end_3/8_cap_array_final_1/cap_final_7/com_x mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# 5.002838f
C517 mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# end_3/8_cap_array_final_1/cap_final_7/com_x 5.002838f
C518 mid_2_0/8_cap_array_final_0/cap_final_0/phi2 VSUBS 4.148705f
C519 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C520 mid_2_0/mid_2_low_0/m4_2410_n9430# VSUBS 3.134649f **FLOATING
C521 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_5/m1_990_n540# VSUBS 3.34045f **FLOATING
C522 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_4/m1_990_n540# VSUBS 3.34039f **FLOATING
C523 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_3/m1_990_n540# VSUBS 3.340337f **FLOATING
C524 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_2/m1_990_n540# VSUBS 3.340289f **FLOATING
C525 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_1/m1_990_n540# VSUBS 3.33782f **FLOATING
C526 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/m1_990_n540# VSUBS 3.340238f **FLOATING
C527 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2_n VSUBS 19.2161f
C528 mid_2_0/8_cap_array_final_0/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C529 mid_2_0/m4_2410_n9430# VSUBS 3.134649f **FLOATING
C530 mid_2_0/8_cap_array_final_0/cap_final_5/m1_990_n540# VSUBS 3.34045f **FLOATING
C531 mid_2_0/8_cap_array_final_0/cap_final_4/m1_990_n540# VSUBS 3.34039f **FLOATING
C532 mid_2_0/8_cap_array_final_0/cap_final_3/m1_990_n540# VSUBS 3.340337f **FLOATING
C533 mid_2_0/8_cap_array_final_0/cap_final_2/m1_990_n540# VSUBS 3.340289f **FLOATING
C534 mid_2_0/8_cap_array_final_0/cap_final_1/m1_990_n540# VSUBS 3.33782f **FLOATING
C535 mid_2_0/8_cap_array_final_0/cap_final_0/m1_990_n540# VSUBS 3.340237f **FLOATING
C536 mid_2_0/8_cap_array_final_0/cap_final_0/phi1 VSUBS 6.571877f
C537 mid_2_0/8_cap_array_final_0/cap_final_0/phi1_n VSUBS 6.322745f
C538 mid_2_0/8_cap_array_final_0/cap_final_0/phi2_n VSUBS 10.678959f
C539 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_7/m1_990_n540# VSUBS 3.340289f **FLOATING
C540 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_6/m1_990_n540# VSUBS 3.340337f **FLOATING
C541 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_5/m1_990_n540# VSUBS 3.340391f **FLOATING
C542 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_4/m1_990_n540# VSUBS 3.34045f **FLOATING
C543 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_3/m1_990_n540# VSUBS 3.34045f **FLOATING
C544 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C545 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/m1_990_n540# VSUBS 3.340247f **FLOATING
C546 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_1/phi1 VSUBS 2.085098f
C547 mid_2_0/mid_2_up_left_1/8_cap_array_final_1/cap_final_0/m1_990_n540# VSUBS 3.475442f **FLOATING
C548 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi2 VSUBS 7.202928f
C549 mid_2_0/8_cap_array_final_0/cap_final_2/phi2 VSUBS 10.852775f
C550 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_7/m1_990_n540# VSUBS 3.340289f **FLOATING
C551 mid_2_0/8_cap_array_final_0/cap_final_2/phi1 VSUBS 13.563651f
C552 mid_2_0/8_cap_array_final_0/cap_final_2/phi1_n VSUBS 17.198885f
C553 mid_2_0/8_cap_array_final_0/cap_final_2/phi2_n VSUBS 17.720972f
C554 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_6/m1_990_n540# VSUBS 3.340337f **FLOATING
C555 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_5/m1_990_n540# VSUBS 3.340391f **FLOATING
C556 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_4/m1_990_n540# VSUBS 3.34045f **FLOATING
C557 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_3/m1_990_n540# VSUBS 3.34045f **FLOATING
C558 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C559 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_1/m1_990_n540# VSUBS 3.340247f **FLOATING
C560 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1 VSUBS 10.206014f
C561 mid_2_0/mid_2_low_0/8_cap_array_final_0/cap_final_0/phi1_n VSUBS 14.554255f
C562 mid_2_0/mid_2_up_left_0/8_cap_array_final_1/cap_final_0/m1_990_n540# VSUBS 3.475442f **FLOATING
C563 mid_6to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C564 mid_6to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# VSUBS 3.340515f **FLOATING
C565 mid_6to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# VSUBS 3.340515f **FLOATING
C566 mid_6to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# VSUBS 3.34045f **FLOATING
C567 mid_6to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# VSUBS 3.34045f **FLOATING
C568 mid_6to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# VSUBS 3.34045f **FLOATING
C569 mid_6to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# VSUBS 3.337859f **FLOATING
C570 mid_6to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# VSUBS 3.34045f **FLOATING
C571 mid_6to8_3/8_cap_array_final_1/m1_n130_1630# VSUBS 6.903774f
C572 mid_6to8_3/8_cap_array_final_1/m1_n130_1750# VSUBS 2.161829f
C573 mid_6to8_3/8_cap_array_final_1/m1_n130_1870# VSUBS 2.166234f
C574 mid_6to8_3/8_cap_array_final_1/m1_n130_1990# VSUBS 2.174879f
C575 mid_6to8_3/8_cap_array_final_1/m1_n130_2110# VSUBS 2.193039f
C576 mid_6to8_3/8_cap_array_final_1/m1_n130_3980# VSUBS 2.15064f
C577 mid_6to8_3/8_cap_array_final_1/m1_n130_4100# VSUBS 2.15295f
C578 mid_6to8_3/8_cap_array_final_1/m1_n130_4220# VSUBS 2.15295f
C579 mid_6to8_3/8_cap_array_final_1/m1_n130_4340# VSUBS 2.15295f
C580 mid_6to8_3/8_cap_array_final_1/m1_n130_4460# VSUBS 6.89743f
C581 mid_6to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# VSUBS 3.34045f **FLOATING
C582 mid_6to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# VSUBS 3.34045f **FLOATING
C583 mid_6to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# VSUBS 3.34045f **FLOATING
C584 mid_6to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# VSUBS 3.340515f **FLOATING
C585 mid_6to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# VSUBS 3.340515f **FLOATING
C586 mid_6to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C587 mid_6to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# VSUBS 3.34045f **FLOATING
C588 mid_6to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# VSUBS 3.47539f **FLOATING
C589 end_3/8_cap_array_final_1/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C590 end_3/8_cap_array_final_1/cap_final_6/m1_990_n540# VSUBS 3.340515f **FLOATING
C591 end_3/8_cap_array_final_1/cap_final_5/m1_990_n540# VSUBS 3.340515f **FLOATING
C592 end_3/8_cap_array_final_1/cap_final_4/m1_990_n540# VSUBS 3.340515f **FLOATING
C593 end_3/8_cap_array_final_1/cap_final_3/m1_990_n540# VSUBS 3.340515f **FLOATING
C594 end_3/8_cap_array_final_1/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C595 end_3/8_cap_array_final_1/cap_final_1/m1_990_n540# VSUBS 3.337859f **FLOATING
C596 end_3/8_cap_array_final_1/cap_final_0/m1_990_n540# VSUBS 3.340514f **FLOATING
C597 end_3/8_cap_array_final_1/m1_n130_1630# VSUBS 6.903774f
C598 end_3/8_cap_array_final_1/m1_n130_1750# VSUBS 2.161829f
C599 end_3/8_cap_array_final_1/m1_n130_1870# VSUBS 2.166234f
C600 end_3/8_cap_array_final_1/m1_n130_1990# VSUBS 2.174879f
C601 end_3/8_cap_array_final_1/m1_n130_2110# VSUBS 2.195349f
C602 end_3/8_cap_array_final_1/m1_n130_2230# VSUBS 3.840402f
C603 end_3/8_cap_array_final_1/m1_n130_3860# VSUBS 3.732141f
C604 end_3/8_cap_array_final_1/m1_n130_3980# VSUBS 2.15295f
C605 end_3/8_cap_array_final_1/m1_n130_4100# VSUBS 2.15295f
C606 end_3/8_cap_array_final_1/m1_n130_4220# VSUBS 2.15295f
C607 end_3/8_cap_array_final_1/m1_n130_4340# VSUBS 2.15295f
C608 end_3/8_cap_array_final_1/m1_n130_4460# VSUBS 6.89743f
C609 end_3/8_cap_array_final_0/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C610 end_3/8_cap_array_final_0/cap_final_6/m1_990_n540# VSUBS 3.340515f **FLOATING
C611 end_3/8_cap_array_final_0/cap_final_5/m1_990_n540# VSUBS 3.340515f **FLOATING
C612 end_3/8_cap_array_final_0/cap_final_4/m1_990_n540# VSUBS 3.340515f **FLOATING
C613 end_3/8_cap_array_final_0/cap_final_3/m1_990_n540# VSUBS 3.340515f **FLOATING
C614 end_3/8_cap_array_final_0/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C615 end_3/8_cap_array_final_0/cap_final_1/m1_990_n540# VSUBS 3.340514f **FLOATING
C616 end_3/8_cap_array_final_0/cap_final_0/m1_990_n540# VSUBS 3.47539f **FLOATING
C617 end_2/8_cap_array_final_1/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C618 end_2/8_cap_array_final_1/cap_final_6/m1_990_n540# VSUBS 3.340515f **FLOATING
C619 end_2/8_cap_array_final_1/cap_final_5/m1_990_n540# VSUBS 3.340515f **FLOATING
C620 end_2/8_cap_array_final_1/cap_final_4/m1_990_n540# VSUBS 3.340515f **FLOATING
C621 end_2/8_cap_array_final_1/cap_final_3/m1_990_n540# VSUBS 3.340515f **FLOATING
C622 end_2/8_cap_array_final_1/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C623 end_2/8_cap_array_final_1/cap_final_1/m1_990_n540# VSUBS 3.337859f **FLOATING
C624 end_2/8_cap_array_final_1/cap_final_0/m1_990_n540# VSUBS 3.340514f **FLOATING
C625 end_2/8_cap_array_final_1/m1_n130_1630# VSUBS 6.903774f
C626 end_2/8_cap_array_final_1/m1_n130_1750# VSUBS 2.161829f
C627 end_2/8_cap_array_final_1/m1_n130_1870# VSUBS 2.166234f
C628 end_2/8_cap_array_final_1/m1_n130_1990# VSUBS 2.174879f
C629 end_2/8_cap_array_final_1/m1_n130_2110# VSUBS 2.195349f
C630 end_2/8_cap_array_final_1/m1_n130_2230# VSUBS 3.840402f
C631 end_2/8_cap_array_final_1/m1_n130_3860# VSUBS 3.732141f
C632 end_2/8_cap_array_final_1/m1_n130_3980# VSUBS 2.15295f
C633 end_2/8_cap_array_final_1/m1_n130_4100# VSUBS 2.15295f
C634 end_2/8_cap_array_final_1/m1_n130_4220# VSUBS 2.15295f
C635 end_2/8_cap_array_final_1/m1_n130_4340# VSUBS 2.15295f
C636 end_2/8_cap_array_final_1/m1_n130_4460# VSUBS 6.89743f
C637 end_2/8_cap_array_final_0/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C638 end_2/8_cap_array_final_0/cap_final_6/m1_990_n540# VSUBS 3.340515f **FLOATING
C639 end_2/8_cap_array_final_0/cap_final_5/m1_990_n540# VSUBS 3.340515f **FLOATING
C640 end_2/8_cap_array_final_0/cap_final_4/m1_990_n540# VSUBS 3.340515f **FLOATING
C641 end_2/8_cap_array_final_0/cap_final_3/m1_990_n540# VSUBS 3.340515f **FLOATING
C642 end_2/8_cap_array_final_0/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C643 end_2/8_cap_array_final_0/cap_final_1/m1_990_n540# VSUBS 3.340514f **FLOATING
C644 end_2/8_cap_array_final_0/cap_final_0/m1_990_n540# VSUBS 3.47539f **FLOATING
C645 mid_6to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C646 mid_6to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# VSUBS 3.340515f **FLOATING
C647 mid_6to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# VSUBS 3.340515f **FLOATING
C648 mid_6to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# VSUBS 3.34045f **FLOATING
C649 mid_6to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# VSUBS 3.34045f **FLOATING
C650 mid_6to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# VSUBS 3.34045f **FLOATING
C651 mid_6to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# VSUBS 3.337859f **FLOATING
C652 mid_6to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# VSUBS 3.34045f **FLOATING
C653 mid_6to8_2/8_cap_array_final_1/m1_n130_1630# VSUBS 6.903774f
C654 mid_6to8_2/8_cap_array_final_1/m1_n130_1750# VSUBS 2.161829f
C655 mid_6to8_2/8_cap_array_final_1/m1_n130_1870# VSUBS 2.166234f
C656 mid_6to8_2/8_cap_array_final_1/m1_n130_1990# VSUBS 2.174879f
C657 mid_6to8_2/8_cap_array_final_1/m1_n130_2110# VSUBS 2.193039f
C658 mid_6to8_2/8_cap_array_final_1/m1_n130_3980# VSUBS 2.15064f
C659 mid_6to8_2/8_cap_array_final_1/m1_n130_4100# VSUBS 2.15295f
C660 mid_6to8_2/8_cap_array_final_1/m1_n130_4220# VSUBS 2.15295f
C661 mid_6to8_2/8_cap_array_final_1/m1_n130_4340# VSUBS 2.15295f
C662 mid_6to8_2/8_cap_array_final_1/m1_n130_4460# VSUBS 6.89743f
C663 mid_6to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# VSUBS 3.34045f **FLOATING
C664 mid_6to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# VSUBS 3.34045f **FLOATING
C665 mid_6to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# VSUBS 3.34045f **FLOATING
C666 mid_6to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# VSUBS 3.340515f **FLOATING
C667 mid_6to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# VSUBS 3.340515f **FLOATING
C668 mid_6to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C669 mid_6to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# VSUBS 3.34045f **FLOATING
C670 mid_6to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# VSUBS 3.47539f **FLOATING
C671 end_1/8_cap_array_final_1/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C672 end_1/8_cap_array_final_1/cap_final_6/m1_990_n540# VSUBS 3.340515f **FLOATING
C673 end_1/8_cap_array_final_1/cap_final_5/m1_990_n540# VSUBS 3.340515f **FLOATING
C674 end_1/8_cap_array_final_1/cap_final_4/m1_990_n540# VSUBS 3.340515f **FLOATING
C675 end_1/8_cap_array_final_1/cap_final_3/m1_990_n540# VSUBS 3.340515f **FLOATING
C676 end_1/8_cap_array_final_1/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C677 end_1/8_cap_array_final_1/cap_final_1/m1_990_n540# VSUBS 3.337859f **FLOATING
C678 end_1/8_cap_array_final_1/cap_final_0/m1_990_n540# VSUBS 3.340514f **FLOATING
C679 end_1/8_cap_array_final_1/m1_n130_1630# VSUBS 6.903774f
C680 end_1/8_cap_array_final_1/m1_n130_1750# VSUBS 2.161829f
C681 end_1/8_cap_array_final_1/m1_n130_1870# VSUBS 2.166234f
C682 end_1/8_cap_array_final_1/m1_n130_1990# VSUBS 2.174879f
C683 end_1/8_cap_array_final_1/m1_n130_2110# VSUBS 2.195349f
C684 end_1/8_cap_array_final_1/m1_n130_2230# VSUBS 3.840402f
C685 end_1/8_cap_array_final_1/m1_n130_3860# VSUBS 3.732141f
C686 end_1/8_cap_array_final_1/m1_n130_3980# VSUBS 2.15295f
C687 end_1/8_cap_array_final_1/m1_n130_4100# VSUBS 2.15295f
C688 end_1/8_cap_array_final_1/m1_n130_4220# VSUBS 2.15295f
C689 end_1/8_cap_array_final_1/m1_n130_4340# VSUBS 2.15295f
C690 end_1/8_cap_array_final_1/m1_n130_4460# VSUBS 6.89743f
C691 end_1/8_cap_array_final_0/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C692 end_1/8_cap_array_final_0/cap_final_6/m1_990_n540# VSUBS 3.340515f **FLOATING
C693 end_1/8_cap_array_final_0/cap_final_5/m1_990_n540# VSUBS 3.340515f **FLOATING
C694 end_1/8_cap_array_final_0/cap_final_4/m1_990_n540# VSUBS 3.340515f **FLOATING
C695 end_1/8_cap_array_final_0/cap_final_3/m1_990_n540# VSUBS 3.340515f **FLOATING
C696 end_1/8_cap_array_final_0/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C697 end_1/8_cap_array_final_0/cap_final_1/m1_990_n540# VSUBS 3.340514f **FLOATING
C698 end_1/8_cap_array_final_0/cap_final_0/m1_990_n540# VSUBS 3.47539f **FLOATING
C699 mid_6to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C700 mid_6to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# VSUBS 3.340515f **FLOATING
C701 mid_6to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# VSUBS 3.340515f **FLOATING
C702 mid_6to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# VSUBS 3.34045f **FLOATING
C703 mid_6to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# VSUBS 3.34045f **FLOATING
C704 mid_6to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# VSUBS 3.34045f **FLOATING
C705 mid_6to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# VSUBS 3.337859f **FLOATING
C706 mid_6to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# VSUBS 3.34045f **FLOATING
C707 mid_6to8_1/8_cap_array_final_1/m1_n130_1630# VSUBS 6.903774f
C708 mid_6to8_1/8_cap_array_final_1/m1_n130_1750# VSUBS 2.161829f
C709 mid_6to8_1/8_cap_array_final_1/m1_n130_1870# VSUBS 2.166234f
C710 mid_6to8_1/8_cap_array_final_1/m1_n130_1990# VSUBS 2.174879f
C711 mid_6to8_1/8_cap_array_final_1/m1_n130_2110# VSUBS 2.193039f
C712 mid_6to8_1/8_cap_array_final_1/m1_n130_3980# VSUBS 2.15064f
C713 mid_6to8_1/8_cap_array_final_1/m1_n130_4100# VSUBS 2.15295f
C714 mid_6to8_1/8_cap_array_final_1/m1_n130_4220# VSUBS 2.15295f
C715 mid_6to8_1/8_cap_array_final_1/m1_n130_4340# VSUBS 2.15295f
C716 mid_6to8_1/8_cap_array_final_1/m1_n130_4460# VSUBS 6.89743f
C717 mid_6to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# VSUBS 3.34045f **FLOATING
C718 mid_6to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# VSUBS 3.34045f **FLOATING
C719 mid_6to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# VSUBS 3.34045f **FLOATING
C720 mid_6to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# VSUBS 3.340515f **FLOATING
C721 mid_6to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# VSUBS 3.340515f **FLOATING
C722 mid_6to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C723 mid_6to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# VSUBS 3.34045f **FLOATING
C724 mid_6to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# VSUBS 3.47539f **FLOATING
C725 end_0/8_cap_array_final_1/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C726 end_0/8_cap_array_final_1/cap_final_6/m1_990_n540# VSUBS 3.340515f **FLOATING
C727 end_0/8_cap_array_final_1/cap_final_5/m1_990_n540# VSUBS 3.340515f **FLOATING
C728 end_0/8_cap_array_final_1/cap_final_4/m1_990_n540# VSUBS 3.340515f **FLOATING
C729 end_0/8_cap_array_final_1/cap_final_3/m1_990_n540# VSUBS 3.340515f **FLOATING
C730 end_0/8_cap_array_final_1/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C731 end_0/8_cap_array_final_1/cap_final_1/m1_990_n540# VSUBS 3.337859f **FLOATING
C732 end_0/8_cap_array_final_1/cap_final_0/m1_990_n540# VSUBS 3.340514f **FLOATING
C733 end_0/8_cap_array_final_1/m1_n130_1630# VSUBS 6.903774f
C734 end_0/8_cap_array_final_1/m1_n130_1750# VSUBS 2.161829f
C735 end_0/8_cap_array_final_1/m1_n130_1870# VSUBS 2.166234f
C736 end_0/8_cap_array_final_1/m1_n130_1990# VSUBS 2.174879f
C737 end_0/8_cap_array_final_1/m1_n130_2110# VSUBS 2.195349f
C738 end_0/8_cap_array_final_1/m1_n130_2230# VSUBS 3.840402f
C739 end_0/8_cap_array_final_1/m1_n130_3860# VSUBS 3.732141f
C740 end_0/8_cap_array_final_1/m1_n130_3980# VSUBS 2.15295f
C741 end_0/8_cap_array_final_1/m1_n130_4100# VSUBS 2.15295f
C742 end_0/8_cap_array_final_1/m1_n130_4220# VSUBS 2.15295f
C743 end_0/8_cap_array_final_1/m1_n130_4340# VSUBS 2.15295f
C744 end_0/8_cap_array_final_1/m1_n130_4460# VSUBS 6.89743f
C745 end_0/8_cap_array_final_0/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C746 end_0/8_cap_array_final_0/cap_final_6/m1_990_n540# VSUBS 3.340515f **FLOATING
C747 end_0/8_cap_array_final_0/cap_final_5/m1_990_n540# VSUBS 3.340515f **FLOATING
C748 end_0/8_cap_array_final_0/cap_final_4/m1_990_n540# VSUBS 3.340515f **FLOATING
C749 end_0/8_cap_array_final_0/cap_final_3/m1_990_n540# VSUBS 3.340515f **FLOATING
C750 end_3/8_cap_array_final_1/cap_final_7/phi2 VSUBS 0.349631p
C751 end_3/8_cap_array_final_1/cap_final_7/phi2_n VSUBS 68.62323f
C752 end_3/8_cap_array_final_1/cap_final_7/com_x VSUBS 0.124438p
C753 end_0/8_cap_array_final_0/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C754 end_3/8_cap_array_final_1/cap_final_7/Vin VSUBS 0.115036p
C755 end_3/8_cap_array_final_1/cap_final_7/Vdd VSUBS 0.491736p
C756 end_3/8_cap_array_final_1/cap_final_7/GND VSUBS 0.126217p
C757 end_0/8_cap_array_final_0/cap_final_1/m1_990_n540# VSUBS 3.340514f **FLOATING
C758 end_0/8_cap_array_final_0/cap_final_0/m1_990_n540# VSUBS 3.47539f **FLOATING
C759 end_3/8_cap_array_final_1/cap_final_7/phi1 VSUBS 0.137739p
C760 end_3/8_cap_array_final_1/cap_final_7/phi1_n VSUBS 95.42289f
C761 mid_6to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C762 mid_6to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# VSUBS 3.340515f **FLOATING
C763 mid_6to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# VSUBS 3.340515f **FLOATING
C764 mid_6to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# VSUBS 3.34045f **FLOATING
C765 mid_6to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# VSUBS 3.34045f **FLOATING
C766 mid_6to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# VSUBS 3.34045f **FLOATING
C767 mid_6to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# VSUBS 3.337859f **FLOATING
C768 mid_6to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# VSUBS 3.34045f **FLOATING
C769 mid_6to8_0/8_cap_array_final_1/m1_n130_1630# VSUBS 6.903774f
C770 mid_6to8_0/8_cap_array_final_1/m1_n130_1750# VSUBS 2.161829f
C771 mid_6to8_0/8_cap_array_final_1/m1_n130_1870# VSUBS 2.166234f
C772 mid_6to8_0/8_cap_array_final_1/m1_n130_1990# VSUBS 2.174879f
C773 mid_6to8_0/8_cap_array_final_1/m1_n130_2110# VSUBS 2.193039f
C774 mid_2_0/8_cap_array_final_0/cap_final_6/phi2_n VSUBS 60.79054f
C775 mid_6to8_0/8_cap_array_final_1/m1_n130_3980# VSUBS 2.15064f
C776 mid_6to8_0/8_cap_array_final_1/m1_n130_4100# VSUBS 2.15295f
C777 mid_6to8_0/8_cap_array_final_1/m1_n130_4220# VSUBS 2.15295f
C778 mid_6to8_0/8_cap_array_final_1/m1_n130_4340# VSUBS 2.15295f
C779 mid_6to8_0/8_cap_array_final_1/m1_n130_4460# VSUBS 6.89743f
C780 mid_6to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# VSUBS 3.34045f **FLOATING
C781 mid_6to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# VSUBS 3.34045f **FLOATING
C782 mid_6to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# VSUBS 3.34045f **FLOATING
C783 mid_2_0/8_cap_array_final_0/cap_final_6/phi1 VSUBS 60.502262f
C784 mid_2_0/8_cap_array_final_0/cap_final_6/phi1_n VSUBS 53.56026f
C785 mid_2_0/8_cap_array_final_0/cap_final_6/phi2 VSUBS 75.70891f
C786 mid_6to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# VSUBS 3.340515f **FLOATING
C787 mid_6to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# VSUBS 3.340515f **FLOATING
C788 mid_6to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C789 mid_6to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# VSUBS 3.34045f **FLOATING
C790 mid_6to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# VSUBS 3.47539f **FLOATING
C791 mid_2to4__1/8_cap_array_final_1/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C792 mid_2to4__1/8_cap_array_final_1/cap_final_6/m1_990_n540# VSUBS 3.34045f **FLOATING
C793 mid_2to4__1/8_cap_array_final_1/cap_final_5/m1_990_n540# VSUBS 3.34045f **FLOATING
C794 mid_2to4__1/8_cap_array_final_1/cap_final_4/m1_990_n540# VSUBS 3.34039f **FLOATING
C795 mid_2to4__1/8_cap_array_final_1/cap_final_3/m1_990_n540# VSUBS 3.340337f **FLOATING
C796 mid_2to4__1/8_cap_array_final_1/cap_final_2/m1_990_n540# VSUBS 3.340289f **FLOATING
C797 mid_2to4__1/8_cap_array_final_1/cap_final_1/m1_990_n540# VSUBS 3.337859f **FLOATING
C798 mid_2to4__1/8_cap_array_final_1/cap_final_0/m1_990_n540# VSUBS 3.340247f **FLOATING
C799 mid_2to4__1/8_cap_array_final_1/m1_n130_1630# VSUBS 6.902235f
C800 mid_2to4__1/8_cap_array_final_1/m1_n130_4460# VSUBS 6.89589f
C801 mid_2to4__1/8_cap_array_final_0/cap_final_7/m1_990_n540# VSUBS 3.340289f **FLOATING
C802 mid_2to4__1/8_cap_array_final_0/cap_final_6/m1_990_n540# VSUBS 3.340337f **FLOATING
C803 mid_2to4__1/8_cap_array_final_0/cap_final_5/m1_990_n540# VSUBS 3.34039f **FLOATING
C804 mid_2to4__1/8_cap_array_final_0/cap_final_4/m1_990_n540# VSUBS 3.34045f **FLOATING
C805 mid_2to4__1/8_cap_array_final_0/cap_final_3/m1_990_n540# VSUBS 3.34045f **FLOATING
C806 mid_2to4__1/8_cap_array_final_0/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C807 mid_2to4__1/8_cap_array_final_0/cap_final_1/m1_990_n540# VSUBS 3.340247f **FLOATING
C808 mid_2to4__1/8_cap_array_final_0/cap_final_0/m1_990_n540# VSUBS 3.47539f **FLOATING
C809 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2 VSUBS 6.866877f
C810 mid_2to4__0/8_cap_array_final_1/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C811 mid_2to4__0/8_cap_array_final_1/cap_final_6/m1_990_n540# VSUBS 3.34045f **FLOATING
C812 mid_2to4__0/8_cap_array_final_1/cap_final_5/m1_990_n540# VSUBS 3.34045f **FLOATING
C813 mid_2to4__0/8_cap_array_final_1/cap_final_4/m1_990_n540# VSUBS 3.34039f **FLOATING
C814 mid_2to4__0/8_cap_array_final_1/cap_final_3/m1_990_n540# VSUBS 3.340337f **FLOATING
C815 mid_2to4__0/8_cap_array_final_1/cap_final_2/m1_990_n540# VSUBS 3.340289f **FLOATING
C816 mid_2to4__0/8_cap_array_final_1/cap_final_1/m1_990_n540# VSUBS 3.337859f **FLOATING
C817 mid_2to4__0/8_cap_array_final_1/cap_final_0/m1_990_n540# VSUBS 3.340247f **FLOATING
C818 mid_2to4__0/8_cap_array_final_1/m1_n130_1630# VSUBS 6.902235f
C819 mid_2to4__0/8_cap_array_final_1/m1_n130_4460# VSUBS 6.89589f
C820 mid_2to4__0/8_cap_array_final_0/cap_final_7/m1_990_n540# VSUBS 3.340289f **FLOATING
C821 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1 VSUBS 6.695977f
C822 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi1_n VSUBS 11.111129f
C823 mid_2to4__1/8_cap_array_final_1/cap_final_2/phi2_n VSUBS 10.412113f
C824 mid_2to4__0/8_cap_array_final_0/cap_final_6/m1_990_n540# VSUBS 3.340337f **FLOATING
C825 mid_2to4__0/8_cap_array_final_0/cap_final_5/m1_990_n540# VSUBS 3.34039f **FLOATING
C826 mid_2to4__0/8_cap_array_final_0/cap_final_4/m1_990_n540# VSUBS 3.34045f **FLOATING
C827 mid_2to4__0/8_cap_array_final_0/cap_final_3/m1_990_n540# VSUBS 3.34045f **FLOATING
C828 mid_2to4__0/8_cap_array_final_0/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C829 mid_2to4__0/8_cap_array_final_0/cap_final_1/m1_990_n540# VSUBS 3.340247f **FLOATING
C830 mid_2to4__0/8_cap_array_final_0/cap_final_0/m1_990_n540# VSUBS 3.47539f **FLOATING
C831 mid_4to8_2/8_cap_array_final_1/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C832 mid_4to8_2/8_cap_array_final_1/cap_final_6/m1_990_n540# VSUBS 3.34045f **FLOATING
C833 mid_4to8_2/8_cap_array_final_1/cap_final_5/m1_990_n540# VSUBS 3.34045f **FLOATING
C834 mid_4to8_2/8_cap_array_final_1/cap_final_4/m1_990_n540# VSUBS 3.34039f **FLOATING
C835 mid_4to8_2/8_cap_array_final_1/cap_final_3/m1_990_n540# VSUBS 3.340337f **FLOATING
C836 mid_4to8_2/8_cap_array_final_1/cap_final_2/m1_990_n540# VSUBS 3.340337f **FLOATING
C837 mid_4to8_2/8_cap_array_final_1/cap_final_1/m1_990_n540# VSUBS 3.337859f **FLOATING
C838 mid_4to8_2/8_cap_array_final_1/cap_final_0/m1_990_n540# VSUBS 3.340337f **FLOATING
C839 mid_4to8_2/8_cap_array_final_1/m1_n130_1630# VSUBS 6.903774f
C840 mid_4to8_2/8_cap_array_final_1/m1_n130_1750# VSUBS 2.161829f
C841 mid_4to8_2/8_cap_array_final_1/m1_n130_1870# VSUBS 2.163925f
C842 mid_4to8_2/8_cap_array_final_1/m1_n130_4220# VSUBS 2.15064f
C843 mid_4to8_2/8_cap_array_final_1/m1_n130_4340# VSUBS 2.15295f
C844 mid_4to8_2/8_cap_array_final_1/m1_n130_4460# VSUBS 6.89743f
C845 mid_4to8_2/8_cap_array_final_0/cap_final_7/m1_990_n540# VSUBS 3.340337f **FLOATING
C846 mid_4to8_2/8_cap_array_final_0/cap_final_6/m1_990_n540# VSUBS 3.340337f **FLOATING
C847 mid_4to8_2/8_cap_array_final_0/cap_final_5/m1_990_n540# VSUBS 3.34039f **FLOATING
C848 mid_4to8_2/8_cap_array_final_0/cap_final_4/m1_990_n540# VSUBS 3.34045f **FLOATING
C849 mid_4to8_2/8_cap_array_final_0/cap_final_3/m1_990_n540# VSUBS 3.34045f **FLOATING
C850 mid_4to8_2/8_cap_array_final_0/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C851 mid_4to8_2/8_cap_array_final_0/cap_final_1/m1_990_n540# VSUBS 3.340337f **FLOATING
C852 mid_4to8_2/8_cap_array_final_0/cap_final_0/m1_990_n540# VSUBS 3.47539f **FLOATING
C853 mid_4to8_3/8_cap_array_final_1/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C854 mid_4to8_3/8_cap_array_final_1/cap_final_6/m1_990_n540# VSUBS 3.34045f **FLOATING
C855 mid_4to8_3/8_cap_array_final_1/cap_final_5/m1_990_n540# VSUBS 3.34045f **FLOATING
C856 mid_4to8_3/8_cap_array_final_1/cap_final_4/m1_990_n540# VSUBS 3.34039f **FLOATING
C857 mid_4to8_3/8_cap_array_final_1/cap_final_3/m1_990_n540# VSUBS 3.340337f **FLOATING
C858 mid_4to8_3/8_cap_array_final_1/cap_final_2/m1_990_n540# VSUBS 3.340337f **FLOATING
C859 mid_4to8_3/8_cap_array_final_1/cap_final_1/m1_990_n540# VSUBS 3.337859f **FLOATING
C860 mid_4to8_3/8_cap_array_final_1/cap_final_0/m1_990_n540# VSUBS 3.340337f **FLOATING
C861 mid_4to8_3/8_cap_array_final_1/m1_n130_1630# VSUBS 6.903774f
C862 mid_4to8_3/8_cap_array_final_1/m1_n130_1750# VSUBS 2.161829f
C863 mid_4to8_3/8_cap_array_final_1/m1_n130_1870# VSUBS 2.163925f
C864 mid_4to8_3/8_cap_array_final_1/m1_n130_4220# VSUBS 2.15064f
C865 mid_4to8_3/8_cap_array_final_1/m1_n130_4340# VSUBS 2.15295f
C866 mid_4to8_3/8_cap_array_final_1/m1_n130_4460# VSUBS 6.89743f
C867 mid_4to8_3/8_cap_array_final_0/cap_final_7/m1_990_n540# VSUBS 3.340337f **FLOATING
C868 mid_4to8_3/8_cap_array_final_0/cap_final_6/m1_990_n540# VSUBS 3.340337f **FLOATING
C869 mid_4to8_3/8_cap_array_final_0/cap_final_5/m1_990_n540# VSUBS 3.34039f **FLOATING
C870 mid_4to8_3/8_cap_array_final_0/cap_final_4/m1_990_n540# VSUBS 3.34045f **FLOATING
C871 mid_4to8_3/8_cap_array_final_0/cap_final_3/m1_990_n540# VSUBS 3.34045f **FLOATING
C872 mid_4to8_3/8_cap_array_final_0/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C873 mid_4to8_3/8_cap_array_final_0/cap_final_1/m1_990_n540# VSUBS 3.340337f **FLOATING
C874 mid_4to8_3/8_cap_array_final_0/cap_final_0/m1_990_n540# VSUBS 3.47539f **FLOATING
C875 mid_4to8_1/8_cap_array_final_1/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C876 mid_4to8_1/8_cap_array_final_1/cap_final_6/m1_990_n540# VSUBS 3.34045f **FLOATING
C877 mid_4to8_1/8_cap_array_final_1/cap_final_5/m1_990_n540# VSUBS 3.34045f **FLOATING
C878 mid_4to8_1/8_cap_array_final_1/cap_final_4/m1_990_n540# VSUBS 3.34039f **FLOATING
C879 mid_4to8_1/8_cap_array_final_1/cap_final_3/m1_990_n540# VSUBS 3.340337f **FLOATING
C880 mid_4to8_1/8_cap_array_final_1/cap_final_2/m1_990_n540# VSUBS 3.340337f **FLOATING
C881 mid_4to8_1/8_cap_array_final_1/cap_final_1/m1_990_n540# VSUBS 3.337859f **FLOATING
C882 mid_4to8_1/8_cap_array_final_1/cap_final_0/m1_990_n540# VSUBS 3.340337f **FLOATING
C883 mid_4to8_1/8_cap_array_final_1/m1_n130_1630# VSUBS 6.903774f
C884 mid_4to8_1/8_cap_array_final_1/m1_n130_1750# VSUBS 2.161829f
C885 mid_4to8_1/8_cap_array_final_1/m1_n130_1870# VSUBS 2.163925f
C886 mid_4to8_1/8_cap_array_final_1/m1_n130_4220# VSUBS 2.15064f
C887 mid_4to8_1/8_cap_array_final_1/m1_n130_4340# VSUBS 2.15295f
C888 mid_4to8_1/8_cap_array_final_1/m1_n130_4460# VSUBS 6.89743f
C889 mid_4to8_1/8_cap_array_final_0/cap_final_7/m1_990_n540# VSUBS 3.340337f **FLOATING
C890 mid_4to8_1/8_cap_array_final_0/cap_final_6/m1_990_n540# VSUBS 3.340337f **FLOATING
C891 mid_4to8_1/8_cap_array_final_0/cap_final_5/m1_990_n540# VSUBS 3.34039f **FLOATING
C892 mid_4to8_1/8_cap_array_final_0/cap_final_4/m1_990_n540# VSUBS 3.34045f **FLOATING
C893 mid_4to8_1/8_cap_array_final_0/cap_final_3/m1_990_n540# VSUBS 3.34045f **FLOATING
C894 mid_4to8_1/8_cap_array_final_0/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C895 mid_4to8_1/8_cap_array_final_0/cap_final_1/m1_990_n540# VSUBS 3.340337f **FLOATING
C896 mid_4to8_1/8_cap_array_final_0/cap_final_0/m1_990_n540# VSUBS 3.47539f **FLOATING
C897 mid_2_0/8_cap_array_final_0/cap_final_4/phi2 VSUBS 34.161232f
C898 mid_2_0/8_cap_array_final_0/cap_final_3/phi2_n VSUBS 23.373602f
C899 mid_2_0/8_cap_array_final_0/cap_final_4/phi2_n VSUBS 28.795658f
C900 mid_4to8_0/8_cap_array_final_1/cap_final_7/m1_990_n540# VSUBS 3.340515f **FLOATING
C901 mid_4to8_0/8_cap_array_final_1/cap_final_6/m1_990_n540# VSUBS 3.34045f **FLOATING
C902 mid_4to8_0/8_cap_array_final_1/cap_final_5/m1_990_n540# VSUBS 3.34045f **FLOATING
C903 mid_4to8_0/8_cap_array_final_1/cap_final_4/m1_990_n540# VSUBS 3.34039f **FLOATING
C904 mid_4to8_0/8_cap_array_final_1/cap_final_3/m1_990_n540# VSUBS 3.340337f **FLOATING
C905 mid_4to8_0/8_cap_array_final_1/cap_final_2/m1_990_n540# VSUBS 3.340337f **FLOATING
C906 mid_4to8_0/8_cap_array_final_1/cap_final_1/m1_990_n540# VSUBS 3.337859f **FLOATING
C907 mid_4to8_0/8_cap_array_final_1/cap_final_0/m1_990_n540# VSUBS 3.340337f **FLOATING
C908 mid_4to8_0/8_cap_array_final_1/m1_n130_1630# VSUBS 6.903774f
C909 mid_4to8_0/8_cap_array_final_1/m1_n130_1750# VSUBS 2.161829f
C910 mid_4to8_0/8_cap_array_final_1/m1_n130_1870# VSUBS 2.163925f
C911 mid_2_0/8_cap_array_final_0/cap_final_3/phi2 VSUBS 22.839111f
C912 mid_4to8_0/8_cap_array_final_1/m1_n130_4220# VSUBS 2.15064f
C913 mid_4to8_0/8_cap_array_final_1/m1_n130_4340# VSUBS 2.15295f
C914 mid_4to8_0/8_cap_array_final_1/m1_n130_4460# VSUBS 6.89743f
C915 mid_4to8_0/8_cap_array_final_0/cap_final_7/m1_990_n540# VSUBS 3.340337f **FLOATING
C916 mid_4to8_0/8_cap_array_final_0/cap_final_6/m1_990_n540# VSUBS 3.340337f **FLOATING
C917 mid_2_0/8_cap_array_final_0/cap_final_4/phi1 VSUBS 33.817f
C918 mid_2_0/8_cap_array_final_0/cap_final_4/phi1_n VSUBS 34.07063f
C919 mid_4to8_0/8_cap_array_final_0/cap_final_5/m1_990_n540# VSUBS 3.34039f **FLOATING
C920 mid_2_0/8_cap_array_final_0/cap_final_3/phi1 VSUBS 20.157578f
C921 mid_2_0/8_cap_array_final_0/cap_final_3/phi1_n VSUBS 22.736082f
C922 mid_4to8_0/8_cap_array_final_0/cap_final_4/m1_990_n540# VSUBS 3.34045f **FLOATING
C923 mid_4to8_0/8_cap_array_final_0/cap_final_3/m1_990_n540# VSUBS 3.34045f **FLOATING
C924 mid_4to8_0/8_cap_array_final_0/cap_final_2/m1_990_n540# VSUBS 3.340515f **FLOATING
C925 mid_4to8_0/8_cap_array_final_0/cap_final_1/m1_990_n540# VSUBS 3.340337f **FLOATING
C926 mid_4to8_0/8_cap_array_final_0/cap_final_0/m1_990_n540# VSUBS 3.47539f **FLOATING
