magic
tech sky130A
timestamp 1730665161
<< metal1 >>
rect 4760 2180 4765 2195
rect 0 2165 4685 2180
rect 4715 2165 4765 2180
rect 4795 2180 4800 2195
rect 5615 2180 5620 2195
rect 4795 2165 5540 2180
rect 5570 2165 5620 2180
rect 5650 2180 5655 2195
rect 6470 2180 6475 2195
rect 5650 2165 6395 2180
rect 6425 2165 6475 2180
rect 6505 2180 6510 2195
rect 7325 2180 7330 2195
rect 6505 2165 7250 2180
rect 7280 2165 7330 2180
rect 7360 2180 7365 2195
rect 8180 2180 8185 2195
rect 7360 2165 8105 2180
rect 8135 2165 8185 2180
rect 8215 2180 8220 2195
rect 9035 2180 9040 2195
rect 8215 2165 8960 2180
rect 8990 2165 9040 2180
rect 9070 2180 9075 2195
rect 9070 2165 13680 2180
rect 3905 2120 3910 2135
rect 0 2105 3830 2120
rect 3860 2105 3910 2120
rect 3940 2120 3945 2135
rect 9890 2120 9895 2135
rect 3940 2105 4685 2120
rect 4715 2105 5540 2120
rect 5570 2105 6395 2120
rect 6425 2105 7250 2120
rect 7280 2105 8105 2120
rect 8135 2105 8960 2120
rect 8990 2105 9815 2120
rect 9845 2105 9895 2120
rect 9925 2120 9930 2135
rect 9925 2105 13680 2120
rect 2195 2060 2200 2075
rect 0 2045 2200 2060
rect 2230 2060 2235 2075
rect 3050 2060 3055 2075
rect 2230 2045 3055 2060
rect 3085 2060 3090 2075
rect 10740 2060 10745 2075
rect 3085 2045 3830 2060
rect 3860 2045 4685 2060
rect 4715 2045 5540 2060
rect 5570 2045 6395 2060
rect 6425 2045 7250 2060
rect 7280 2045 8105 2060
rect 8135 2045 8960 2060
rect 8990 2045 9815 2060
rect 9845 2045 10670 2060
rect 10700 2045 10745 2060
rect 10775 2060 10780 2075
rect 11600 2060 11605 2075
rect 10775 2045 11525 2060
rect 11555 2045 11605 2060
rect 11635 2060 11640 2075
rect 11635 2045 13680 2060
rect 485 2000 490 2015
rect 0 1985 490 2000
rect 520 2000 525 2015
rect 1340 2000 1345 2015
rect 520 1985 1345 2000
rect 1375 2000 1380 2015
rect 12455 2000 12460 2015
rect 1375 1985 4685 2000
rect 4715 1985 5540 2000
rect 5570 1985 6395 2000
rect 6425 1985 7250 2000
rect 7280 1985 8105 2000
rect 8135 1985 8960 2000
rect 8990 1985 9815 2000
rect 9845 1985 10670 2000
rect 10700 1985 11525 2000
rect 11555 1985 12380 2000
rect 12410 1985 12460 2000
rect 12490 2000 12495 2015
rect 13310 2000 13315 2015
rect 12490 1985 13235 2000
rect 13265 1985 13315 2000
rect 13345 2000 13350 2015
rect 13345 1985 13680 2000
rect 485 1275 490 1305
rect 520 1275 525 1305
rect 1180 1290 1345 1305
rect 1340 1275 1345 1290
rect 1375 1275 1380 1305
rect 12295 1290 12460 1305
rect 12455 1275 12460 1290
rect 12490 1275 12495 1305
rect 13150 1290 13315 1305
rect 13310 1275 13315 1290
rect 13345 1275 13350 1305
rect 2035 1230 2200 1245
rect 2195 1215 2200 1230
rect 2230 1215 2235 1245
rect 2890 1230 3055 1245
rect 3050 1215 3055 1230
rect 3085 1215 3090 1245
rect 10580 1230 10745 1245
rect 10740 1215 10745 1230
rect 10775 1215 10780 1245
rect 11440 1230 11605 1245
rect 11600 1215 11605 1230
rect 11635 1230 13680 1245
rect 11635 1215 11640 1230
rect 0 1170 3910 1185
rect 3905 1155 3910 1170
rect 3940 1155 3945 1185
rect 9730 1170 9895 1185
rect 9890 1155 9895 1170
rect 9925 1170 13680 1185
rect 9925 1155 9930 1170
rect 0 1110 4070 1125
rect 4600 1110 4765 1125
rect 4760 1095 4765 1110
rect 4795 1095 4800 1125
rect 5455 1110 5620 1125
rect 5615 1095 5620 1110
rect 5650 1095 5655 1125
rect 6310 1110 6475 1125
rect 6470 1095 6475 1110
rect 6505 1095 6510 1125
rect 7165 1110 7330 1125
rect 7325 1095 7330 1110
rect 7360 1095 7365 1125
rect 8020 1110 8185 1125
rect 8180 1095 8185 1110
rect 8215 1095 8220 1125
rect 8875 1110 9040 1125
rect 9035 1095 9040 1110
rect 9070 1110 9175 1125
rect 9070 1095 9075 1110
<< via1 >>
rect 4765 2165 4795 2195
rect 5620 2165 5650 2195
rect 6475 2165 6505 2195
rect 7330 2165 7360 2195
rect 8185 2165 8215 2195
rect 9040 2165 9070 2195
rect 3910 2105 3940 2135
rect 9895 2105 9925 2135
rect 2200 2045 2230 2075
rect 3055 2045 3085 2075
rect 10745 2045 10775 2075
rect 11605 2045 11635 2075
rect 490 1985 520 2015
rect 1345 1985 1375 2015
rect 12460 1985 12490 2015
rect 13315 1985 13345 2015
rect 490 1275 520 1305
rect 1345 1275 1375 1305
rect 12460 1275 12490 1305
rect 13315 1275 13345 1305
rect 2200 1215 2230 1245
rect 3055 1215 3085 1245
rect 10745 1215 10775 1245
rect 11605 1215 11635 1245
rect 3910 1155 3940 1185
rect 9895 1155 9925 1185
rect 4765 1095 4795 1125
rect 5620 1095 5650 1125
rect 6475 1095 6505 1125
rect 7330 1095 7360 1125
rect 8185 1095 8215 1125
rect 9040 1095 9070 1125
<< metal2 >>
rect 4600 2200 4640 2205
rect 4600 2180 4605 2200
rect 0 2170 4605 2180
rect 4635 2170 4640 2200
rect 5455 2200 5495 2205
rect 0 2165 4640 2170
rect 4760 2165 4765 2195
rect 4795 2165 4800 2195
rect 5455 2170 5460 2200
rect 5490 2170 5495 2200
rect 6310 2200 6350 2205
rect 5455 2165 5495 2170
rect 5615 2165 5620 2195
rect 5650 2165 5655 2195
rect 6310 2170 6315 2200
rect 6345 2170 6350 2200
rect 7165 2200 7205 2205
rect 6310 2165 6350 2170
rect 6470 2165 6475 2195
rect 6505 2165 6510 2195
rect 7165 2170 7170 2200
rect 7200 2170 7205 2200
rect 8020 2200 8060 2205
rect 7165 2165 7205 2170
rect 7325 2165 7330 2195
rect 7360 2165 7365 2195
rect 8020 2170 8025 2200
rect 8055 2170 8060 2200
rect 8875 2200 8915 2205
rect 8020 2165 8060 2170
rect 8180 2165 8185 2195
rect 8215 2165 8220 2195
rect 8875 2170 8880 2200
rect 8910 2170 8915 2200
rect 9135 2200 9175 2205
rect 8875 2165 8915 2170
rect 9035 2165 9040 2195
rect 9070 2165 9075 2195
rect 9135 2170 9140 2200
rect 9170 2180 9175 2200
rect 9170 2170 13680 2180
rect 9135 2165 13680 2170
rect 3745 2140 3785 2145
rect 3745 2120 3750 2140
rect 0 2110 3750 2120
rect 3780 2110 3785 2140
rect 0 2105 3785 2110
rect 3905 2105 3910 2135
rect 3940 2105 3945 2135
rect 2035 2080 2075 2085
rect 2035 2060 2040 2080
rect 0 2050 2040 2060
rect 2070 2050 2075 2080
rect 2890 2080 2930 2085
rect 0 2045 2075 2050
rect 2195 2045 2200 2075
rect 2230 2045 2235 2075
rect 2890 2050 2895 2080
rect 2925 2050 2930 2080
rect 2890 2045 2930 2050
rect 3050 2045 3055 2075
rect 3085 2045 3090 2075
rect 325 2020 365 2025
rect 325 2000 330 2020
rect 0 1990 330 2000
rect 360 1990 365 2020
rect 1180 2020 1220 2025
rect 0 1985 365 1990
rect 485 1985 490 2015
rect 520 1985 525 2015
rect 1180 1990 1185 2020
rect 1215 1990 1220 2020
rect 1180 1985 1220 1990
rect 1340 1985 1345 2015
rect 1375 1985 1380 2015
rect 340 1970 355 1985
rect 495 1970 510 1985
rect 1195 1970 1210 1985
rect 1350 1970 1365 1985
rect 2050 1970 2065 2045
rect 2205 1970 2220 2045
rect 2905 1970 2920 2045
rect 3060 1970 3075 2045
rect 3760 1970 3775 2105
rect 3915 1970 3930 2105
rect 4615 1970 4630 2165
rect 4770 1970 4785 2165
rect 5470 1970 5485 2165
rect 5625 1970 5640 2165
rect 6325 1970 6340 2165
rect 6480 1970 6495 2165
rect 7180 1970 7195 2165
rect 7335 1970 7350 2165
rect 8035 1970 8050 2165
rect 8190 1970 8205 2165
rect 8890 1970 8905 2165
rect 9045 1970 9060 2165
rect 9730 2140 9770 2145
rect 9730 2110 9735 2140
rect 9765 2110 9770 2140
rect 9990 2140 10030 2145
rect 9730 2105 9770 2110
rect 9890 2105 9895 2135
rect 9925 2105 9930 2135
rect 9990 2110 9995 2140
rect 10025 2120 10030 2140
rect 10025 2110 13680 2120
rect 9990 2105 13680 2110
rect 9745 1970 9760 2105
rect 9900 1970 9915 2105
rect 10580 2080 10620 2085
rect 10580 2050 10585 2080
rect 10615 2050 10620 2080
rect 11440 2080 11480 2085
rect 10580 2045 10620 2050
rect 10740 2045 10745 2075
rect 10775 2045 10780 2075
rect 11440 2050 11445 2080
rect 11475 2050 11480 2080
rect 11700 2080 11740 2085
rect 11440 2045 11480 2050
rect 11600 2045 11605 2075
rect 11635 2045 11640 2075
rect 11700 2050 11705 2080
rect 11735 2060 11740 2080
rect 11735 2050 13680 2060
rect 11700 2045 13680 2050
rect 10600 1970 10615 2045
rect 10755 1970 10770 2045
rect 11455 1970 11470 2045
rect 11610 1970 11625 2045
rect 12295 2020 12335 2025
rect 12295 1990 12300 2020
rect 12330 1990 12335 2020
rect 13150 2020 13190 2025
rect 12295 1985 12335 1990
rect 12455 1985 12460 2015
rect 12490 1985 12495 2015
rect 13150 1990 13155 2020
rect 13185 1990 13190 2020
rect 13410 2020 13450 2025
rect 13150 1985 13190 1990
rect 13310 1985 13315 2015
rect 13345 1985 13350 2015
rect 13410 1990 13415 2020
rect 13445 2000 13450 2020
rect 13445 1990 13680 2000
rect 13410 1985 13680 1990
rect 12310 1970 12325 1985
rect 12465 1970 12480 1985
rect 13165 1970 13180 1985
rect 13320 1970 13335 1985
rect 340 1305 355 1310
rect 495 1305 510 1310
rect 1195 1305 1210 1310
rect 1350 1305 1365 1310
rect 0 1300 365 1305
rect 0 1290 330 1300
rect 325 1270 330 1290
rect 360 1270 365 1300
rect 485 1275 490 1305
rect 520 1275 525 1305
rect 1180 1300 1220 1305
rect 325 1265 365 1270
rect 1180 1270 1185 1300
rect 1215 1270 1220 1300
rect 1340 1275 1345 1305
rect 1375 1275 1380 1305
rect 1180 1265 1220 1270
rect 2050 1245 2065 1310
rect 2205 1245 2220 1310
rect 2905 1245 2920 1310
rect 3060 1245 3075 1310
rect 0 1240 2075 1245
rect 0 1230 2040 1240
rect 2035 1210 2040 1230
rect 2070 1210 2075 1240
rect 2195 1215 2200 1245
rect 2230 1215 2235 1245
rect 2890 1240 2930 1245
rect 2035 1205 2075 1210
rect 2890 1210 2895 1240
rect 2925 1210 2930 1240
rect 3050 1215 3055 1245
rect 3085 1215 3090 1245
rect 2890 1205 2930 1210
rect 3760 1185 3775 1310
rect 3915 1185 3930 1310
rect 0 1180 3785 1185
rect 0 1170 3750 1180
rect 3745 1150 3750 1170
rect 3780 1150 3785 1180
rect 3905 1155 3910 1185
rect 3940 1155 3945 1185
rect 3745 1145 3785 1150
rect 4615 1125 4630 1310
rect 4770 1125 4785 1310
rect 5470 1125 5485 1310
rect 5625 1125 5640 1310
rect 6325 1125 6340 1310
rect 6480 1125 6495 1310
rect 7180 1125 7195 1310
rect 7335 1125 7350 1310
rect 8035 1125 8050 1310
rect 8190 1125 8205 1310
rect 8890 1125 8905 1310
rect 9045 1125 9060 1310
rect 9745 1185 9760 1310
rect 9900 1185 9915 1310
rect 10600 1245 10615 1310
rect 10755 1245 10770 1310
rect 11455 1245 11470 1310
rect 11610 1245 11625 1310
rect 12310 1305 12325 1310
rect 12465 1305 12480 1310
rect 13165 1305 13180 1310
rect 13320 1305 13335 1310
rect 12295 1300 12335 1305
rect 12295 1270 12300 1300
rect 12330 1270 12335 1300
rect 12455 1275 12460 1305
rect 12490 1275 12495 1305
rect 13150 1300 13190 1305
rect 12295 1265 12335 1270
rect 13150 1270 13155 1300
rect 13185 1270 13190 1300
rect 13310 1275 13315 1305
rect 13345 1275 13350 1305
rect 13410 1300 13680 1305
rect 13150 1265 13190 1270
rect 13410 1270 13415 1300
rect 13445 1290 13680 1300
rect 13445 1270 13450 1290
rect 13410 1265 13450 1270
rect 10580 1240 10620 1245
rect 10580 1210 10585 1240
rect 10615 1210 10620 1240
rect 10740 1215 10745 1245
rect 10775 1215 10780 1245
rect 11440 1240 11480 1245
rect 10580 1205 10620 1210
rect 11440 1210 11445 1240
rect 11475 1210 11480 1240
rect 11600 1215 11605 1245
rect 11635 1215 11640 1245
rect 11700 1240 13680 1245
rect 11440 1205 11480 1210
rect 11700 1210 11705 1240
rect 11735 1230 13680 1240
rect 11735 1210 11740 1230
rect 11700 1205 11740 1210
rect 9730 1180 9770 1185
rect 9730 1150 9735 1180
rect 9765 1150 9770 1180
rect 9890 1155 9895 1185
rect 9925 1155 9930 1185
rect 9990 1180 13680 1185
rect 9730 1145 9770 1150
rect 9990 1150 9995 1180
rect 10025 1170 13680 1180
rect 10025 1150 10030 1170
rect 9990 1145 10030 1150
rect 0 1120 4640 1125
rect 0 1110 4605 1120
rect 4600 1090 4605 1110
rect 4635 1090 4640 1120
rect 4760 1095 4765 1125
rect 4795 1095 4800 1125
rect 5455 1120 5495 1125
rect 4600 1085 4640 1090
rect 5455 1090 5460 1120
rect 5490 1090 5495 1120
rect 5615 1095 5620 1125
rect 5650 1095 5655 1125
rect 6310 1120 6350 1125
rect 5455 1085 5495 1090
rect 6310 1090 6315 1120
rect 6345 1090 6350 1120
rect 6470 1095 6475 1125
rect 6505 1095 6510 1125
rect 7165 1120 7205 1125
rect 6310 1085 6350 1090
rect 7165 1090 7170 1120
rect 7200 1090 7205 1120
rect 7325 1095 7330 1125
rect 7360 1095 7365 1125
rect 8020 1120 8060 1125
rect 7165 1085 7205 1090
rect 8020 1090 8025 1120
rect 8055 1090 8060 1120
rect 8180 1095 8185 1125
rect 8215 1095 8220 1125
rect 8875 1120 8915 1125
rect 8020 1085 8060 1090
rect 8875 1090 8880 1120
rect 8910 1090 8915 1120
rect 9035 1095 9040 1125
rect 9070 1095 9075 1125
rect 9135 1120 13680 1125
rect 8875 1085 8915 1090
rect 9135 1090 9140 1120
rect 9170 1110 13680 1120
rect 9170 1090 9175 1110
rect 9135 1085 9175 1090
<< via2 >>
rect 4605 2170 4635 2200
rect 5460 2170 5490 2200
rect 6315 2170 6345 2200
rect 7170 2170 7200 2200
rect 8025 2170 8055 2200
rect 8880 2170 8910 2200
rect 9140 2170 9170 2200
rect 3750 2110 3780 2140
rect 2040 2050 2070 2080
rect 2895 2050 2925 2080
rect 330 1990 360 2020
rect 1185 1990 1215 2020
rect 9735 2110 9765 2140
rect 9995 2110 10025 2140
rect 10585 2050 10615 2080
rect 11445 2050 11475 2080
rect 11705 2050 11735 2080
rect 12300 1990 12330 2020
rect 13155 1990 13185 2020
rect 13415 1990 13445 2020
rect 330 1270 360 1300
rect 1185 1270 1215 1300
rect 2040 1210 2070 1240
rect 2895 1210 2925 1240
rect 3750 1150 3780 1180
rect 12300 1270 12330 1300
rect 13155 1270 13185 1300
rect 13415 1270 13445 1300
rect 10585 1210 10615 1240
rect 11445 1210 11475 1240
rect 11705 1210 11735 1240
rect 9735 1150 9765 1180
rect 9995 1150 10025 1180
rect 4605 1090 4635 1120
rect 5460 1090 5490 1120
rect 6315 1090 6345 1120
rect 7170 1090 7200 1120
rect 8025 1090 8055 1120
rect 8880 1090 8910 1120
rect 9140 1090 9170 1120
<< metal3 >>
rect 4600 2200 4640 2205
rect 4600 2170 4605 2200
rect 4635 2195 4640 2200
rect 5455 2200 5495 2205
rect 5455 2195 5460 2200
rect 4635 2170 5460 2195
rect 5490 2195 5495 2200
rect 6310 2200 6350 2205
rect 6310 2195 6315 2200
rect 5490 2170 6315 2195
rect 6345 2195 6350 2200
rect 7165 2200 7205 2205
rect 7165 2195 7170 2200
rect 6345 2170 7170 2195
rect 7200 2195 7205 2200
rect 8020 2200 8060 2205
rect 8020 2195 8025 2200
rect 7200 2170 8025 2195
rect 8055 2195 8060 2200
rect 8875 2200 8915 2205
rect 8875 2195 8880 2200
rect 8055 2170 8880 2195
rect 8910 2195 8915 2200
rect 9135 2200 9175 2205
rect 9135 2195 9140 2200
rect 8910 2170 9140 2195
rect 9170 2170 9175 2200
rect 4600 2165 9175 2170
rect 3745 2140 3785 2145
rect 3745 2110 3750 2140
rect 3780 2135 3785 2140
rect 9730 2140 9770 2145
rect 9730 2135 9735 2140
rect 3780 2110 9735 2135
rect 9765 2135 9770 2140
rect 9990 2140 10030 2145
rect 9990 2135 9995 2140
rect 9765 2110 9995 2135
rect 10025 2110 10030 2140
rect 3745 2105 10030 2110
rect 2035 2080 2075 2085
rect 2035 2050 2040 2080
rect 2070 2075 2075 2080
rect 2890 2080 2930 2085
rect 2890 2075 2895 2080
rect 2070 2050 2895 2075
rect 2925 2075 2930 2080
rect 10580 2080 10620 2085
rect 10580 2075 10585 2080
rect 2925 2050 10585 2075
rect 10615 2075 10620 2080
rect 11440 2080 11480 2085
rect 11440 2075 11445 2080
rect 10615 2050 11445 2075
rect 11475 2075 11480 2080
rect 11700 2080 11740 2085
rect 11700 2075 11705 2080
rect 11475 2050 11705 2075
rect 11735 2050 11740 2080
rect 2035 2045 11740 2050
rect 325 2020 365 2025
rect 325 1990 330 2020
rect 360 2015 365 2020
rect 1180 2020 1220 2025
rect 1180 2015 1185 2020
rect 360 1990 1185 2015
rect 1215 2015 1220 2020
rect 12295 2020 12335 2025
rect 12295 2015 12300 2020
rect 1215 1990 12300 2015
rect 12330 2015 12335 2020
rect 13150 2020 13190 2025
rect 13150 2015 13155 2020
rect 12330 1990 13155 2015
rect 13185 2015 13190 2020
rect 13410 2020 13450 2025
rect 13410 2015 13415 2020
rect 13185 1990 13415 2015
rect 13445 1990 13450 2020
rect 325 1985 13450 1990
rect 325 1300 13450 1305
rect 325 1270 330 1300
rect 360 1275 1185 1300
rect 360 1270 365 1275
rect 325 1265 365 1270
rect 1180 1270 1185 1275
rect 1215 1275 12300 1300
rect 1215 1270 1220 1275
rect 1180 1265 1220 1270
rect 12295 1270 12300 1275
rect 12330 1275 13155 1300
rect 12330 1270 12335 1275
rect 12295 1265 12335 1270
rect 13150 1270 13155 1275
rect 13185 1275 13415 1300
rect 13185 1270 13190 1275
rect 13150 1265 13190 1270
rect 13410 1270 13415 1275
rect 13445 1270 13450 1300
rect 13410 1265 13450 1270
rect 2035 1240 11740 1245
rect 2035 1210 2040 1240
rect 2070 1215 2895 1240
rect 2070 1210 2075 1215
rect 2035 1205 2075 1210
rect 2890 1210 2895 1215
rect 2925 1215 10585 1240
rect 2925 1210 2930 1215
rect 2890 1205 2930 1210
rect 10580 1210 10585 1215
rect 10615 1215 11445 1240
rect 10615 1210 10620 1215
rect 10580 1205 10620 1210
rect 11440 1210 11445 1215
rect 11475 1215 11705 1240
rect 11475 1210 11480 1215
rect 11440 1205 11480 1210
rect 11700 1210 11705 1215
rect 11735 1210 11740 1240
rect 11700 1205 11740 1210
rect 3745 1180 10030 1185
rect 3745 1150 3750 1180
rect 3780 1155 9735 1180
rect 3780 1150 3785 1155
rect 3745 1145 3785 1150
rect 9730 1150 9735 1155
rect 9765 1155 9995 1180
rect 9765 1150 9770 1155
rect 9730 1145 9770 1150
rect 9990 1150 9995 1155
rect 10025 1150 10030 1180
rect 9990 1145 10030 1150
rect 4600 1120 9175 1125
rect 4600 1090 4605 1120
rect 4635 1095 5460 1120
rect 4635 1090 4640 1095
rect 4600 1085 4640 1090
rect 5455 1090 5460 1095
rect 5490 1095 6315 1120
rect 5490 1090 5495 1095
rect 5455 1085 5495 1090
rect 6310 1090 6315 1095
rect 6345 1095 7170 1120
rect 6345 1090 6350 1095
rect 6310 1085 6350 1090
rect 7165 1090 7170 1095
rect 7200 1095 8025 1120
rect 7200 1090 7205 1095
rect 7165 1085 7205 1090
rect 8020 1090 8025 1095
rect 8055 1095 8880 1120
rect 8055 1090 8060 1095
rect 8020 1085 8060 1090
rect 8875 1090 8880 1095
rect 8910 1095 9140 1120
rect 8910 1090 8915 1095
rect 8875 1085 8915 1090
rect 9135 1090 9140 1095
rect 9170 1090 9175 1120
rect 9135 1085 9175 1090
use 8_cap_array_final  8_cap_array_final_0
timestamp 1730665161
transform 1 0 65 0 1 115
box -65 -115 6775 2245
use 8_cap_array_final  8_cap_array_final_1
timestamp 1730665161
transform 1 0 6905 0 1 115
box -65 -115 6775 2245
<< end >>
