magic
tech sky130A
timestamp 1730665161
<< metal1 >>
rect 3905 2060 3910 2075
rect 0 2045 3910 2060
rect 3940 2045 3945 2075
rect 4760 2060 4765 2075
rect 4600 2045 4765 2060
rect 4795 2045 4800 2075
rect 5615 2060 5620 2075
rect 5455 2045 5620 2060
rect 5650 2045 5655 2075
rect 6470 2060 6475 2075
rect 6310 2045 6475 2060
rect 6505 2045 6510 2075
rect 7325 2060 7330 2075
rect 7165 2045 7330 2060
rect 7360 2045 7365 2075
rect 8180 2060 8185 2075
rect 8020 2045 8185 2060
rect 8215 2045 8220 2075
rect 9035 2060 9040 2075
rect 8875 2045 9040 2060
rect 9070 2045 9075 2075
rect 9890 2060 9895 2075
rect 9730 2045 9895 2060
rect 9925 2045 9930 2075
rect 485 2000 490 2015
rect 325 1985 490 2000
rect 520 1985 525 2015
rect 1340 2000 1345 2015
rect 1180 1985 1345 2000
rect 1375 1985 1380 2015
rect 2195 2000 2200 2015
rect 2035 1985 2200 2000
rect 2230 1985 2235 2015
rect 3050 2000 3055 2015
rect 2890 1985 3055 2000
rect 3085 1985 3090 2015
rect 10745 2000 10750 2015
rect 10585 1985 10750 2000
rect 10780 1985 10785 2015
rect 11600 2000 11605 2015
rect 11440 1985 11605 2000
rect 11635 1985 11640 2015
rect 12455 2000 12460 2015
rect 12295 1985 12460 2000
rect 12490 1985 12495 2015
rect 13310 1985 13315 2015
rect 13345 1985 13350 2015
rect 0 1290 490 1305
rect 485 1275 490 1290
rect 520 1290 1345 1305
rect 520 1275 525 1290
rect 1340 1275 1345 1290
rect 1375 1290 2200 1305
rect 1375 1275 1380 1290
rect 2195 1275 2200 1290
rect 2230 1290 3055 1305
rect 2230 1275 2235 1290
rect 3050 1275 3055 1290
rect 3085 1290 10750 1305
rect 3085 1275 3090 1290
rect 10745 1275 10750 1290
rect 10780 1290 11605 1305
rect 10780 1275 10785 1290
rect 11600 1275 11605 1290
rect 11635 1290 12460 1305
rect 11635 1275 11640 1290
rect 12455 1275 12460 1290
rect 12490 1290 13315 1305
rect 12490 1275 12495 1290
rect 13310 1275 13315 1290
rect 13345 1290 13680 1305
rect 13345 1275 13350 1290
rect 0 1230 3910 1245
rect 3905 1215 3910 1230
rect 3940 1230 4765 1245
rect 3940 1215 3945 1230
rect 4760 1215 4765 1230
rect 4795 1230 5620 1245
rect 4795 1215 4800 1230
rect 5615 1215 5620 1230
rect 5650 1230 6475 1245
rect 5650 1215 5655 1230
rect 6470 1215 6475 1230
rect 6505 1230 7330 1245
rect 6505 1215 6510 1230
rect 7325 1215 7330 1230
rect 7360 1230 8185 1245
rect 7360 1215 7365 1230
rect 8180 1215 8185 1230
rect 8215 1230 9040 1245
rect 8215 1215 8220 1230
rect 9035 1215 9040 1230
rect 9070 1230 9895 1245
rect 9070 1215 9075 1230
rect 9890 1215 9895 1230
rect 9925 1230 13680 1245
rect 9925 1215 9930 1230
<< via1 >>
rect 3910 2045 3940 2075
rect 4765 2045 4795 2075
rect 5620 2045 5650 2075
rect 6475 2045 6505 2075
rect 7330 2045 7360 2075
rect 8185 2045 8215 2075
rect 9040 2045 9070 2075
rect 9895 2045 9925 2075
rect 490 1985 520 2015
rect 1345 1985 1375 2015
rect 2200 1985 2230 2015
rect 3055 1985 3085 2015
rect 10750 1985 10780 2015
rect 11605 1985 11635 2015
rect 12460 1985 12490 2015
rect 13315 1985 13345 2015
rect 490 1275 520 1305
rect 1345 1275 1375 1305
rect 2200 1275 2230 1305
rect 3055 1275 3085 1305
rect 10750 1275 10780 1305
rect 11605 1275 11635 1305
rect 12460 1275 12490 1305
rect 13315 1275 13345 1305
rect 3910 1215 3940 1245
rect 4765 1215 4795 1245
rect 5620 1215 5650 1245
rect 6475 1215 6505 1245
rect 7330 1215 7360 1245
rect 8185 1215 8215 1245
rect 9040 1215 9070 1245
rect 9895 1215 9925 1245
<< metal2 >>
rect 3745 2080 3785 2085
rect 3745 2060 3750 2080
rect 0 2050 3750 2060
rect 3780 2050 3785 2080
rect 4600 2080 4640 2085
rect 0 2045 3785 2050
rect 3905 2045 3910 2075
rect 3940 2045 3945 2075
rect 4600 2050 4605 2080
rect 4635 2050 4640 2080
rect 5455 2080 5495 2085
rect 4600 2045 4640 2050
rect 4760 2045 4765 2075
rect 4795 2045 4800 2075
rect 5455 2050 5460 2080
rect 5490 2050 5495 2080
rect 6310 2080 6350 2085
rect 5455 2045 5495 2050
rect 5615 2045 5620 2075
rect 5650 2045 5655 2075
rect 6310 2050 6315 2080
rect 6345 2050 6350 2080
rect 7165 2080 7205 2085
rect 6310 2045 6350 2050
rect 6470 2045 6475 2075
rect 6505 2045 6510 2075
rect 7165 2050 7170 2080
rect 7200 2050 7205 2080
rect 8020 2080 8060 2085
rect 7165 2045 7205 2050
rect 7325 2045 7330 2075
rect 7360 2045 7365 2075
rect 8020 2050 8025 2080
rect 8055 2050 8060 2080
rect 8875 2080 8915 2085
rect 8020 2045 8060 2050
rect 8180 2045 8185 2075
rect 8215 2045 8220 2075
rect 8875 2050 8880 2080
rect 8910 2050 8915 2080
rect 9730 2080 9770 2085
rect 8875 2045 8915 2050
rect 9035 2045 9040 2075
rect 9070 2045 9075 2075
rect 9730 2050 9735 2080
rect 9765 2050 9770 2080
rect 9990 2080 10030 2085
rect 9730 2045 9770 2050
rect 9890 2045 9895 2075
rect 9925 2045 9930 2075
rect 9990 2050 9995 2080
rect 10025 2060 10030 2080
rect 10025 2050 13680 2060
rect 9990 2045 13680 2050
rect 325 2020 365 2025
rect 325 2000 330 2020
rect 0 1990 330 2000
rect 360 1990 365 2020
rect 1180 2020 1220 2025
rect 0 1985 365 1990
rect 485 1985 490 2015
rect 520 1985 525 2015
rect 1180 1990 1185 2020
rect 1215 1990 1220 2020
rect 2035 2020 2075 2025
rect 1180 1985 1220 1990
rect 1340 1985 1345 2015
rect 1375 1985 1380 2015
rect 2035 1990 2040 2020
rect 2070 1990 2075 2020
rect 2890 2020 2930 2025
rect 2035 1985 2075 1990
rect 2195 1985 2200 2015
rect 2230 1985 2235 2015
rect 2890 1990 2895 2020
rect 2925 1990 2930 2020
rect 2890 1985 2930 1990
rect 3050 1985 3055 2015
rect 3085 1985 3090 2015
rect 340 1980 355 1985
rect 495 1980 510 1985
rect 1195 1980 1210 1985
rect 1350 1980 1365 1985
rect 2050 1980 2065 1985
rect 2205 1980 2220 1985
rect 2905 1980 2920 1985
rect 3060 1980 3075 1985
rect 3760 1980 3775 2045
rect 3915 1980 3930 2045
rect 4615 1980 4630 2045
rect 4770 1980 4785 2045
rect 5470 1980 5485 2045
rect 5625 1980 5640 2045
rect 6325 1980 6340 2045
rect 6480 1980 6495 2045
rect 7180 1980 7195 2045
rect 7335 1980 7350 2045
rect 8035 1980 8050 2045
rect 8190 1980 8205 2045
rect 8890 1980 8905 2045
rect 9045 1980 9060 2045
rect 9745 1980 9760 2045
rect 9900 1980 9915 2045
rect 10585 2020 10625 2025
rect 10585 1990 10590 2020
rect 10620 1990 10625 2020
rect 11440 2020 11480 2025
rect 10585 1985 10625 1990
rect 10745 1985 10750 2015
rect 10780 1985 10785 2015
rect 11440 1990 11445 2020
rect 11475 1990 11480 2020
rect 12295 2020 12335 2025
rect 11440 1985 11480 1990
rect 11600 1985 11605 2015
rect 11635 1985 11640 2015
rect 12295 1990 12300 2020
rect 12330 1990 12335 2020
rect 13150 2020 13190 2025
rect 12295 1985 12335 1990
rect 12455 1985 12460 2015
rect 12490 1985 12495 2015
rect 13150 1990 13155 2020
rect 13185 1990 13190 2020
rect 13410 2020 13450 2025
rect 13150 1985 13190 1990
rect 13310 1985 13315 2015
rect 13345 1985 13350 2015
rect 13410 1990 13415 2020
rect 13445 2000 13450 2020
rect 13445 1990 13680 2000
rect 13410 1985 13680 1990
rect 10600 1980 10615 1985
rect 10755 1980 10770 1985
rect 11455 1980 11470 1985
rect 11610 1980 11625 1985
rect 12310 1980 12325 1985
rect 12465 1980 12480 1985
rect 13165 1980 13180 1985
rect 13320 1980 13335 1985
rect 340 1305 355 1320
rect 495 1305 510 1320
rect 1195 1305 1210 1320
rect 1350 1305 1365 1320
rect 2050 1305 2065 1320
rect 2205 1305 2220 1320
rect 2905 1305 2920 1320
rect 3060 1305 3075 1320
rect 0 1300 365 1305
rect 0 1290 330 1300
rect 325 1270 330 1290
rect 360 1270 365 1300
rect 485 1275 490 1305
rect 520 1275 525 1305
rect 1180 1300 1220 1305
rect 325 1265 365 1270
rect 1180 1270 1185 1300
rect 1215 1270 1220 1300
rect 1340 1275 1345 1305
rect 1375 1275 1380 1305
rect 2035 1300 2075 1305
rect 1180 1265 1220 1270
rect 2035 1270 2040 1300
rect 2070 1270 2075 1300
rect 2195 1275 2200 1305
rect 2230 1275 2235 1305
rect 2890 1300 2930 1305
rect 2035 1265 2075 1270
rect 2890 1270 2895 1300
rect 2925 1270 2930 1300
rect 3050 1275 3055 1305
rect 3085 1275 3090 1305
rect 2890 1265 2930 1270
rect 3760 1245 3775 1320
rect 3915 1245 3930 1320
rect 4615 1245 4630 1320
rect 4770 1245 4785 1320
rect 5470 1245 5485 1320
rect 5625 1245 5640 1320
rect 6325 1245 6340 1320
rect 6480 1245 6495 1320
rect 7180 1245 7195 1320
rect 7335 1245 7350 1320
rect 8035 1245 8050 1320
rect 8190 1245 8205 1320
rect 8890 1245 8905 1320
rect 9045 1245 9060 1320
rect 9745 1245 9760 1320
rect 9900 1245 9915 1320
rect 10600 1305 10615 1320
rect 10755 1305 10770 1320
rect 11455 1305 11470 1320
rect 11610 1305 11625 1320
rect 12310 1305 12325 1320
rect 12465 1305 12480 1320
rect 13165 1305 13180 1320
rect 13320 1305 13335 1320
rect 10585 1300 10625 1305
rect 10585 1270 10590 1300
rect 10620 1270 10625 1300
rect 10745 1275 10750 1305
rect 10780 1275 10785 1305
rect 11440 1300 11480 1305
rect 10585 1265 10625 1270
rect 11440 1270 11445 1300
rect 11475 1270 11480 1300
rect 11600 1275 11605 1305
rect 11635 1275 11640 1305
rect 12295 1300 12335 1305
rect 11440 1265 11480 1270
rect 12295 1270 12300 1300
rect 12330 1270 12335 1300
rect 12455 1275 12460 1305
rect 12490 1275 12495 1305
rect 13150 1300 13190 1305
rect 12295 1265 12335 1270
rect 13150 1270 13155 1300
rect 13185 1270 13190 1300
rect 13310 1275 13315 1305
rect 13345 1275 13350 1305
rect 13410 1300 13680 1305
rect 13150 1265 13190 1270
rect 13410 1270 13415 1300
rect 13445 1290 13680 1300
rect 13445 1270 13450 1290
rect 13410 1265 13450 1270
rect 0 1240 3785 1245
rect 0 1230 3750 1240
rect 3745 1210 3750 1230
rect 3780 1210 3785 1240
rect 3905 1215 3910 1245
rect 3940 1215 3945 1245
rect 4600 1240 4640 1245
rect 3745 1205 3785 1210
rect 4600 1210 4605 1240
rect 4635 1210 4640 1240
rect 4760 1215 4765 1245
rect 4795 1215 4800 1245
rect 5455 1240 5495 1245
rect 4600 1205 4640 1210
rect 5455 1210 5460 1240
rect 5490 1210 5495 1240
rect 5615 1215 5620 1245
rect 5650 1215 5655 1245
rect 6310 1240 6350 1245
rect 5455 1205 5495 1210
rect 6310 1210 6315 1240
rect 6345 1210 6350 1240
rect 6470 1215 6475 1245
rect 6505 1215 6510 1245
rect 7165 1240 7205 1245
rect 6310 1205 6350 1210
rect 7165 1210 7170 1240
rect 7200 1210 7205 1240
rect 7325 1215 7330 1245
rect 7360 1215 7365 1245
rect 8020 1240 8060 1245
rect 7165 1205 7205 1210
rect 8020 1210 8025 1240
rect 8055 1210 8060 1240
rect 8180 1215 8185 1245
rect 8215 1215 8220 1245
rect 8875 1240 8915 1245
rect 8020 1205 8060 1210
rect 8875 1210 8880 1240
rect 8910 1210 8915 1240
rect 9035 1215 9040 1245
rect 9070 1215 9075 1245
rect 9730 1240 9770 1245
rect 8875 1205 8915 1210
rect 9730 1210 9735 1240
rect 9765 1210 9770 1240
rect 9890 1215 9895 1245
rect 9925 1215 9930 1245
rect 9990 1240 13680 1245
rect 9730 1205 9770 1210
rect 9990 1210 9995 1240
rect 10025 1230 13680 1240
rect 10025 1210 10030 1230
rect 9990 1205 10030 1210
<< via2 >>
rect 3750 2050 3780 2080
rect 4605 2050 4635 2080
rect 5460 2050 5490 2080
rect 6315 2050 6345 2080
rect 7170 2050 7200 2080
rect 8025 2050 8055 2080
rect 8880 2050 8910 2080
rect 9735 2050 9765 2080
rect 9995 2050 10025 2080
rect 330 1990 360 2020
rect 1185 1990 1215 2020
rect 2040 1990 2070 2020
rect 2895 1990 2925 2020
rect 10590 1990 10620 2020
rect 11445 1990 11475 2020
rect 12300 1990 12330 2020
rect 13155 1990 13185 2020
rect 13415 1990 13445 2020
rect 330 1270 360 1300
rect 1185 1270 1215 1300
rect 2040 1270 2070 1300
rect 2895 1270 2925 1300
rect 10590 1270 10620 1300
rect 11445 1270 11475 1300
rect 12300 1270 12330 1300
rect 13155 1270 13185 1300
rect 13415 1270 13445 1300
rect 3750 1210 3780 1240
rect 4605 1210 4635 1240
rect 5460 1210 5490 1240
rect 6315 1210 6345 1240
rect 7170 1210 7200 1240
rect 8025 1210 8055 1240
rect 8880 1210 8910 1240
rect 9735 1210 9765 1240
rect 9995 1210 10025 1240
<< metal3 >>
rect 3745 2080 3785 2085
rect 3745 2050 3750 2080
rect 3780 2075 3785 2080
rect 4600 2080 4640 2085
rect 4600 2075 4605 2080
rect 3780 2050 4605 2075
rect 4635 2075 4640 2080
rect 5455 2080 5495 2085
rect 5455 2075 5460 2080
rect 4635 2050 5460 2075
rect 5490 2075 5495 2080
rect 6310 2080 6350 2085
rect 6310 2075 6315 2080
rect 5490 2050 6315 2075
rect 6345 2075 6350 2080
rect 7165 2080 7205 2085
rect 7165 2075 7170 2080
rect 6345 2050 7170 2075
rect 7200 2075 7205 2080
rect 8020 2080 8060 2085
rect 8020 2075 8025 2080
rect 7200 2050 8025 2075
rect 8055 2075 8060 2080
rect 8875 2080 8915 2085
rect 8875 2075 8880 2080
rect 8055 2050 8880 2075
rect 8910 2075 8915 2080
rect 9730 2080 9770 2085
rect 9730 2075 9735 2080
rect 8910 2050 9735 2075
rect 9765 2075 9770 2080
rect 9990 2080 10030 2085
rect 9990 2075 9995 2080
rect 9765 2050 9995 2075
rect 10025 2050 10030 2080
rect 3745 2045 10030 2050
rect 325 2020 365 2025
rect 325 1990 330 2020
rect 360 2015 365 2020
rect 1180 2020 1220 2025
rect 1180 2015 1185 2020
rect 360 1990 1185 2015
rect 1215 2015 1220 2020
rect 2035 2020 2075 2025
rect 2035 2015 2040 2020
rect 1215 1990 2040 2015
rect 2070 2015 2075 2020
rect 2890 2020 2930 2025
rect 2890 2015 2895 2020
rect 2070 1990 2895 2015
rect 2925 2015 2930 2020
rect 10585 2020 10625 2025
rect 10585 2015 10590 2020
rect 2925 1990 10590 2015
rect 10620 2015 10625 2020
rect 11440 2020 11480 2025
rect 11440 2015 11445 2020
rect 10620 1990 11445 2015
rect 11475 2015 11480 2020
rect 12295 2020 12335 2025
rect 12295 2015 12300 2020
rect 11475 1990 12300 2015
rect 12330 2015 12335 2020
rect 13150 2020 13190 2025
rect 13150 2015 13155 2020
rect 12330 1990 13155 2015
rect 13185 2015 13190 2020
rect 13410 2020 13450 2025
rect 13410 2015 13415 2020
rect 13185 1990 13415 2015
rect 13445 1990 13450 2020
rect 325 1985 13450 1990
rect 325 1300 13450 1305
rect 325 1270 330 1300
rect 360 1275 1185 1300
rect 360 1270 365 1275
rect 325 1265 365 1270
rect 1180 1270 1185 1275
rect 1215 1275 2040 1300
rect 1215 1270 1220 1275
rect 1180 1265 1220 1270
rect 2035 1270 2040 1275
rect 2070 1275 2895 1300
rect 2070 1270 2075 1275
rect 2035 1265 2075 1270
rect 2890 1270 2895 1275
rect 2925 1275 10590 1300
rect 2925 1270 2930 1275
rect 2890 1265 2930 1270
rect 10585 1270 10590 1275
rect 10620 1275 11445 1300
rect 10620 1270 10625 1275
rect 10585 1265 10625 1270
rect 11440 1270 11445 1275
rect 11475 1275 12300 1300
rect 11475 1270 11480 1275
rect 11440 1265 11480 1270
rect 12295 1270 12300 1275
rect 12330 1275 13155 1300
rect 12330 1270 12335 1275
rect 12295 1265 12335 1270
rect 13150 1270 13155 1275
rect 13185 1275 13415 1300
rect 13185 1270 13190 1275
rect 13150 1265 13190 1270
rect 13410 1270 13415 1275
rect 13445 1270 13450 1300
rect 13410 1265 13450 1270
rect 3745 1240 10030 1245
rect 3745 1210 3750 1240
rect 3780 1215 4605 1240
rect 3780 1210 3785 1215
rect 3745 1205 3785 1210
rect 4600 1210 4605 1215
rect 4635 1215 5460 1240
rect 4635 1210 4640 1215
rect 4600 1205 4640 1210
rect 5455 1210 5460 1215
rect 5490 1215 6315 1240
rect 5490 1210 5495 1215
rect 5455 1205 5495 1210
rect 6310 1210 6315 1215
rect 6345 1215 7170 1240
rect 6345 1210 6350 1215
rect 6310 1205 6350 1210
rect 7165 1210 7170 1215
rect 7200 1215 8025 1240
rect 7200 1210 7205 1215
rect 7165 1205 7205 1210
rect 8020 1210 8025 1215
rect 8055 1215 8880 1240
rect 8055 1210 8060 1215
rect 8020 1205 8060 1210
rect 8875 1210 8880 1215
rect 8910 1215 9735 1240
rect 8910 1210 8915 1215
rect 8875 1205 8915 1210
rect 9730 1210 9735 1215
rect 9765 1215 9995 1240
rect 9765 1210 9770 1215
rect 9730 1205 9770 1210
rect 9990 1210 9995 1215
rect 10025 1210 10030 1240
rect 9990 1205 10030 1210
use 8_cap_array_final  8_cap_array_final_0
timestamp 1730665161
transform 1 0 65 0 1 115
box -65 -115 6775 2245
use 8_cap_array_final  8_cap_array_final_1
timestamp 1730665161
transform 1 0 6905 0 1 115
box -65 -115 6775 2245
<< end >>
