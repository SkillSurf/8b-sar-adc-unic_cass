magic
tech sky130A
timestamp 1730665161
<< metal1 >>
rect 485 1985 490 2015
rect 520 1985 525 2015
rect 1340 2000 1345 2015
rect 1180 1985 1345 2000
rect 1375 1985 1380 2015
rect 2195 2000 2200 2015
rect 2035 1985 2200 2000
rect 2230 1985 2235 2015
rect 3050 2000 3055 2015
rect 2890 1985 3055 2000
rect 3085 1985 3090 2015
rect 3905 2000 3910 2015
rect 3745 1985 3910 2000
rect 3940 1985 3945 2015
rect 4760 2000 4765 2015
rect 4600 1985 4765 2000
rect 4795 1985 4800 2015
rect 5615 2000 5620 2015
rect 5455 1985 5620 2000
rect 5650 1985 5655 2015
rect 6470 2000 6475 2015
rect 6310 1985 6475 2000
rect 6505 1985 6510 2015
rect 7325 2000 7330 2015
rect 7165 1985 7330 2000
rect 7360 1985 7365 2015
rect 8180 2000 8185 2015
rect 8020 1985 8185 2000
rect 8215 1985 8220 2015
rect 9035 2000 9040 2015
rect 8875 1985 9040 2000
rect 9070 1985 9075 2015
rect 9890 2000 9895 2015
rect 9730 1985 9895 2000
rect 9925 1985 9930 2015
rect 10745 2000 10750 2015
rect 10585 1985 10750 2000
rect 10780 1985 10785 2015
rect 11600 2000 11605 2015
rect 11440 1985 11605 2000
rect 11635 1985 11640 2015
rect 12455 2000 12460 2015
rect 12295 1985 12460 2000
rect 12490 1985 12495 2015
rect 13310 2000 13315 2015
rect 13150 1985 13315 2000
rect 13345 1985 13350 2015
rect 0 1290 490 1305
rect 485 1275 490 1290
rect 520 1290 1345 1305
rect 520 1275 525 1290
rect 1340 1275 1345 1290
rect 1375 1290 2200 1305
rect 1375 1275 1380 1290
rect 2195 1275 2200 1290
rect 2230 1290 3055 1305
rect 2230 1275 2235 1290
rect 3050 1275 3055 1290
rect 3085 1290 3910 1305
rect 3085 1275 3090 1290
rect 3905 1275 3910 1290
rect 3940 1290 4765 1305
rect 3940 1275 3945 1290
rect 4760 1275 4765 1290
rect 4795 1290 5620 1305
rect 4795 1275 4800 1290
rect 5615 1275 5620 1290
rect 5650 1290 6475 1305
rect 5650 1275 5655 1290
rect 6470 1275 6475 1290
rect 6505 1290 7330 1305
rect 6505 1275 6510 1290
rect 7325 1275 7330 1290
rect 7360 1290 8185 1305
rect 7360 1275 7365 1290
rect 8180 1275 8185 1290
rect 8215 1290 9040 1305
rect 8215 1275 8220 1290
rect 9035 1275 9040 1290
rect 9070 1290 9895 1305
rect 9070 1275 9075 1290
rect 9890 1275 9895 1290
rect 9925 1290 10750 1305
rect 9925 1275 9930 1290
rect 10745 1275 10750 1290
rect 10780 1290 11605 1305
rect 10780 1275 10785 1290
rect 11600 1275 11605 1290
rect 11635 1290 12460 1305
rect 11635 1275 11640 1290
rect 12455 1275 12460 1290
rect 12490 1290 13315 1305
rect 12490 1275 12495 1290
rect 13310 1275 13315 1290
rect 13345 1290 13680 1305
rect 13345 1275 13350 1290
<< via1 >>
rect 490 1985 520 2015
rect 1345 1985 1375 2015
rect 2200 1985 2230 2015
rect 3055 1985 3085 2015
rect 3910 1985 3940 2015
rect 4765 1985 4795 2015
rect 5620 1985 5650 2015
rect 6475 1985 6505 2015
rect 7330 1985 7360 2015
rect 8185 1985 8215 2015
rect 9040 1985 9070 2015
rect 9895 1985 9925 2015
rect 10750 1985 10780 2015
rect 11605 1985 11635 2015
rect 12460 1985 12490 2015
rect 13315 1985 13345 2015
rect 490 1275 520 1305
rect 1345 1275 1375 1305
rect 2200 1275 2230 1305
rect 3055 1275 3085 1305
rect 3910 1275 3940 1305
rect 4765 1275 4795 1305
rect 5620 1275 5650 1305
rect 6475 1275 6505 1305
rect 7330 1275 7360 1305
rect 8185 1275 8215 1305
rect 9040 1275 9070 1305
rect 9895 1275 9925 1305
rect 10750 1275 10780 1305
rect 11605 1275 11635 1305
rect 12460 1275 12490 1305
rect 13315 1275 13345 1305
<< metal2 >>
rect 325 2020 365 2025
rect 325 2000 330 2020
rect 0 1990 330 2000
rect 360 1990 365 2020
rect 1180 2020 1220 2025
rect 0 1985 365 1990
rect 485 1985 490 2015
rect 520 1985 525 2015
rect 1180 1990 1185 2020
rect 1215 1990 1220 2020
rect 2035 2020 2075 2025
rect 1180 1985 1220 1990
rect 1340 1985 1345 2015
rect 1375 1985 1380 2015
rect 2035 1990 2040 2020
rect 2070 1990 2075 2020
rect 2890 2020 2930 2025
rect 2035 1985 2075 1990
rect 2195 1985 2200 2015
rect 2230 1985 2235 2015
rect 2890 1990 2895 2020
rect 2925 1990 2930 2020
rect 3745 2020 3785 2025
rect 2890 1985 2930 1990
rect 3050 1985 3055 2015
rect 3085 1985 3090 2015
rect 3745 1990 3750 2020
rect 3780 1990 3785 2020
rect 4600 2020 4640 2025
rect 3745 1985 3785 1990
rect 3905 1985 3910 2015
rect 3940 1985 3945 2015
rect 4600 1990 4605 2020
rect 4635 1990 4640 2020
rect 5455 2020 5495 2025
rect 4600 1985 4640 1990
rect 4760 1985 4765 2015
rect 4795 1985 4800 2015
rect 5455 1990 5460 2020
rect 5490 1990 5495 2020
rect 6310 2020 6350 2025
rect 5455 1985 5495 1990
rect 5615 1985 5620 2015
rect 5650 1985 5655 2015
rect 6310 1990 6315 2020
rect 6345 1990 6350 2020
rect 7165 2020 7205 2025
rect 6310 1985 6350 1990
rect 6470 1985 6475 2015
rect 6505 1985 6510 2015
rect 7165 1990 7170 2020
rect 7200 1990 7205 2020
rect 8020 2020 8060 2025
rect 7165 1985 7205 1990
rect 7325 1985 7330 2015
rect 7360 1985 7365 2015
rect 8020 1990 8025 2020
rect 8055 1990 8060 2020
rect 8875 2020 8915 2025
rect 8020 1985 8060 1990
rect 8180 1985 8185 2015
rect 8215 1985 8220 2015
rect 8875 1990 8880 2020
rect 8910 1990 8915 2020
rect 9730 2020 9770 2025
rect 8875 1985 8915 1990
rect 9035 1985 9040 2015
rect 9070 1985 9075 2015
rect 9730 1990 9735 2020
rect 9765 1990 9770 2020
rect 10585 2020 10625 2025
rect 9730 1985 9770 1990
rect 9890 1985 9895 2015
rect 9925 1985 9930 2015
rect 10585 1990 10590 2020
rect 10620 1990 10625 2020
rect 11440 2020 11480 2025
rect 10585 1985 10625 1990
rect 10745 1985 10750 2015
rect 10780 1985 10785 2015
rect 11440 1990 11445 2020
rect 11475 1990 11480 2020
rect 12295 2020 12335 2025
rect 11440 1985 11480 1990
rect 11600 1985 11605 2015
rect 11635 1985 11640 2015
rect 12295 1990 12300 2020
rect 12330 1990 12335 2020
rect 13150 2020 13190 2025
rect 12295 1985 12335 1990
rect 12455 1985 12460 2015
rect 12490 1985 12495 2015
rect 13150 1990 13155 2020
rect 13185 1990 13190 2020
rect 13410 2020 13450 2025
rect 13150 1985 13190 1990
rect 13310 1985 13315 2015
rect 13345 1985 13350 2015
rect 13410 1990 13415 2020
rect 13445 2000 13450 2020
rect 13445 1990 13680 2000
rect 13410 1985 13680 1990
rect 340 1980 355 1985
rect 495 1980 510 1985
rect 1195 1980 1210 1985
rect 1350 1980 1365 1985
rect 2050 1980 2065 1985
rect 2205 1980 2220 1985
rect 2905 1980 2920 1985
rect 3060 1980 3075 1985
rect 3760 1980 3775 1985
rect 3915 1980 3930 1985
rect 4615 1980 4630 1985
rect 4770 1980 4785 1985
rect 5470 1980 5485 1985
rect 5625 1980 5640 1985
rect 6325 1980 6340 1985
rect 6480 1980 6495 1985
rect 7180 1980 7195 1985
rect 7335 1980 7350 1985
rect 8035 1980 8050 1985
rect 8190 1980 8205 1985
rect 8890 1980 8905 1985
rect 9045 1980 9060 1985
rect 9745 1980 9760 1985
rect 9900 1980 9915 1985
rect 10600 1980 10615 1985
rect 10755 1980 10770 1985
rect 11455 1980 11470 1985
rect 11610 1980 11625 1985
rect 12310 1980 12325 1985
rect 12465 1980 12480 1985
rect 13165 1980 13180 1985
rect 13320 1980 13335 1985
rect 340 1305 355 1320
rect 495 1305 510 1320
rect 1195 1305 1210 1320
rect 1350 1305 1365 1320
rect 2050 1305 2065 1320
rect 2205 1305 2220 1320
rect 2905 1305 2920 1320
rect 3060 1305 3075 1320
rect 3760 1305 3775 1320
rect 3915 1305 3930 1320
rect 4615 1305 4630 1320
rect 4770 1305 4785 1320
rect 5470 1305 5485 1320
rect 5625 1305 5640 1320
rect 6325 1305 6340 1320
rect 6480 1305 6495 1320
rect 7180 1305 7195 1320
rect 7335 1305 7350 1320
rect 8035 1305 8050 1320
rect 8190 1305 8205 1320
rect 8890 1305 8905 1320
rect 9045 1305 9060 1320
rect 9745 1305 9760 1320
rect 9900 1305 9915 1320
rect 10600 1305 10615 1320
rect 10755 1305 10770 1320
rect 11455 1305 11470 1320
rect 11610 1305 11625 1320
rect 12310 1305 12325 1320
rect 12465 1305 12480 1320
rect 13165 1305 13180 1320
rect 13320 1305 13335 1320
rect 0 1300 365 1305
rect 0 1290 330 1300
rect 325 1270 330 1290
rect 360 1270 365 1300
rect 485 1275 490 1305
rect 520 1275 525 1305
rect 1180 1300 1220 1305
rect 325 1265 365 1270
rect 1180 1270 1185 1300
rect 1215 1270 1220 1300
rect 1340 1275 1345 1305
rect 1375 1275 1380 1305
rect 2035 1300 2075 1305
rect 1180 1265 1220 1270
rect 2035 1270 2040 1300
rect 2070 1270 2075 1300
rect 2195 1275 2200 1305
rect 2230 1275 2235 1305
rect 2890 1300 2930 1305
rect 2035 1265 2075 1270
rect 2890 1270 2895 1300
rect 2925 1270 2930 1300
rect 3050 1275 3055 1305
rect 3085 1275 3090 1305
rect 3745 1300 3785 1305
rect 2890 1265 2930 1270
rect 3745 1270 3750 1300
rect 3780 1270 3785 1300
rect 3905 1275 3910 1305
rect 3940 1275 3945 1305
rect 4600 1300 4640 1305
rect 3745 1265 3785 1270
rect 4600 1270 4605 1300
rect 4635 1270 4640 1300
rect 4760 1275 4765 1305
rect 4795 1275 4800 1305
rect 5455 1300 5495 1305
rect 4600 1265 4640 1270
rect 5455 1270 5460 1300
rect 5490 1270 5495 1300
rect 5615 1275 5620 1305
rect 5650 1275 5655 1305
rect 6310 1300 6350 1305
rect 5455 1265 5495 1270
rect 6310 1270 6315 1300
rect 6345 1270 6350 1300
rect 6470 1275 6475 1305
rect 6505 1275 6510 1305
rect 7165 1300 7205 1305
rect 6310 1265 6350 1270
rect 7165 1270 7170 1300
rect 7200 1270 7205 1300
rect 7325 1275 7330 1305
rect 7360 1275 7365 1305
rect 8020 1300 8060 1305
rect 7165 1265 7205 1270
rect 8020 1270 8025 1300
rect 8055 1270 8060 1300
rect 8180 1275 8185 1305
rect 8215 1275 8220 1305
rect 8875 1300 8915 1305
rect 8020 1265 8060 1270
rect 8875 1270 8880 1300
rect 8910 1270 8915 1300
rect 9035 1275 9040 1305
rect 9070 1275 9075 1305
rect 9730 1300 9770 1305
rect 8875 1265 8915 1270
rect 9730 1270 9735 1300
rect 9765 1270 9770 1300
rect 9890 1275 9895 1305
rect 9925 1275 9930 1305
rect 10585 1300 10625 1305
rect 9730 1265 9770 1270
rect 10585 1270 10590 1300
rect 10620 1270 10625 1300
rect 10745 1275 10750 1305
rect 10780 1275 10785 1305
rect 11440 1300 11480 1305
rect 10585 1265 10625 1270
rect 11440 1270 11445 1300
rect 11475 1270 11480 1300
rect 11600 1275 11605 1305
rect 11635 1275 11640 1305
rect 12295 1300 12335 1305
rect 11440 1265 11480 1270
rect 12295 1270 12300 1300
rect 12330 1270 12335 1300
rect 12455 1275 12460 1305
rect 12490 1275 12495 1305
rect 13150 1300 13190 1305
rect 12295 1265 12335 1270
rect 13150 1270 13155 1300
rect 13185 1270 13190 1300
rect 13310 1275 13315 1305
rect 13345 1275 13350 1305
rect 13410 1300 13680 1305
rect 13150 1265 13190 1270
rect 13410 1270 13415 1300
rect 13445 1290 13680 1300
rect 13445 1270 13450 1290
rect 13410 1265 13450 1270
<< via2 >>
rect 330 1990 360 2020
rect 1185 1990 1215 2020
rect 2040 1990 2070 2020
rect 2895 1990 2925 2020
rect 3750 1990 3780 2020
rect 4605 1990 4635 2020
rect 5460 1990 5490 2020
rect 6315 1990 6345 2020
rect 7170 1990 7200 2020
rect 8025 1990 8055 2020
rect 8880 1990 8910 2020
rect 9735 1990 9765 2020
rect 10590 1990 10620 2020
rect 11445 1990 11475 2020
rect 12300 1990 12330 2020
rect 13155 1990 13185 2020
rect 13415 1990 13445 2020
rect 330 1270 360 1300
rect 1185 1270 1215 1300
rect 2040 1270 2070 1300
rect 2895 1270 2925 1300
rect 3750 1270 3780 1300
rect 4605 1270 4635 1300
rect 5460 1270 5490 1300
rect 6315 1270 6345 1300
rect 7170 1270 7200 1300
rect 8025 1270 8055 1300
rect 8880 1270 8910 1300
rect 9735 1270 9765 1300
rect 10590 1270 10620 1300
rect 11445 1270 11475 1300
rect 12300 1270 12330 1300
rect 13155 1270 13185 1300
rect 13415 1270 13445 1300
<< metal3 >>
rect 325 2020 365 2025
rect 325 1990 330 2020
rect 360 2015 365 2020
rect 1180 2020 1220 2025
rect 1180 2015 1185 2020
rect 360 1990 1185 2015
rect 1215 2015 1220 2020
rect 2035 2020 2075 2025
rect 2035 2015 2040 2020
rect 1215 1990 2040 2015
rect 2070 2015 2075 2020
rect 2890 2020 2930 2025
rect 2890 2015 2895 2020
rect 2070 1990 2895 2015
rect 2925 2015 2930 2020
rect 3745 2020 3785 2025
rect 3745 2015 3750 2020
rect 2925 1990 3750 2015
rect 3780 2015 3785 2020
rect 4600 2020 4640 2025
rect 4600 2015 4605 2020
rect 3780 1990 4605 2015
rect 4635 2015 4640 2020
rect 5455 2020 5495 2025
rect 5455 2015 5460 2020
rect 4635 1990 5460 2015
rect 5490 2015 5495 2020
rect 6310 2020 6350 2025
rect 6310 2015 6315 2020
rect 5490 1990 6315 2015
rect 6345 2015 6350 2020
rect 7165 2020 7205 2025
rect 7165 2015 7170 2020
rect 6345 1990 7170 2015
rect 7200 2015 7205 2020
rect 8020 2020 8060 2025
rect 8020 2015 8025 2020
rect 7200 1990 8025 2015
rect 8055 2015 8060 2020
rect 8875 2020 8915 2025
rect 8875 2015 8880 2020
rect 8055 1990 8880 2015
rect 8910 2015 8915 2020
rect 9730 2020 9770 2025
rect 9730 2015 9735 2020
rect 8910 1990 9735 2015
rect 9765 2015 9770 2020
rect 10585 2020 10625 2025
rect 10585 2015 10590 2020
rect 9765 1990 10590 2015
rect 10620 2015 10625 2020
rect 11440 2020 11480 2025
rect 11440 2015 11445 2020
rect 10620 1990 11445 2015
rect 11475 2015 11480 2020
rect 12295 2020 12335 2025
rect 12295 2015 12300 2020
rect 11475 1990 12300 2015
rect 12330 2015 12335 2020
rect 13150 2020 13190 2025
rect 13150 2015 13155 2020
rect 12330 1990 13155 2015
rect 13185 2015 13190 2020
rect 13410 2020 13450 2025
rect 13410 2015 13415 2020
rect 13185 1990 13415 2015
rect 13445 1990 13450 2020
rect 325 1985 13450 1990
rect 325 1300 13450 1305
rect 325 1270 330 1300
rect 360 1275 1185 1300
rect 360 1270 365 1275
rect 325 1265 365 1270
rect 1180 1270 1185 1275
rect 1215 1275 2040 1300
rect 1215 1270 1220 1275
rect 1180 1265 1220 1270
rect 2035 1270 2040 1275
rect 2070 1275 2895 1300
rect 2070 1270 2075 1275
rect 2035 1265 2075 1270
rect 2890 1270 2895 1275
rect 2925 1275 3750 1300
rect 2925 1270 2930 1275
rect 2890 1265 2930 1270
rect 3745 1270 3750 1275
rect 3780 1275 4605 1300
rect 3780 1270 3785 1275
rect 3745 1265 3785 1270
rect 4600 1270 4605 1275
rect 4635 1275 5460 1300
rect 4635 1270 4640 1275
rect 4600 1265 4640 1270
rect 5455 1270 5460 1275
rect 5490 1275 6315 1300
rect 5490 1270 5495 1275
rect 5455 1265 5495 1270
rect 6310 1270 6315 1275
rect 6345 1275 7170 1300
rect 6345 1270 6350 1275
rect 6310 1265 6350 1270
rect 7165 1270 7170 1275
rect 7200 1275 8025 1300
rect 7200 1270 7205 1275
rect 7165 1265 7205 1270
rect 8020 1270 8025 1275
rect 8055 1275 8880 1300
rect 8055 1270 8060 1275
rect 8020 1265 8060 1270
rect 8875 1270 8880 1275
rect 8910 1275 9735 1300
rect 8910 1270 8915 1275
rect 8875 1265 8915 1270
rect 9730 1270 9735 1275
rect 9765 1275 10590 1300
rect 9765 1270 9770 1275
rect 9730 1265 9770 1270
rect 10585 1270 10590 1275
rect 10620 1275 11445 1300
rect 10620 1270 10625 1275
rect 10585 1265 10625 1270
rect 11440 1270 11445 1275
rect 11475 1275 12300 1300
rect 11475 1270 11480 1275
rect 11440 1265 11480 1270
rect 12295 1270 12300 1275
rect 12330 1275 13155 1300
rect 12330 1270 12335 1275
rect 12295 1265 12335 1270
rect 13150 1270 13155 1275
rect 13185 1275 13415 1300
rect 13185 1270 13190 1275
rect 13150 1265 13190 1270
rect 13410 1270 13415 1275
rect 13445 1270 13450 1300
rect 13410 1265 13450 1270
use 8_cap_array_final  8_cap_array_final_0
timestamp 1730665161
transform 1 0 65 0 1 115
box -65 -115 6775 2245
use 8_cap_array_final  8_cap_array_final_1
timestamp 1730665161
transform 1 0 6905 0 1 115
box -65 -115 6775 2245
<< end >>
