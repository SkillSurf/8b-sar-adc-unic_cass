magic
tech sky130A
magscale 1 2
timestamp 1728894068
<< pwell >>
rect 1326 -1043 1408 -1037
rect 1326 -1111 1408 -1049
<< locali >>
rect 1120 -56 1610 -40
rect 1120 -91 1183 -56
rect 1559 -91 1610 -56
rect 1120 -178 1610 -91
rect 1120 -422 1240 -178
rect 1505 -425 1610 -178
rect 1120 -1139 1241 -931
rect 1501 -1139 1610 -929
rect 1120 -1216 1610 -1139
rect 1120 -1252 1155 -1216
rect 1561 -1252 1610 -1216
rect 1120 -1260 1610 -1252
<< viali >>
rect 1183 -91 1559 -56
rect 1155 -1252 1561 -1216
<< metal1 >>
rect 1330 81 1410 90
rect 1330 28 1338 81
rect 1400 28 1410 81
rect 1330 22 1410 28
rect 1120 -56 1610 -40
rect 1120 -91 1183 -56
rect 1559 -91 1610 -56
rect 1120 -100 1610 -91
rect 1320 -219 1420 -210
rect 1320 -272 1336 -219
rect 1402 -272 1420 -219
rect 1320 -280 1420 -272
rect 1300 -630 1345 -504
rect 1387 -510 1432 -504
rect 1387 -570 1430 -510
rect 1270 -700 1345 -630
rect 1300 -830 1345 -700
rect 1386 -630 1430 -570
rect 1386 -700 1460 -630
rect 1386 -770 1430 -700
rect 1387 -830 1430 -770
rect 1328 -1049 1407 -1045
rect 1328 -1050 1335 -1049
rect 1320 -1102 1335 -1050
rect 1401 -1050 1407 -1049
rect 1401 -1102 1410 -1050
rect 1320 -1110 1410 -1102
rect 1120 -1216 1610 -1200
rect 1120 -1252 1155 -1216
rect 1561 -1252 1610 -1216
rect 1120 -1260 1610 -1252
rect 1330 -1324 1400 -1316
rect 1330 -1381 1335 -1324
rect 1398 -1381 1400 -1324
rect 1330 -1390 1400 -1381
<< via1 >>
rect 1338 28 1400 81
rect 1336 -272 1402 -219
rect 1335 -1102 1401 -1049
rect 1335 -1381 1398 -1324
<< metal2 >>
rect 1330 81 1410 90
rect 1330 28 1338 81
rect 1400 28 1410 81
rect 1330 20 1410 28
rect 1350 -210 1380 20
rect 1320 -219 1420 -210
rect 1320 -272 1336 -219
rect 1402 -272 1420 -219
rect 1320 -280 1420 -272
rect 1324 -1049 1410 -1042
rect 1324 -1050 1335 -1049
rect 1320 -1102 1335 -1050
rect 1401 -1102 1410 -1049
rect 1320 -1110 1410 -1102
rect 1350 -1310 1380 -1110
rect 1330 -1324 1400 -1310
rect 1330 -1381 1335 -1324
rect 1398 -1381 1400 -1324
rect 1330 -1390 1400 -1381
use sky130_fd_pr__pfet_01v8_NKK3FE  XM1 ~/saf
timestamp 1728654492
transform 1 0 1369 0 1 -380
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_5WP7M2  XM2 ~/saf
timestamp 1728654492
transform -1 0 1366 0 1 -948
box -211 -279 211 279
<< labels >>
flabel metal1 1330 -1390 1335 -1316 0 FreeSans 256 0 0 0 clk
port 0 nsew
flabel metal1 1386 -770 1430 -570 0 FreeSans 256 0 0 0 vout
port 2 nsew
flabel metal1 1300 -769 1345 -569 0 FreeSans 256 0 0 0 vin
port 3 nsew
flabel metal1 1330 22 1338 90 0 FreeSans 256 0 0 0 clk_b
port 5 nsew
flabel metal1 1120 -100 1178 -40 0 FreeSans 256 0 0 0 vdd
port 4 nsew
flabel metal1 1120 -1260 1180 -1200 0 FreeSans 256 0 0 0 sub
port 1 nsew
<< end >>
